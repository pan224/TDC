

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IyCaF6+6roRR/z73FG9YaF0d7dULyJHX+GoNBLXm93HBP9lCLRfrto6vEw3iGCXzK5VqUo8LUzXz
LNIjSmykCQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ars/zU9oYJUMCyRasaGmgdFnCUXaN3o1oQ0fks4+dXZBJExbjObt0eQ4bTm1Oe0kx7bwkjVYQOv+
UQ7LSA8+pLx+dSrw76W+fhwmbjv8NHk8HXyQr62gS6pGtiXKgK736w7+XTNBA1vQ12Yb/XlI+UNz
IEXEAHZPmFtNRS82+9s=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ypT22bO1Sgj7GXF62sjMcbzRg1ae280bxZhy4N2bQAjzULe/jSsJYy+PGhgDbzqrDKTpXiyDtZkt
oD02eLDdRTGllWcMLfmAbMcheBPHnKTXt9HAhXv063PgOy3UnY+4gioTKkh80haiBvLJgatSPifi
YQpeTG2uJk2s6avI9DDuJWf5ytesbOIq8rdjhkKeFXOVJkRrosfyEugTvccoc1Vbfz7A4F2wgM+D
zQAdcf6ITFXwFESPDeWg0jBH/8FT/oGTumoj/JU8XybS9R37MtI+EqSG5OCB5UPfR7kygCRxMdqx
w9C2YvXXr8F4xw6pVMAzGqjHHzZitlsy10wY2A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iUt+lAN3QxnHPLXCGVB/8iLwL0mQDxrC2eKEtZRQ3tSttWm8FZZIS+L6sXzOYBFdcvxa9yav+Skk
gH0KYhQwN9nPnbBmvq+pv0OWmlNAuJl9BKYeCRvvHDm6ZFmplDtVldoTwk3H3W89FxmDdhSnrp8p
y+EZ4Sey0JKCjHzhKDLb9aiV4K1RcLnUYIHkxt5NRemjZPNHJtaHYmmTYfrufApExkwl0g97mMJh
/9bAzlLXFYd5iRY8cWYOanmNtNy8XdgpYQ9x9FO0bReaxTyYk8KeTd2hcuaOnipXIq1dnLyNcsQ3
oacpKj3c+OCD0yKkipipeAUExSzqLkMixzBzew==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JjEJ4N/hIu1WBDUjIMq9s1GMccDmtrtckrJO9KM4FgsQ0FVnrvs7XLEtH7w3vJEH6mnZFK6gx+Zp
Z6sD/j5+c1FsEF5qvoz8DFaJv1SA0e6R+wJt9JWLiNHRgEY4FWJuMy4GeEzK+JXZXpK3GXkLR7a+
1Q6HsnbRSckp2PGMKP0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KZqHvWv65FrttYAd5GXAxNF6M7H4sPlwsazq1nKQJNzvqECgNuEcm+ZAEJdmD/ayAjxuoA6PeUTI
0DfZA6W/dyVpZBZL701cNaCalR4P8jm9gUNIdKoK9h5ACM0wpchU/5peA9dkp8Q71W1JfJhVf6wV
Pfq6P6zpkxEHamzXVJgMfDIbIUtVkFo5jpozvANXGvZy4NvDF+IkDqh9n1WhJSFw2vSTSWwOc6Os
YPCyiHHgK6fUeo5HsDm8nUZX9YA0YMDCcn+IsvxAoCbVnB8MyuhCLYXxAuS9RlY1JV6hAzEQMCpq
3UPMC6tAiYJyvnJO2Ue+HpfWovjSQbxzMY99PA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vdoPlvKWn5Ji3Xo88zOn99MOAqtEoxjAhuAza+l5LAfqRqsliwhzcGFkAJK4ugd9gKm/M3nHnHPi
/PzAE8cF+f+Utbn8D4EMwG4W0Hif+wOLC02e4qH1wSqAV6WWUm8H7NgadjCJBzXMdZZG7gjGozFv
hvjCKrn45bL0EmR7wl2Q8vZe6J7uihKTYiousdVwB8VF1FLUjPpp6Af2cQmPK82eSrVw0IFHIKqJ
Y/a7ujGEnXPRmoENXb8yibx2IfMb6P5x8SvBxbWHb/Z6q10od4kw4eQyCm6rPn5iaTS1SDweCTJ2
LVJYDuUcJm0TAZrXENpQQfojrfHxe1bol/kUPg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lmo1O/nWVfjvEnWKtJ3RCiwGaUnm3M24qPwY+KlvzkKo4sOFoccG5hcg/sL3BguT2Fqs6upec+/P
lgkR9EpxAHK53ySSYK2Gk+/zJ6wPEAQODMbLtASGTteC4atByoS7g+bnqTV2RCzwQJ8IeLVm63oC
q/A1HmQVWMT63Dha7RRPAWhUKfbQ6Gcxxbrt178CMgNEF8fK64fGKwpKWWGSTZdOuCI6JYCt31CH
jLLgd8XhBzNkjXVlUX1wvTnpXb+ZIkY6TeEL8T+DC3/ZFeM7LEjbf1gPEnDR55V2FW99uqAyh9B+
/sRPnmh44cDlw55G3HMOOIAM5c5/ybP6C+lmBw==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ByXNDvTKDI6gFflyODyOtNqLQFU3tDtRuDnI1QTYGEkfXSRy0PtPqdzLUwZOdH6S+7qVRr5I7hia
BIzMOSTXTbSUeFMET0ea5G6/osyZGxD3vhMq5mc07fbIvonlLCBhXZc9zsxWxmrQIUImWH2twnpK
slu9Wg50/fudlPoBjMVmVGo1w8qzoBi/BwnTzF3og4Q8HdJMlsbKVZ96oAGGsWVhVVGjpde8xZC+
GvqB6jQ2vMmNZJNkyZ47uC4C7nyRet9HhKhT7lFrpKi/HydIDNj30XFaozPxFCtHrnxgGQ0dtM+E
UDFL1fGQBdh4xbe+5S2zrlJKxZ83MLUKUmpM6w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
FQ6jaaUCHb2f5pwzRov4i+aUIFiMKPimy8OY+o+gUz//jjiIaOpD6Fb2xgk2Okc8YooDCJrDYjPb
BF/sRJXAJYwuNhWotzpIrvL2LnFXSbQNxuA2G5QfJ/L3VVwBRS4Erpw4CO/XnekwlWm+Hemw7lmg
TSh+g/2UQMuo1I11X1pur/r2msaXY0AebX28C9COEc0JATSc01E/YXHA+fLu8n+caFcCXRP3+2MP
IlEkaLsCCfoK4ORo/kEhW+F3Bm0Uh54NNOKjxM+QUfzVq9DytNjSvqeZuGQymxo7ErwVBGBpRYA+
ajlSUM37upzcVCH3RfMYB7EutHRnPKlf9eOlUDntgNM120FQd7XBo52pyvu5RMrgjPJDcafK66GF
roZJa7mN8ibREUD/LFm4ey27+sUEgefgixYd25JkaD+lQjTpDGzIcGu6dj/0wIsIwHonuivhvMJT
0hasbkCvom5AvzD3yH9e3VMRBn41Fsy93r+X2Y2u1dn3aR4YrybdDN2do1trqiqbKZ3bWwx7XEZO
EmmPQVaP4kL6P9mVKz6DBxhN9Yl8NVIZhNVwfRmnXpTpIbIFrjIptBkqE/ZhgwepYCslf6K5UfmN
3lp5pBvj+hmlku09FLpFZmlYC4hTUAja6GrdbnPHXwu4CZz5an83bAM50hyawnYUoG8ukdLbUCPu
JOcgeOsjDn6fQggXhE59++WTJX/0S+w5rZ6hjKxolaxrbHng2fr9hippQyAaQ55yMqw8kCIBAYiq
0q1uJPMtorm/BOxYvsubvK1irvXRK2712GZFaCCliO9vF8vjCo1QYonLYXM5Xx38j/31Q8i6xetQ
43FfrNO/8wmfORxW7voqeuJVR1HjU6B4/2cbiCJnBSZv0RekqbuziGtiY7KHmVCxkazDp8Usci2R
QwfcnMkECBuaI12Mrx5EyBXdCWFtyN8AtyoBevYfrbWiuzXFjoCCBCK9XfuG/9D39guhTwVmhCoj
3c4oT6ognOLt8eCp5xVjqgezY4+DLTxGEE1E/PoDOYaS1Mn7bpR+GiPp25tBe8/6MtE4DFlZTdnZ
2trO1KpQM4s4NEPAtx9tNBfO6hfawivn6XCntGPw5/1d7UGx9vKDXbeNEtrkskwetuXNWYvDoydo
tlNjVpxWtW3x0RgOqLtDiVua/x4l399Xcd6ndLWU2OlUMQdC51aPG9+HihiV0G5WKqToO7PArDOV
EUyK4ktWT362dKm72tzgsQeiFWEGCQHm37w60Hh2L0mI+y04Zw/39X+lRAeOrG5xxqKA799RuQnq
ncd/YpPhHthHTHsGsd6SJ1EoEuGoYXatBDhT6oYzriBtg2eKbijCaxENBzY6vIPhwMqvIF/9uAhZ
7hJVGv0eWVUO9EQCpfSvZHxAA6xGaZzI3rnb9xKlYzEBvPEmdZjoj/KszfaRj53O92ei/Tay6Qih
EpAK7NCdIhZS+5VX7GCwoamNGcOGCyzRDG0Qn9uP2fC5CcfPaQ2Y8Sc3ve+4e/CJFZ3Y1XEZWNcl
CP+9Hra1+yjoNpCn3909G/0tr5axIHwbu16cY96rag+uyMvRqWaaySRn6gJnptvTZr/NO5ffury8
ATI/qZxxPe4hPEcrTc9R82kQTcW4YvJYnW3lIePDFL6JZbXygZUxcNU+fIdqU5gm3I1mwt2nrEY3
6YvjFmTit+mwrvWoSGIzyXVnyhImGYZR/zLRXLd80AYrRY18gmhT3nlksPy8PXlDW1U64UZ3E544
UUXHEkine21O90muxW0W5xZ1gVtYl0w39tQ/94s4Jw2WSCvDEhK05YHwj64xgBhZlSDsNpqx1Uqj
FkyxobC56x8UvBEiprWOBDqil0oGs2yFlj9dXnsgCLTaUkLBxXR3Niq9/9hdiOBM29clBHpV/+rd
49ox2jb+x4BQNktuauGObYriSuh/kLcfmImTUMzmq1uXV1hDut6C8U+60c+cD9UnyEe5KVQFNIJD
Vfm9MP4q5k8ihHzf8tZbfLp8KFQky8lq6t8Un4Cq4nC8ZnGjAdQ18BhG/15mYppPfIPuOazuKVCD
FMaCqXbKh+/lRKbJwacNmdJAm4PteK9EYqfydn6V35afDv/0r0yB/pG9fHzcgR7gaC0Q7IsobW9V
m8aLz7PF/QfYMaEEGfH9Uj7MazdsMNZmY9vWRCPR1HffA3VYYFJJP+hzmAHugYcfHXWMnJtUUKPU
m6hZSIzu6B64DFX+MdmEKdt6c4B0EvtpmulX9BmLEtBtnTR2TOaefUENKbinD++xAZ+9aAT6Xq1G
ZEXJ/QgwPHswu0gkmzPMLuEl8zYpmAAsWys/3VAFTLAJit1e0JjHyyK117vDQePcn2A3x4uGPLbp
Vh0NKqZkCaZ5tXXvlfelo4Qy7qcxck1zV7eSyEnXjUt3u3zFi80UTKzk5DGA8CQvg9vrAhRJWLDF
w3vS68P4f17o73wk8YozM+ZPYHa1u24ib6ngpsXDzi234jrmVgzrNvFE8VNCTfUXCc77fkhZa8Aa
e1M1km4y9N1/OqJsmgFb5bPeFBpskkySTTPxgY8xKyXhx4q4f5dIo80YebpOOwupH6KFDH5Sty82
33mNJG4xsyXauseLU8iwvAvkY9+jYBAmgDI7wo6q/uxD0PUuIal77p3voaH9xvWkjkS6Sz61wI3d
iY/rZmZDmga2gewurXNBxgEySwVFnWabFfMFtdgsbo6Xr5SjynSh2ijIE96jicolw1taPDKtSi/U
xh0Zx6oJn3fO6+gL9iSFt0rB+H+N6ZDCK0Vkq8IQ2CdLBA26lDqzJiQZlAYxNG52RQigdm2DJcEK
BY/wBFdkaM84PdcPLYFH8eETR2n/pQcWf7EyoJEVCFmzxfEewLX1zLWmbDvhrKgRXtFSlFXtjbi1
4tjCdGwuuwTofrCa4mZbz9qP3l2h85tYnCenyi5uLwPAyCFnK6OqxIn29ZBLa31Fh38tFjjHH4Gl
0pyB/Sgp64mzZvdtdCr5eB6K+YRDHD2eyIiePeC1+KkTBIk8aRHiBsQRKghf+TglXDf1Y/+yt2u2
kA+o2vEQVLQ9sRwfVsSS6SR1Z32Kdx0tiX7jFJAniHL1XQRfbRm7aSnfT6KvaOuAv6G1tIDcOdtw
8reX2Ig2qSMldmQUPv4PaxCewnWkQ9mWjDRoaAaToI4A977PYfuZBUZuUJxFmOjBK5uU1m4X3pWo
nDieWy8IRdfKpN3oU9K/oTyVMnL46p5KhXJxm/vz9zzBmeHW0J5KxzyGgWXstBskFTppoKTpc+Gx
WFNVAqpJXO+jqCh6KmKvZxSR2SaPKPP0ktPtPasVyoKW5uXul7UW0uxqy1OuOUHyjT9sQwgGG31O
iGpfCZirmrzXdU/w990yhGWyxkh9W5z7hNQ8n74liZSNZtaocRuR9Z60Cd9v32iqMGu2ichgAK3/
0+XUnzEh2ADzxrx8WS4adgUOrQ93NC6lg02GQHXeAqRI1WETK0hjk1mnaKrI2+dqunvfo7dhAx58
qrxoVp1KRtZvIch1EzZIUm8JPL8wqnp/dm6H3NNULV0b7URgm6XeIA4qvzciZYdl7KCYANt3n0qw
mgyRliO7llXxYPqOrHkWCl0l9KjOfDIOhohVaDOqzywIkP3xmOFB0mw1olxtov0x9i89DHVUi/eJ
azcGtkgQnBEeyog/GnUlUfm3hlUUhyxu+d4uO2+2L9ydZoTYCRkeoG4Ho+GUTPIq6WhpJiQI2w5E
GWKV5aVNges3yVq4Pa4Hp3XmrtYzFP3S8hRYbAwnU69nwic0wqfwNhOdlo522z4xeYCmcJTXOM9Y
PY6uhnioqR0tPwh/sElI9UMMQpAXAqTaXf0V2LrX3F9Z6HMgQW+roJjDt6jVHR/pFI8/pJZx1srN
0scLOL+lq1JQRDEsWXon7OLsD2wrg2jrXp6cvD9oQ1X7mgyn8gQYKilnE537BbLoc3ToEgqoU8d9
nrKgkrojtrzSGr6Le6FlWf+bxiLH0AibxzGljWAl8HO7ai9PTL0rnBjE1r7SDNsDwn3FEoscoi8C
9AeMst505xKZpr+UsNS4hnCyqrgSp2LbO4NzfMwRzvKRSjGG79cUxmWKT9RrobFWK6nNT/4G2sL1
bZAfWOO2A20UFZi9pv1QqEwWCF84IlzhtitzMalhEGwoN6KLdPCelPHekqtIetlom1Ek4gqop/rc
XeRjZcH/gNtt7YciJOuQsA5Uv5iVhwYi7wkusnUpVLIal+qdPYOGwlGbHlk7n6Y9S1ochqc32FjP
jYk5l31/yIXnqTSAp6csd/0i7lozbwkP4pbZ/09u3/So5JzwJDWiYX+AdLmNu58HaVppqVImOSIE
Qc7vsSlQw9leATz3Za+Rr/y28b+3a44FBJJocT9UryLTCTg4Leo6OUIOKTKAejtECV5ChcwtC4Aa
COF/8EZUY8wTddlULoNBuAH81tr5Fji+ITGhbBv+plwacK7uYpDGtkk4demV42EKqsgaNj7QODuC
jRIu7BPvw1Paf1hNfkeoEo/fRdTDqQrIP5Mv9yQhl4dG3ZfaiAyzCU/gf2+orzHXV7udIVm8HjuM
Avz/tGuVUb1xM2dsTZbeA1nAgWFyfsYMaQFH8WTnwvxqpiMOEDkrNig9EQeR9W67Ll15wAH2slR9
X+CtzgnTyKUCt4BtOlgzIGLDgc+iyKtZsA/DXut0kxl3dQZZ1tQFkpAMoWXwRlHnmuFsdX8G7Vmq
2QJUxsGLpGa2tCGGKhCcBPh0YFHGeClWxchh50+vbVOCyRtOnm8cr1iM6xjDQPTI8ytrW65SE6l3
KTH6E2hncoIqZWEH9I073/e+lfEwmpNIqBHqZ/Bm9p7F6LPx3uFa+ATcqO/qgF78a5GfkPBNg3rA
EX5QslA1yOOt74zlw1UYj1xZFfCqi74wYGPnOKde9SJ2yiLf9qRH/26WESROkLNTNdVn0Z6GiteC
0tzA2IIzvMLKdz/yJ3ZCpuadYW0+6gm4ZOvaXTqi/GPIvc8EluYk/pRLjN10PRtLyyStzRlaCWgl
0YL2D8xLuSAWPmeM2tXIA26WWRL4N85mg8rOr1m0JelR80Ji3nBMxGJSTl1Hq8oPm7o4NiAYTjEE
9QXcl6Tr5nTR81h2qHjfFesepVmcOoPml1Tgxs+OpqNvY7DWElRFwXmMnSySNsftn74xcfbvzMHH
nt4fMElOkF5yLZb4+/OlJH9R7xOolW0Biq0KzTUrc4C9tAPGOI/12feaBYXMpcGYnAc3u9MqzMm6
FNf6COFHhlWwxmU0Rk25MO7DIjHMS0ij1LC7QA8v3C53q+7X1V7ifictrtzh8kOx+7cQuN4ao0vb
ZQQgvlJgJUN6sHn0xYgBOrVSHG8iTu2r2rolhJQAjXv2Fixu/VMmPS8lWcktReVMXK4eT8s5sgz6
OO0QeB43Z1dg2bHXXZF83bQB16wJJzRuEzwZLpTqFLWPtyPfgA0PnhXe3lLGe7RyFSG3af2RLrGg
lxdvA80l3vRctfn7XRjGKGqOLn5DtnUYj8ETlJKIWQmC+m0tfLBX9bRUqwrezUKTpgz1haXauXHW
YGqACaeFo2ECzUnfRT9ACAKJQGweNVYeweLLeRNWEnO/6K2mcZbrp8kmsT+B4txze17EoSRiFIN+
l4Zo8rExtqNghVWbmOJwUf1OVKa9fOq7s6lBN79pWNNlQQUJsLDYwtdElmIaEaD8w6ZO4WXklSLw
So81/SecoWFjlv+KkgffmbB+9AaeR85Ej6hizp6UbyNBpFIMllKBwhAoou6DNyuz356rRMZRvMfg
Ol/GIzmV6a1LUKkG+Sb0cmq5OgAVuPHnHnd3HolHrVqTcsL914ESwwBPJaA94gCs2LY2CnzQ0kI/
ufdJk3cEHEXe8k5t6YWvCB0hkMZTEsR5kb+lM9PKvD0B1KbI1Ra5G6lhM8VrPK7p+fR/zKTgnYKI
IAW44glg5T6EjGJ8b0EssNuqTaVoNkH+NU7LrTbZQ1ZgXH8hTRT17qEEwnpYQlcNhqplOfD0MANw
wUShm1bVddORNJqs8EO2N66euWe3a1z2Uu6ilUC3/5Od7gCaZtJtqZNMy+QBeJ2DEvaDGVvqtzmH
Y3lgpM+2vV0pJWHAcJTrXbSlrBfnezlKDdAUTO46dor3OouUobPb88Yv6ttdGoiFSDeLd9jEyBIX
Ox2CLturjrnmz8c7lKnsacgyZ4QG8MXW2/xuWIZ/tMhX9SSpUVxMNtkfunr5zLahvDwDSeF6vLAx
hhrCFA8Uhs2NmDT9okz5Bt3elKRCtT4PhGYSVCdtLpAazUKTsLyv1pWb+Y+cNyhhE640IrKsPc3z
fy/3QiKlRkdISOGOVjJwzSTcNCWgIRHzVxa0V4YNl+8FlaPKv9uOFg4z0rlJyGmj8Q7jE3muHons
HL6OyzDx4TPpkwaupP/F5IKsc1zn8CvGFJke1lZcvEALizgeePfFGzNbUp8N6rQOhOLkdEtJqJMq
y4mUQpgOO7//78cxpbHfS8ZroOJF5+oFnBbcbNsLxzP8cUX76AcqxP1KNKbWs1eVenJg0jdkkmJC
yfGulZyuUiVeoF5g+Qb9nBeK73XrQxHZcvp1k2Fh97QRpdF02U3pX+lwRSHSvIasn489S1SHVJ+1
OTzbre+II8/bfKBpKOSYTbt7S6uJroAi+AQXFs5RsVRFDv06iWSW/L5bvL9Y7P7Ntqlb+22Y/LeH
Ryw77EVkWw2fANcZxPeU2eYh99zdG3Sm6ioIA93qKyTd3YapHjAQn8vQCC9ZxrtwWNgmvxaDNSSJ
ks0HOfj9mMrVd7XB692qYcF+UyTh4uTMy8jp++MQbDh1qrbBklO+0SOxXI1lQyD1UPX/ltkfVHoL
HzmT/yauSICThT7so9Y27BBVNQY81jn3mI4r2gervf7meTis8DWJSglv4pHhIW0tfN8JzPjpb8i9
5T/YecW3z/9Kix4O45cKeHTIaocJE4h3ZGZQytd2uu1pA4GosDOuoNPXwVNphv4yFbKwh0qV8hFb
X7k9Jzrq0B9k4BnKwcY9T4XNeTz1CkM8MalphSMnWGDWTUvLNkxaNXIKxO67gKtPbCzNIMp8Zs7+
2FevQuZf7KQPfVazg7rCD1aAiEcgy9R1qO5epAX1z8fIwSqKoUg1MuPDE+cvLPsPd8ABJqX8FGXJ
Jiel+hi+Z1XF5udgDqJnyI7ESYHP2B/I73R9hBtiAOrb4slUvPlbk6OPbZzvNSxItz0yTwGJa4MY
Ije6lvKcCvv024XcLhNJ3g9RDl0VXmfH7/CA4VI5bGWpaJ722EbuStrd65mNGes4Z/J8tRe7+kSS
39zvv+gTCr2MEAQYIBJAT5CTdzbIdYXKJ2rWUWfKXh0eQq4UnHJh8LVK+0UOQxms5afZumnGULXa
n82Br1fiKqTrGic41IvnsE6fHr1FnkNx5Yq8ajNu5brnmkwq0rb/RlpUmI14hKt0jGMEvzsgiumx
jxq1jpPU2aHUypIO4aXYcLVzt93Fwy6av6rykXREg1WN0q42Gle6khQORgH4WufH/TvXLkS3Ote+
rZn71PrQwBUR2jDoHd7fOyqanLAvGK4X4NdVBGu89hlFDkzYPhczH7WkssStSIxe2SxpmqpEmfhG
HhE6Hdc/8m6Zy5Un53cb8Mlbb4AvDCJMQHpxjbS6YcMEtwc9lENUMP7s2weiUmllRdb+F/zUkAxJ
t2FmWSX0wQcfqR9rrSDGTTnem4G0w29p7Z2+yKCoH29CTv1ZQ3XAmv12SjFeiRBcmCE4VUPLj1+2
LdwoNcOkbalPOhLx9gwC1b3YU8gZjhyTtQtkWBPXtwxywaesYX1aYXetfpwC6tB9sAEMYxJwzWiQ
BE4LLNsbACAK9b99jeoRcYli4f2TbqaGFrT7P9kKR3Rmil8owPRZ8eWH5FBlh4XPnZrpc3fBvAQt
qhVW/W9xYIyj8naUe2lmlOn+NfUVQIRucKKc2VRyjYO9gLUiDA1UmWePwkcLjI+78k/oeWVOkfaT
UzF2yGbx/Pgok+f2Bd9BEmmIVVY7r6LujsAYavEaI/Ahn4kZKCY+pHPqus8fs/q+AxpybJo+Wgxp
q2UhqSMdj/BWo8fq+KhIa2rIGfCgzEjH+q/XKQQQPkt0Gm5lo9a2ZMuDa90uVZ8FJWIfwyebp7RU
9YEPS3xFPRLscd2wSUkDbedUGtaeKoss9mLOrzv7kxK6O7qvKeg6epZsCbediZQ2oyshbtgdFy5p
+1yJgwqSjeGDs6cvV2Zq6QnyXc8Z/72uPzvDUbmRuY+yBCBcrorDzJBbQgiQSkjrjslNQhYv7/13
1ovyfuvpVSNd/oiGyw4bpby30Et/c8qgAtW6uG5bl0zbHc94TS2DkBGv4WPlTKKBgVkK/jP7IMwY
luBXyU9wOgB6QBx6QhEvR+P/Pzgtl6Sbs01CcTMtC/uPE/fBBSmHlFfZhoPyRbqE5Cfi+N17v7of
d+6aU8DezEnALtgsuOMo8mbP9P76Yov9310xGyMmio8ExD5pwFTM37jZNwlqfSU1CfPCaCv4Xh2p
zYaL7WrcKIU9NjLRzLbQphu/c9ZudoK5sbjj9Emfr0qiPzWrTnIoKvK8qbYjNHd8BWBGbbtM6r8R
J4R2rgEliv+nCvmZvgw9rJWIbOIVTnjpOyvU4VWw8lTqnKGBwH7d/4pMlLM6QMM3hmwjxhR9Uii7
yxRaqiECBeqdAiuVb2Y7EAYTgp9IdMVjmvexYZt26PGe7zSnBumlUrTQfaum8cUaK4NehdvPWmXh
/V6eUpFGjTX+t6CGgm/xKUowuxxy3EmMGg/fFrvNnmAT+TBH4IAr6ooxC91pZt2+iFWoAY8sPnCB
2KPthJZ8jFEaAX6tfS/fvAqkpgU5tHKGthRG7Mk1UwGy41b2PS8XEXxQapUXtFwmFYDN+BpD/KQO
I9wvuaUqaUo3uadPIB4lfVdkB6Zm/VckOAqqEydsUeOs3kexYNE/kEBAiMv1i2SU+zbn/P/7AcCC
fwYGa4N9gbwvuDneJBMHB0NqnSEL6oysVKJWEJfw+eIXnZ4whk5eKxAn42/y/Kw3A4azMYlo9rTc
PYqeZO+ZYM2Mw4xDm3LaaT5hwnksJXCfbbHuVTs+7FY4wySQv2pond7shqncIoUco7dNRs30fpsJ
p7Pf2MV0BMmDJeqt5cZuQJQszyDC8em+keAYxqG32PgaKsTgBhAudt+d7PDlQMRhOJRy16H+Pj8e
gc/dBJipeIrFFdkZ1YOL0/LhJmXxW4KTU6QPk5/sWxQ3JVayaR7KQ/vURGBqhmYE0tILC03rcTA7
Jiq7isWXt/hPCQ+AtFToIYB0DTOR26cGl7ZZIfngFTfa59wmm3vBfqPtUj3i+Q0cb4Zfrm+xOK5L
1xcSm5aQo11LiUUzeXUzadKIDjY+RiaSeMMjy/kzRtvuScQEpqal/d5U+w/bk4urZjpnbNbiJDLI
W2UbA8Dfk8nSXKxy4PhRHvxBVnMB19TRzxPWfTeoMP6syskJUR6E6tUJjpFSUj6QC245GMmVPtXo
21a+xr5eMz/8Ose1eZsi3ylZB4B5h3dYg10dAufMztDBue3be42D/JX+4jlOWAQFtG5AqlTSIu53
86dt1r8JSD1AJTP9qp2NvvlUMCDhmgqhSEty+HXBHFXRpDYj8UAoWFVXs2T6cvZFZPZfGPzQX/q+
iJXJJB3gc1MHGGYbgz3dNjdn1XvEjdSJikEccI2SEd9xyoZAXWNAs22ZAf46NB4EBH9myhi5Wyt+
n89CcwLVNE/iD0LeDZ8N2lZoCv6lOR4gILoq5qa0wAU6wD/SkWWDJOQFSCTi5JV6z0vuwdJckSSq
Qr1zwJdXuyd7DYwo5OjCi8hg751vP5zNSz/97Sd1qn2Sxxhy9tO3GCrqVpPtKdWWN9/kZ+raq3T5
1USTn8NZ5kCNSenVE9/UVOCd/N27lqdYOX1jdoqTPbju2rHyWnlewTZc6O7JOArgsOL3mAmj0zlN
U1l4izF9/qjnh+o+FRNv5xrigbnxkKMNZ5TBDPYe7BokYT5LGovRrzT4srWIHL2kr3JSFFED3oAL
B+xVEOIIHCmIGBFwQItFSTcfDckijJwL7kmd3ZnYZqZO8xDNkJDQBv/faJp0nxi24IRGTWXu52vd
yLAQzcVbKMJ+E1z0EIp9uC7UjAEM4roIPQkkS6+M1CuP7NXEG/fMuM/SqaxpvrWe88N849s5U5AT
4dOt2ajTlRCSKym7nHtaf8zVCqwawC2gt1fFYBfyAjvJV2cu/mk3VfTVbLyT43gXtVz/UCy7Idb8
nbFC1SNVle2pTk2s2VFJtz/4r2AAkIebbExEsBd3G4hXRl76jwSf+7CbxO3NRNL1tQQdsEz3rB9Y
RGKeypKlfMWsZVDxDnQz+NkZctwIUaJKDrQ2HMp041zXQBdp/7MUSXRpPd9gSnsUd+3zNS1zm0Ff
wJZHPbXP+X2/wrmYwdir4pdPMrnniLAqyyNxq00ccNI6WmhR+GKWY7eHchaRQkFjynUA1c8ZHewp
R0pzs2a0E0XMZNOCv2/fBOfROD6+aC29gMyIKabhZoG3ENyiO/jYp3DsCM9iTVKMTynkA4v/NpN6
figz0def6HSlVihWIiB96QskyEBEcgG2kUxr0dZXJ5i1jdqIXOwcvNvyJOH0TJIbFxTCofQf0MHf
EzRpRSUhkM6f7WeBnKVql+QUSI81t6GtunvvE9Y/AC1doD2j9JPX7vIqzcqe0fobnaaOieP8yH2d
of2ViPLXkh6gK30HLLqXr9MZZO6HQ6xT7cP6uel50lG6swhUjEuolLy2Vir9qsKkA/RfqDgQkSh4
IcDDY84yI1a4PbQsZIl5ajVulTLC7gQavG1PLjEjQzDa344+GCQiYYFWW4iEM00bw+kjDYQ4L0fq
hZYVP+ogPqRgbeDpy2hdzXG3y6tC27tdx4UqXCKLLItCp8Uxv8Iscj0fjXegtIXq8+1WeEfSy2yH
BlcD0CIOP+lPHTmgeRWBQqed4B21BPFAIMnBfMQZ33eXniZi076rdhnXFWEzyCN3TBh4vFBtYoAq
trRWhMhNzh1ddYXty7F5AZRWNNfDYh2F9mUZ2wd0mq+cUCVNDUkDe0GUGYC2W1rBH70xx1+0Te2/
m0mjWPBnZU18YjtgAcR4VksfqTgw8z6yFLJCSR/ZoEluPMegW/X8UxM2Woa5rpHuL91SfzVnMYzs
ulNIfNHnsGNgfSxzpUkyniWBcM6LlzygsPFnYjPt7Pi5IDSmpkG1gtorqE+/EvUExmcYHKCvtUEM
RBTo/oC32mXwISLH85UXZ3WZ/rGNvM9gvff/nX6j0oHdLqEpOEtovbUEb/Ai8MWy6wTocN8uVwh9
3Am2q6VJE7StqTDbUc3AnlobJzgwyUXUu3u7pfa8Rl+dwLcg4SVYw7ll5aX/90Ve3iN4tTSP/fr4
lxtwZJm/uI1QvBX6njLgakEuSMhBBDSpIey9QKHk32NSJFlMxdN2D8CiLZbo/cxm1TRkX4LjENOH
wrkEnK1rlAj7H3CxweVv61hbrk5wMq5T4Xm4eg+jp7fZtjdhgS8t489yMJY6D5muVjdU4RBQCvGD
/5Y4nlJAijxldkTqs7LuiT619Aa9e6kGOkGSGt45s+S0NnGVNXG8ra7aI1pzY0zPLdsrroE5l7xd
X4U4YPogfWwpEf15bCK4BceiKD+QpVq9U9OxoIzmkVJ5LDuEyRmkt71/Gc8z1D4RpFgACdy3gMuy
9F2YPFYvp3Rzh5fWyRjy0bH9J9CMAH7Jh1NJVIdNDWXNSW5U7FNzq989UXlwrzXCqSDXmlyD0UFd
ZKPPMVwaSnKydjVmz4sfKp7HqnLxqhXZyw7DibLq3MrE3Xv1losG9jUqiJCZurXg2GgBhO95k+tQ
hRW0XoLDjW8AUzFbXa5bCy7DpDv33VcEr/asVq2RyWEe/rLYZ5Ef+uhRVFuahYWoGMbvLtPYQ9D3
L2xhSbICwW9OIVBxWHWBAzLk6S3JWtiTlvGXt9pY8gLNHAh/BKQ+s2AiZZPPfVwy32s8uEtE9e4/
qA3RsFYpL6GVHJV460gBQFqplAg3dFzVK4o0oxYIeiBeJc6a6xDzcRA/WnAMv6SmWA6S3nPQ1LuP
52/s3SSMX4bkFlNtRTkEAdMAoeiM4JN4grRBg9EQgrqW3DZelQbZNwUk0+M7flUM0HrMxMOhymiD
eIXTaXJnXBbyXFiIKMvSx1BGyQm9PH9wM8spC3ELRSFHyv3tx+pAEz5tVjpnldpwBkIVjiVmrXdR
y6d3gaSk3h5zqLjar9ijOXs0EpPhsvwTeAkWg4hL20HXcnYpTuxQEU9TscrHMNJkcU0ba5RNbG+F
I+TBM4298YFo0pRQxHgOZ4Xu54rqd8N56ePTsXKOUpOaE3w8Va/ZaW/o1W+HtWHGeIkr9T7ruZpN
BZj6cyZWY6Ss+HN4dSCPCMqPKGOOnBtIfQ1r/CLD9h8ehe9Xjb2nN0Zpi6604y5JIqSHF/2ADLbz
LLuXo9kZqG4QILJb464Un+zzY8ID6JFjIJeXxOx1Y/ClVNB9k5+pepxvm6cSwImxs4sMjeDrAwnd
dpR9CkCN04yvLOp/so8kg89ZrWyglbBS8TrXclIIOrUuD+TdqhQ9Oh8n2oYux1dpMWRg+G+nuj7T
ClaV9zv9pwU+nvoIVW20Sq5IaXbBrh7iK/H7qF9tMzj0CwVdyQZmU0wmU84vczSck7QNsOWWuCEE
0rBsmQVnEA8Wux6pK3kZFFsQpDkeTaJuQohpR96x1DR/PotwDqsudkzPL7poNxu0Ro7X+oK1hwe7
BXBa4wxlp4YwJ576o53Eb/NCZBmPJMjuXkOpj7C4fmQ8fARcSYA9AO7CxkTNIvkBwBXuWtELCu5b
cyQyAEUpc8zA/mx9hvsyQhiTbLGMWxyzCIeY+kK3HBiv1VnTmXsGlqOTnr1qPKjLVR+SvodQ1Aae
wsfXDjQaZaUyKU2BZ8ozRsbiAuijDvQ+XWG21+bjG5WXvwPOCmBoV7BjWEBPltrlW/0TEgiBM8lW
CSMtHPUyWILnBSPLDqL/TIb4a/YUv9LBElWsh57qmaKFM4r4IF7rfZ1fxWNTlm7WS5v6qahiX942
CMqwzeC2bugvNQoOTOKDCVm8B0mPLSlp9VNNSRpVDca7EwtxgqDUoJMeRGwwJKzGYnh+451+rVYC
FOaq68yIw4rbrqJOFMPTMvZzLJVtG8OFczGgiGvvjhbvzhF0w6Y0jLxtzgCz2DvfvTC1sSX0CFH1
Rk0Znx/ivaxrlqgXBfu6J8l0bK8/8hgV6DJzak/H1UTO30U8d9h8uXRlwHfC7Lp3GYf9MfXcNv2h
MbBMyyU06aela/DEmXMN8m5ZnsYfRHwV0pQ7/1oJlHa0oHXGSaDESH/zlXFG957/48p6INKHDnVO
AsPYqFteP1sCk7obFG8lL9SJvqyqktHbv+N5cj1pnmm3eNic+5XdtASOfVqrDflWLI06dTdDiRiB
epYsksSGxQgV+NXjYZm3UQ0tSLFUTRttifVXGZGR2PDQp+WGLJPDAc5drxiXCuPTWuwoRLAV84eV
pu06O5xU/sr+Me3n3umNDaHf0AV16S+Pf2Q+IMM8lgc/sIlK9QXyMVEpIf5suNZB9/gC40Qmcfbu
AnUD3bJDyoOykaWKU/iOiPG+2dFDKEP58WRONNKl7NLobPfalTods55PTrHh+ix2pCgQvtkFuM1R
9+UZuUWx6OiWD2sUg/muTqxtzL6ihKBsvSd135ApuPESVgtAE+kqOyw6rjlItCLlCyUC9k0jd7sS
sLVpfGrt7B41iQg0e0ULAczSqc+wPkrKltatWVjj5f8jWm+fZqJXYRsMiGilzsFS8lK5Qrf5gMrb
6XHnqigUNsrpghUMuBHI0DyHISNHO9s/LMLMHe/XCRVaypq+zuGoDlo6NxtELcHUIgG2dqgIXwHu
PqujWWDJf8tuKSNsO5pKbzq1ziGUQmToGzxoLT+2e6NASxJ7VcmBmf+KfJRAgtBwxvAqEy5Tcu60
n75pL8LjxqYaWLLNV2G++CBoNjUFQDMvoZyUu3ibxxqhnZj3RR5lSRxJn57eZqv/3+x6fmCibV23
Bn6higkMDggsl7NVRIQ+L8QH/Z0gVBUMU7ARs8USZUvjK7YqxkHG8BnUZCLq74/lN4YAVUYoRiVw
HcV9t4sbpTRWYM7LQ24X7OG3QFmpmH93MD0BYEVvgJD5F5vSvhSQ+iGHlkCx621xxbVa0Ha5kGeM
XT4A8qTPJFXcaHwUBnRsXTvrHngArBSL2YeJGDy/DzFF0ikDCY+09HMG05w0pO8sGo2BdjNoWwEC
8ovAyZDGFAkE0fL4prALlB5f2ve2KSErR6LodDnaxjSCnoHe05tATEed5jL52bAz8/ZgzRPBrNm9
CRKG01vxdWtJcyV6SmqWZdfvEDxwBXjniXsUmiYE5Qit+UEnJcCMnL2U32gutGf8zYjtcA6/3QPh
NwEcpkx/eYIxvAvpe2bJxRPG7wlJjk16D12m+0bor6eySuCFay7sQMLo1snYEE/4YH07wrdu96hO
Gh3yESIFHtXp6h9RM+VmUIpokjF/CrNy2b2yPI8BB7iaPmnswIOOw4LSSpklXJTYXU3idUeo34fm
jBtyNzC6BNFCHifgIyL/RaU7xv2jea18U3zVLdJ5bx1kEwOGXSCWe3UxPFOCVUhCvUw/M/pCQTUq
dIF+bGOjvWRQtYDpi13ppbmRBEd6t8eNqwZni/sOL16AQIsYTRAIdy8bI4BIsG2vmvERapVtLYt7
Ax6awI0rMiRJ6XEvhURaM9T5WDmK9WUIsteQ0YaTRAdXV/dbCXZi3HxOS2HvrXCBEJ6XfvCllD8/
8UUTg6v8UDQIHGmiRWGkOfac6VheWTIGC9pAyFFcowQuczvQbIglJhYFSHI1jh/yWZOVRfwln4o7
Rkcqsvz54B5MSCsYz7JUwGsdb9HMikjoWJrUJ9HZ+av/P86Rf5O5lai6bSUZCoVAxC9UIvSi2LsM
GSnDulOMvErUzTIe9ng6byjWvLB/prgt1YT5IHtvLlDc5KG4TwTXPgCvcrydZ0E/XRH6fmKmVdSx
hYEZr89N3JkgRjsHHUhrYE9Vg+GWIBM3qkeMG9bg4wW3zY/+G/l7Xu21YvrCWKLOntNkdhOq7dWf
7Q7RLAbBH5Yw4mUGH/2ZjdUDeyAXdr+QdIpNozrPvAd0ptY6NmwzkO7+5EINDX8n9+YtyqmMYKue
IJIfaztEfhAdeepJzggvDnliZVdmQOH1666rBkx4hkjU0lxvJ87pW8YWvmb7MGChLiELgrQGDOJW
XKeoJZbSCq+lMgls0gV/Iaq3wu0vd6pNGStTVWXbDA2Ph32Ow6LujDG5h/kKLG9b+eIWu2q+tMc7
shMlQk7trsghwsnymZ2tSJ+OwnMLHA9FyP0rQhYmlI59XwskKHUC7pGY7uC3ISAdiOl3BKPL0SHh
mcs7HpeQ034DElaTexC4+OfvTjWzeYliNmnZTpL+VJV7QaBuLwhtdyq94cD44+j/WTM7iKq3uTBP
iNlSRdbJTDCZN7Ki/t8JMjLoMLzJBeOTsIU8MWCKuhmLPui4qRflPiNYDmHXlQDFlGl9DQDNCIYA
etDEfBR9XebKSF9u5Il/vF9mk5ObYr4t4fr0wgZYqZubzR1orn9Z8W2v1MFSdYlixEcPNgKWkzP6
CIW4yzucn8Xx8Bj+V9d1giGv8mwV3PWVfvSyTbUpHOla3JFovyw0gWhxVjc5F1umGooUXMT2Cvx+
sSuwe5Yuu4TO9fD+bIkS7lklOpPoUdUgOxt4kUExD9pgGPHx03DxRz0E5LJFSA/bxe5tUjUUIulr
pqelJek9xIrStwM9P6HHxLYAbP54r+k7jB23wi0oqLA8YSLXzzlRDO3Q+aN2LnaO8HJlIl7XPgdU
hrK/BYNtAVohOOqS3GUPOuxCe6aPQorBrk+oEzh6r31NQqZDVPSNBTs3A09hTEfna5RNa3Ep/3TQ
OyGRMtqb9I9QcldNoX92WKZmCLPj+wKM1jDWTXDTAR5S5VAT92u8AG4OS46NXX6tda9KzcmHpYBm
CVqdjKFaCqRHOinlqYLDfW2fXVKeE/D2hvoEyJRhSN0fxoWuOGC+SfBUQAxBXvueE88RcaLdPZzc
yypSRXRfn+qCNuf0egEhWopmBKxclg4CMPOiPunw8T7vjbxrfBlzq9s/JmrXaCn5ISRtn2JGVlc3
szxS0wD7xcEDfJfThKRctpEGlT0OngX+xIh/7JS0PQ8kyVFsLGqXf84WGADEpTXlfK8Q+LDjuavI
+l/wzYWQ262eE1oAsnKSfWX6LVA2O3ywx/nOsH/Ml9AJpYu9A1zOz8n6Cda+fuHCFcmf8CAkBtji
q68p/uReJB5Qaj3073Y7bIhgiP2vJX798OTAyRH6nLk0n7sjpqbaN93wQYhXxILEwWlEsuZfZCse
rIWtl74wFBXVbOHs4mO36GYLKDarXxAB1hbTD1KxwsW4rlkdlghDY/J2Gst5CDLDSThRbn218KLh
vbnDRSHUizdrCLY+qTd3yjCH3aMA9YNG3yjWBbnwDNGUCk6VWkNXmXQ+tPOU375taVOdL+rzdlZ1
xil+ydoAJYgjaCglcdpmzhb44uTEYyfOD1PjDrpZFF+VtCflSj529sr35wulDBEI5cJPS0s5eOAe
GdEKyYoJ6QVrNPyaXt4Q20fDutvfZh3AXYwMKaAFQwX3rf7zGcN/E5Bn3nekgSgerRJLYK7PYd9u
zzgqP72T65lUrY5QWyNbzOIh/xmrIAGO6MosKi5PJAUno14yiVXoJJepximlXi8LLyTjCOii67dn
hgZgedRTu4EZiyFfppJbssVGRH8WSyy4NIrDaupCEUBwGPnKklwMBurHLmsxpdRufT6NLCOVf69C
YQJDGsfUHD3nfEyMYQWYp0UnA7kF/4jdX/ut/AhIbI1Yet5KXm4CO0z6rRNtpDzAo0S0uqiwC9TZ
4tTWxWSl3mqra0nzUBEtHp3TvtCECqs0N38iOOMnnFWRDH3mqb/0mLW17j5P+74zfCFHX2I2EGf3
XLU+myvvJSPNnxjnW15G37xLjmss0llEube4tskdxlNFxvsy9r9mh9EIkCLGmzk0QDevJ92V2Hhg
SR93y+26/FjJ+kTVxrs4jbjyGYwIsniZjSs8RkY/LruEeOry55umPfxUlVIkbkJ2bilLUcYbvGd6
QaS1eEDcEkHqOr0JisRkzQih7HDxx6xutRnnEn6/PBxISySVqxiXiGbVY3fnktutfCvmQOWlJnnJ
QSpaxix0x2BzAhYyb6GypU+5DOmXH8sosu4lNrHr27xXkR9JJ5KgAy76dnsyLr5ueyhEkNv4kuPz
FwVFqsQTJiqt85L3W9T4cnXXHVNDTezMib+/l5BGd9rolLtDGF3EZzkfoE0CBGcYicVnw0iIALwa
TWHxu7Oq79RYeW/hhRzgyLGNQBF3bg/cYOQbRt70+At5bZyEMHnIEJqJXvlk3e6YL0gXmJilLUNF
QM/MXzqpqauSRaw9h4QBYGzaNo2hW1/jaoKkv4A9hXhYUDNyyDzn1TN8kiCpoT/Ht8SQdA9GoLW0
0rPbdGoFqps0fDcra3tC8B0zmiFmGf2XfvCdlKUW0UBbW8x1+hBz6FMn+wS2Si6cr3EMTC4icZnQ
dNEHW4R2v3LcZwfvPparkuhENy4Iv3LQ9ewxn/zP9ewA93c9DnetABWlza6swm6e8FiDHAcQQyx4
CYw8H0bPODbG0BFNVvUMHDDRiiC6wVw6GxfyhI1oLdluWuxSOsuX5p6x4xPk0W0qEbaSQxyv0Q7h
JJAVJe3lKAio8YBhIqB+cqEuQdw0c43xwluWhm6MnqqlJ+KVaLnFXuP4nh9a2uUwuNT9f5muP+wU
ABqZ5DmMRNlaKnrR4wbnyuZKLyzFcfFKD2+hLFjuDaVQl8X9iYaZe4hd8x/3ikUxkyy1zN1IZM+B
9TPgM4Hs0RQO+CCEF8zrdOWEXcHd6bnFv6r7tVdPTKkkIsm9+kvyU16Px/lZOv/+GNdOkS9yuRfM
mQkozvdfVZFx/IVBz9LKkyhb5yIS5YC1su3Zr+p24/UwTbtxE4+e7q4gXqYkjMhfZ0OmMU5ksAk2
UAw0+8fp7RUCIsihZtN+NML2K8JLoRsQ3hzkjx1i9RTFO3Qj2oFmlel1BM1TsZylVXxLB9rIPB+0
PyfSJsjdwCCWX0HUK2tl1REvQVYdnaTvvRlroAaUU8lcBMAITFvJMIXk+7tkj2cT3ThMVh7G8K6l
uG+OQ/n9iw2GYiONwO1U1tAdBQlwZR2Lhu/URJ7+5ZFtZWIEe+onKoKAkf0sK0nm1HBlVWt6KJew
8ii5LZo58k1oQE8zJNs11F7cUW0y6m94ex4eIMy1PNsatCX1DF4QrPmKy9THPHwhMbJGt3usus4f
i8AFoxXt9ZfoDkv6vUA3dJv4mnxmcRlhCwpQuWc1bRq1KUwkXFe3TCA9GJQxdslOYC1bv1M/6WB3
+jmEK9dvCXUz+sW0aRavvric6dK4wTZv5R1srcSj2Wwmg4bnlzE/ptSWpT+OrUxMmIxyly/bOvOr
nDrzIhsQuLyr3G64M+IuM/yKqnhUA928QGYZRm29oo+cWZpTvEAbebr4/AgMYc+yBWaVxhZQ8gPM
pBylw5545YZEN680utyRQ19VOgY+i/F5B9KvUs/ZW/a1DU8erXxFsaS80fNSfh5GQkX6SCLOQ4VY
F0jcGJl9a9/WtcWjkgk1OLS7PSXTzvgGTT0mSTM8anF+VpmJeOrMLWSCEZ2OyrtvP4540gVynaef
VuThF/zShOJKGx3wnOe/ensc7gHpg5cyPepHQKX+UTYxmgXu3367aR902Ne3H9eVvwqXj7KVqynH
dnjoitnjv0kL2gS3SGKuFutOyi1Y3W5wwqbj0vrB0hT7uTSujKZwl20UIbvRnzi9HVh8cYE8WWfF
D/tMhmID33lRZ11hnxDWqO/u7wl0/WPuqQwNnl9HSB85xWtO5UqtFMjmR4RK+yr1Jdcl+puExvPo
CPVk2zYd+C+cGnl+dHNXaxHetIxoCorMdRFUFqmN37DMUEOkESGt9RqMqtmFfQxrHRTQdqHQTqVm
ABu13u4u0wrPbdNiabpOoC8pdpW9Y7aQtuYBd80c5y3pJoQyTNh5bhLI0ehDSdGMi5AA/dQyihUg
a1mM0luduPs8b4xE+eLhXSzT6H1V+7ZmgRNBiW6Je4dke+4Trnnrt05qFD8Eh/KHwjLoZvLbF8FV
qauCY60f+b7MsFHL0Fes3bPAvFKMqr41M8mn+HXzHGxH8SMEzkyMDDjyO+YvCGUYZOKOZuol8iXk
VzD18f7YCgG0ZjQ/P8vl00Uj7rvBitssZMUwZlJTl9FAa6wTPe+AjcjPZGta4QSSMSIDMN9vDl2w
CF3QXClecSvDdAzqN3ngvguoMSaOTO41SeApZRRM6XctplZnukvjEqDyXqBaJiT10/dMAN3hq/zB
hi2mproWocgt46DVJaSuD1CcYbN/XPwO2/6M3/E1zEn4HkkzNpClDpQUi57PFyUldycB7AOfQJWx
nvB0hktydX7u2qpQwchAT5lvZxM19xYLrYaWmQJkHAbTFsWvgGrHSYQevg5XtyDEFuVVM3tVNgUO
JQMsMeAUztIFEuNOOOg90BTgS/vwL3osFeRnQimT5N7ltyxQa7nURtMHKjjCJVPyC3mi0ltv16A3
ztQi3ZWsMyUiYbMyzZrV9Q76L1+/9PA29SFDkZ4KgD8Ersx5XEytk29NXZVi+bXBVqXvqPBQ/fLw
B0i0YIliyTHHQswaGNlNrL0mSKeOpGWj4xA/y9fNx900Wwyw7/h4F3kJBDouRvpYe9fiJLUrnp1b
ZOEevAHK8AbnH7QdGoAhXFp18w9uHEftGK53NUcfSIV47BviBJMxFOJgqJxOPFlWUOrGtpI7SAxi
oFqW1U9ZRYvRts/8cDTsJw8EUup9F/FdIIQwzFFCKwy7ObMoRuI83yFdyifEhExMLmk3f2e9nKoe
iNfJVDbriD7kkx3U/t0KX6Jgq6C8HJ9taeaHt239DbTR5OWac8LrwcmcLttb3fANHrrHJP3T8c52
qNzabTJol9Kv2KZMeXho/cdyMYiyORA7FzyCYmkNO1e7MKgbkxSLWrlx/d1ArYCIU8Hszg4phlCz
Px/dsRXDNL1fv3to/Dgiuw0kTg9wlKLIep7kz54MBqtZkSqf8eP0jm5TxI/AL/KFqW4ubZqtZu7i
500e8Pb3emvpcTHapX6t+NA6XGNGErofj5k0evkQODxHxwur+4fRDmmXR024nowinNVmbDInf1NE
tPrvx28Lr25Y8k7U0Hbzg1OJlVGE6h/UWTPFlgV6CGZp0SiJEma8/IdXte6WVi3E65hLmhzcyrG0
jKj3VV5MuvcnoQe6Zj2HsnjdvY/kfaqb5Q/TlGY67MagaVy4MqHgXxrWQl3UVvJqeMIze1uOvzI9
kXMI5XrhdSwC5Iiz+yAi1uH4wHjqWhyp1YB0yusqgnMxF6UeNoUcWO4kOUDz5YGyEZmBoqznDOYS
8qY+0E1FmtBkqBH9apySPrn4bFs3Jq9thWoOY6wQtPFdICtAO1fhpqTKLvwvlyJWnuYd05bfobIM
T1a/W9GLB8cYnP/Bbp141TTz81hK2Q4ZXAMIDv/1XQRql6Uxfn3KXvLWqE5BwAW32cZ4Nd+0sklk
dyJq88MFRUf/obTiwenBek+LUBJkc38dp4e2wxDdetYmkSYIBD6vfzulkBrug/s36ioXmbXJgNup
2QwNXIHZmTN62ADQIeXCwrnCNKtnal2L1MAfK5D5zIL/hc9YfKCtofL34U4PkbMnSW8bIW/Dasbs
AFZrrKAn+Y3QEjuYH4yT8OVk1pqVO4tE9OMEwOqg8FNLNjkeSPsKESltE7sC9J2CUjxzK24KDdeF
81YjwGskaH0FuI1MKBsNTVm9sRT/+LALXZMInd5oTRe9fzpDpUekAnvtJ/tBmRleL9L4wxZw/4EQ
UN56X5ACbprtRNZjcqusw1LGxr3qzgGuaJGE0KJPx4+BSIErzm+RYKZtNYojif+GoPkow9vc9RAQ
KCjcCTwHcgmnFGlRw3Kq1N67WoIwFcaTku0BweRSxNnL895zyp5mmrILi16U1/OTi019GoJZkRTw
WIut/z2wWrGvz64hdT0y/8ZI6nMJxWWOu6ACUiYbQVg7R1dHXajj74OSd0bdvSWM0tZ0DelAg8VY
FW0YXPzi+Tl59SIK9jwpaActDi6k87+mWcvkMBxubiX9ufv+FNlKeZbH+W8YFbAtt5x2UAL6adWc
MRhGd4IBe3YRPRW0mrq1MSMN01Yu4UsnEdkXk24gVow7BlsFsKVOAMjxIKJVXrfeCV4q7hj9t3Q0
4Wc/LdxeOlHXhf2PL0ovBW76QvPWXXtxqI42oDAFn5etmJeiCOWXbmc3PbgpLKH+1etBrUiTGx8Z
Hn2aTG+mozKZ/XwLpfNpcfBLwwOKdFVkvUhWSpZRZXFP1qm5G6hIKFdtvvWz04wwxizkObneI7Db
7zfamM2M27lcS3uKwL0Atab6XkyZn/i4OsBtZeWmVQFdVzUmGFTjcdfwuB8uiICRj3RNLZxlz0N3
JW4UMcl68Kh6HWgALnjTJo1DTaErErvu7Xq4E0GyAdnMGZ7IBFDzP0oL5Wy90+pZ6aBsgikJUw8D
HiUDZgVNWAVs9CJmIaaBGW7fxgQmE86V1HqQNCOxbsTjmwvzaBpO7AhMcELM9a6F8TOYlqFWDSmE
LJuk0A8aYN0nqbjHTCwdyT16dbDZ8TiwvnmCBeMMdrKN/09vkuy81z5mpy/w4C21tkPoCNIu9wQT
pB024tq8/mwEIAEMLev7qk7nvHvlg9BxoUGChSscHiuUurQyvu2B90ez7xaqywD5Wmxr0y3RbLXN
ahasmmUsaGI/e2oEZE1C6p2klBvSoIf/Yp0j8OYeL+sKeVR6jZO+exjX5fp513y1dKuVuvBS9SGm
GP9/HQacLXOVeK+qm50+hJlQdfy9uLt5FRYIGfaw65TnfxDB/TJMOJAMjQbNZHORSzNbG9cs8dtE
7XXZc1RzGmo2z6BnlB06eHpkg4/1oLJLytq8oSOxHP5ZgazU9M3X02FzJvqvJ4e5O1vz1hvzc+Yd
oqruqrHEwzkobLLdNCrwFBfMliVMyqu2jPNYYfApvyY6+WgnR4ETrcL8zAR4vEbWyloi8ygLJeT7
I8YmlkutUKKQLytqdmIC1Nmx+UePFbt+LaVVCiCuF/Q8ElBn77F4ViCw1T8i3AzyFtcdilInaWeg
xXV7zOBlSbr5i7fepMbE7oO/ZlY3zYUpZlednYo9kNkalsrjtUkpkXp6IchGLwQ0c17HPfaLRJiY
fRxp5cQow41n2wKGprmd3RDeJc7iyfBi4OgqHmIKK3/oFGMr9UlTjxXOONMPIkCe64bu9qmnXzSv
klcQAm9c9j9JOR2rca6xw0FIuwvCWQltbdLjXxEj6bd7TQn64gXbComv5H75WQmMLt0AmV3jHgwC
76z5lN7re2AeugXmFcI92fiMbNk80FthyGSBbL8mWN/+uyEByeUG5SA02B8XUpzxAi9Cg1PbFE6w
LqcJQjTHZ+Bkta3cqqjU60+hekFJBgaSZ176HvsSISVX5PXennYORQ6taM5Ymtlwpc7FMA10RXaj
q8pAnvqGYU0uH+ywV9+V9b0FRflbl5hFt46yYChKhyXsGcW46ymdFfBB62cRCEM62+pkVQj9r2Dl
KIc/bNDlGha1hgBgIo3VfqJvU8LFkg6mX8J4TP+qA95/I/vvZlGvfF24e7yyIrPS6wKpOtO6E2u4
JbP5QAeDhZYiaMoC/7nQ6NipHJomMSymShcKBwAXTBAvKsl1hMUla/QSOWS4myP85BUPXLdne3jK
mJD3t1l6r9lEvv9mcPQxgSOEHCzgsDZewfmyusvJ9plswlBXl/rtLFx9/mGERlPH52WErTpJdHuf
14oLC8W1Gv2Qnojn89Z56p20Pe8XTVnYAo1yjDBxw/MNXhO2Ln9fig686OEYDpk8h7jr2HZpz77V
c05tsoE6NuWT2uCd8sapKrSSkt71mwu2xxPRoWJShQGXIQBHQWiF9Res3jO8OM8Gj32Z5qRJlYj/
tgaKvy63LBi5opDugvxTFuOBfjQx18wy9s/fw7B3Xsj/1vK2IIBJnM/mI9MjQXXaD0V8Wgn6r30p
g51y2XvtlCjaFUbMJuJ9qhRLRKZ2xKGShXGT3NLw/0eodSU79+ztA4mhHC9dzxkCaapMz4bcYDMg
T38VIxasQOKvaJCdU9kx9EHTZbIfmiMOtXIi+eH7roPhJIY84BVZr0+jhIlca8SEU6XAFCWkuMOC
VFkI6y7qajSo7hF9qzdGguLFI+HVXrvnjzdmkfxFewHJ536IcgXXTwKaL42Y3ynpQr30zHVlJz/D
lYBPsu0BcZG5sfK829fJfnXSNrxGot24+5NXHud2xYtjl5e9YhDdzSx3L6qclW27f6QhI3KyxS6t
Z2q75LMv6oM4E/XYosp6dQ4GS3b3/P2r2eDgNlKf2/98Dr1kgHkSl5lonZZs7cFsZ3XcENEJOIbN
NkPU4CPoH0mM0x+z53U+sCtN6/7dC9X8Ug9aDsOzcHFa8KHlkiN0MgVWkiCBhRkvYf8IHdE664D/
usgMRbZTXn1BEu5y9oREeeT/87t4amuSi118tiJBd5TTGQ+G2iSjuaOtBLDhMFVUz5+IgCcZGv/7
My4OkZQ3L9ra3yW2OvLJgDs/JSLwYps+Vc4/kOq0bjrcU1b47QADEzinJqXX/VQSjPusAgPWyAwB
6O9kPFJME8g5X/UwopKve8ayxc+4Q0lnihH19iCPMNCpnggY6ahlGqPPwbGg/81SxoMBayRy1WLh
kuqLsA7gnfI6rkjXblOvxRDxVjO9g3Q8SR4affP5AuXIkB712GUHol7IyK9ljc2vCM2gLHNQ+Q7T
n7fQ5UFuTPaz/GOox8A3HQHAoaNICUycaPqgtifJiE3yz+p++N8wnjjS3x4ZQxzrEDWqRVMT1N67
pRslaewUlb2yU1ROUZG3O1cESv4+JO1bwanXuMUS3guuMyr0r0v3Vly57WueKJXxM9cD2r3jQhPe
Arkfxtpv8/+Msf1RZHFwDMunazKN5flW3tsAnZhLS75voJwBbSSY7dV10m8mV3jSftLFgNzaZBue
/26i1mvI8F73rXYAwuQq+DNKViSjQnQjKM/8QAjcNPJevGeQr2a3Jrw4Q3rw8fZ02Gyspe988LdQ
eg9hWdbo5FvNhZZTQpMdWrTQizIcy/+E8mX8RG2pf2fzlvc6Ke4hdqVGyO8voJs8A9wTj8D0MB1Q
tH0HLmiTL1A7CoPsmUYjoBfR7TYGcDgyfjO6YE+7sAaH1/5amNp54IX/9UH19j3CwFBMKvtMrtFh
a8sfYy/fHmfj719L51iAGCVg8dbSNpmEAKsOzL8PxUmNfw+Owc01zY3wteKHwjNTfPBuXxlZJJhk
sB6KxMrN0A5PlgVQC9C330GHGCanqV7OPa2CsFedzVjH68VcelfzwP6kSVC8qWl1OJOQBVQlxdZy
j2VY6L4EjhrCY81jLW3sedRKOK21WCWBrXYxmttKr9+PYEDTGTHSGJtvBkMrrOphNaVJH208ht/4
WpQa1MG72L5/T3DsP5XFVx4tGJYOwOxr36QMlE12O9hqz626F7SleoQUkdH3lobkW8XzS1yTyFpy
gOex5+SEaISHmqbhu0CfWsr1LqXf9T+jj7lYBeqyPugYm24iPtsmLxXybV/bTFsX6YRRZxlN26bL
DbLGwCrKBTIic4bocIgaqHvCc1V3mHOMol8WGHqa7v0/NOspySljWZ2wGftVYWWgKTm0X2MDxREl
oM2SWAF3yNyDI00aSHuTqveAaagXBPW2K36GKRt3nbCeBAERJqoKfxqSnoePowJ9fcV8IrUbtQyn
iRV7svUqAffRXcl1CQ3CHC3MMQYn1PoFjg/05n7la4gXeTlM0holmEF2y8+KYZ13HHb7GbCsxorA
ydfZ1akKnNr+9OJufRaQoKCCGjDgpj0ofrVNstPu1mys8SIic7cIJybRoObFVrHh4IDuKSmA7KOq
wlzt40Ft1I/1TOL0+dd7I7OmfhL1NP5sxzTykMOD6CdjNgyTMdVyhUHnVkK9ndLLY1bq06JffJWp
hGk+Nt8S1WA7knlTbr7OXS0R/nSVYNZiKn3QBKnWr8abjDHMIp3ZfrvXXGgS4JSi3CLmh9Aj4SJp
hLKGYFTGgaGsPl5waOTLcGHOkC2wBLcDohOyfZSGxAOtQ8WQ8sVHlB1jx2lRH5ecxOqq7WsJ8mkx
kBQn0/TQrVdr3FOY+Lo5igOH9LAKfWYgPX2mnZmYjax81uiRaHqvHIoc7CwMLQyCx1V5LLdp1Ppw
SM5F+gxCp61dJ4+2VP2mAL50k+kd+oRQsmYnKswjZVyCTtOhMnfw9N7shnVGWhzUA72i1vX2qhLc
NKRaz2fIForDyLQGqSllPM+cLR6f2yBnistBVExgnu16Kp5JKTaQAo/c6bGAxErKh2SuAqyWIMbu
HY2KwXRni/W5pAxKoLSL/MzbNrV/bxJ6DbaGvnziBd4FhQ4gwLeaofYM0p6tBHjIALGpKTpZ3RHM
g3XHpM0ugW4EekRAjkWJjU3aCZkVRazi3jzAqJ8exlEQpvmXLLhUYz3UDjG0PaOsMWoe0G41Samg
JMxgS8Sx3O5NBmBcEe3F3/9XqyfQNN+FBPt/PK3pjdFXhwcjQsRUxShw54XsNWT16L7vzuuc5AzV
6augQMhlh1vqrR6BG9AsErshFKpk0jZ70TapCm7byIF/NgeTvS6AwHeTyc0547POZnHRm5g95JqL
IigoOT6dIFnhoNM+z4+agQEEnzuVBZbVLldEZHOMeWjp5sLWYi8lQBh+wo62Ka+iz7O/0q5vFE2x
JIrBBnb2ikHcLx33TH/i3ggm9FZz1e0ghGXi02dfZzi1/jm24aMmY8XXnfLgwO2I18u5r4JSb+cd
o9eD4dJli0+TTAnCDpkU7upE2ZmVds9JTC/B8u/wO8lSp29wlGjvA4apZTgxO/qdT9u9/tb5MfBZ
iTMWAEuCLme/PxqqMoXZq1IWe4qAakbeVBamV2FTuje5uBKutUJBuYN4T0iM1N9QP3O5haTFIq8J
YvnT/DSJQM42HHrS7LNVr3nuj8u/s7Yht3U6tEpbCgfyATp3w1qCrBjHc6nqD8J8/qNINuhhnBgG
P1XWC3L41ZMUfWOnNqum9r00AjMT1unxZz1ylw+PE09YEkBqIG0SfL2miFomHV0OUplaiicqz2ql
Em/8WfB7d83vnsetw1JpXWRtgt+Sd/7KDRpnvvGohOlp+KSoJ9Bj5y8pmIrx4Go27HL9kSsRsgod
yOS2jKLYB7494MbI6tVPn8BRQ/rgqja8J3SmCPH+h1w05NqjgXSE/4Ti3dLEjVnutIVLuU9NP8NP
UMZR8gRV53MSy8JhUESsFdr3p+9/u4D/HqDMgmWFXnjK8pVailkIxVgFWbUgWIeNUrKCDVFd9c0w
X5tg7s9vFX8lDi1/+8XGC/peXbpG2bNBGB0iImILCwDtn586XTQwrak+48DGfi1lLd+d2KPwoKox
rOix7NaURQE5ocJag4I/VmNTY/HwljH96ATDQ0OCU/NiGn7eO3zC/xr2UgG9RSFOpCR5+lv0vR54
rc1j0nuxeoVUuGi+LRII3kkV8eG20PkvdaH5L0Di35AVq7kfBbEXy35FsvVnSgJHDQbkZqY70jEN
DGiu1LO53oVIJzciNpO2nbGPA0KosZsG+47ZipiIphIOcmkX/PFeEdjM80ZiSeL73nKjipBKitPQ
c/kIlntcec0aPWCFsLW0fiEkex0EGQPv1Wvu6J55mhnuAxtln5YXigbiPVOqZVCtOGHOddMimvfA
iKdCH2Ty26uOrhdd0E/ERDGfDNAYWWUu4cO+7qgiogxfeieceLxpjKd266KXL/zoFta4Eoly+MFK
Zri1hc2fp7NbQACCi2r5WviZQngb1x4UvEZ6o669RTTkF3PVZcMlSGFgCLqkDNGFk5fmr+uB8Rry
oJyOyIsLbIKzNwOf4Q3TroHbTv1yX7L2KuG4nbQoY/5jRkEq2zklRQwyYX2uJ0AVWOCP29vOo6lh
DD1io1TmGUaFnN2dZHWoypP+qTxh6kiztFapPufvhp+2oraQlZbwGYOFOvljd3BEsDcFZbb+tvII
Tk9NzvguT0hQ/N326QkJIBsbUjdUC/ZeawbzM1ihTeGSqX+hCDhheJKnrXqj+K4x8F0+LIm47cip
njA8xwebbxPXZ9T/iEl3ifi55dm6VN28TfV88EE8E+NFhDHTPfduxijr/Fnex5vbonzDNHxTmapT
jg5jRK3bzNgrSBLz7fJUiqP4pmMTaBYIUhzr/juSC/O2PRvOClEranPAGNMsE1VBuh9zR7pgLBgF
z/4uMgCba2of3UGc0/VNpSjHYcdgEjqLsDXUgNDLVadvbyygRo8MfymbTJsORuuhCxlVpHqCs64K
r4HoeUX1DDHvdQeyRFcL4YxyQFPlTdBcmb723UJobLydwiTwhzWBtMm4dASjKkK6S1zq9jMMfXJ7
23zGpIxQ8Z9AEGKuYwx5bVp34CF9gu+uRid5fkMjaaeD8iI2eXIPRezoquudL/oZeR8OwqwlS8CN
La7ktjn9IhMsSg2r75r3zSbsXQiJzIN/5iX50IaZv9d6XBx0/ljikemKL9G2MvDE4lqRI2VFydNW
ixScq4QFfwGkaTZ15EjSVgaJ6lDuBHcLv1IYZY+sYFE1R78EDb4fGaBhiROlEaY5jRTu39neadJz
r4k/nBnveLH06xbRXQyZp4sC8RxXRYm8okCC9fReph7nW44BR74UVxiKTXZZCNY9fkegZO4W2l/W
SOsGnzAOhZZv8IZVqkkWB5TnT4ARmxKfhxi8ilWJ5KqPZ/30iYL4VQREtQovxaGpLRpcXPdS0kEn
/1ZOkonPwn7RjDPns7BHUhVUUCsZoaiMOCzMEUca9fEm9YTJ3PvuhnlfkD1lDThXBV44bprwNxHN
DOv/5O+20EnRnRRiejG40T6otQqhAwEKdYCvA9yScpjPyLVyzqYYs+rJQRWVgZwg1xqpl8Cbg1i6
JOFlsEBdl6OUC+eeANMK46utm49wnqJF7x6+0AHTLG3XSd2qK3vI2fOBcwcIyiwFi82kUVVEWfyG
SRy1prC24wGmeawvzxXsKUgQQ9MT8JqBFZbX+H9rLdaZatomL3bEZ3CW9B9qaLAaoiPEDRo4i+l8
Qi7yGO9Whkal6SINdoy5q2XrMeSbozv1z7gNLvFzIX8s50iPsq22OHpCVZ6UuYvd8KGrbs3DEt8P
YruD2raPQhPwgPombXfRBMscM2dD0cJIb5ePDYpMn3wlwYpibXWCbz0OBWI+iS9vlfIfm0p5hSM/
zPem3oHEKZ4L1fHvXGp8G5CCDxktuJrOAXN87WTlfJfNSmnopmoIS/Y/+uo3Y+fa+TW8+oonT+P4
JW4D4zxaCAMrhMb4VD1/2PZcKhuIok/3lQ/l2lx22kpMkuag+dkwY1E25Xg7sHriFNVkiEIgD7Ke
5M7jpokuX3DE2ZTil+WSWhELgBs+SwebaZoS/33pwXA+pHfs0kovKfeNP80qBW6WroBwKy08PFQb
UOQm3HdZi0M4hmZnGnqMthks8AIs2ybOaV3VWefLeElttlKu/kSL8fNldBxnR3pLdfjj9Hsfe23f
XuXCfrWs1msH3kWJRlMNOEb3ExxGV7WP8yuEk7IWvlX9o+jKLZGeJE/28hZPFOYyC4tBUoOjdHx2
vouJ3LBjPUmRXyaXPaiSuaO/UPDKiVVtXhkR1Dj5XbIEi6+Ink+Anbq7hX5+LMm8x8GfbQR4/tjr
8wqyhMA/uwvjbo/QMDRyLVQ2bF2q83hCo8DFN6N5f7JApNQivdwUY2cpwsetAiwVpGIbnDDc6a0f
wOD/2LeyBklO5I37lPDexliKcV+wolEpQNyHDvvDZNteK+nanBjn63bhUaEtQWXUjk2ZZIX5hDBa
A10aU7/g2ppnknM1kzQMnUeya09u8m7JdQK5uACtuiJF/j+1bWFTCl/FwqkgHnEHvjn9TXoNkoFp
s+8HKspvqi4Uc/KkjBWmludJAs+V78HUCoXplAjZHLZF3BdjKkZTTkeijD+ynX5dqLxQQlHk0qYx
bD6pw9HFz6XWggquKDuoAohwbzGlPiGwce4T11QgZaMV/C1OOLSavQ2fTeEKa34jnPWmHiD1QAYf
OJUfiC15OqFKE/NQnB0Kt1VKBThmCIWRHR3c/Ce2fo0PioqOKeMVQeKGVuEKbZnIFjRxNK44h7Yj
tDMa8w34YALVEDCu8wg/zI9JU/wcQQP1HeHpToO9EKVJmrAa+LfZZnb/N/1jjYU1uxaYvfHcAQvz
FHOnV74SWPpkF9wdWl7EpdtSPcz1JwgRSolpBP3s9WnwodWa0mZ5MwU+L7G0kAzlsEpGMPa/i7if
l1F1x68JtIkM8z6BDGIJzqRlMzGK3yXh9VDAcx99fy8LSaDVyIrCv2gVKzLIkn7mpnHSdeIJNQxo
BIoR05dTOIBM97fTxwcLcrNsfxROz451X3ezjjT49JIDPgF/4C4nVj2POEEEiClZCOxtN4KUCI6S
WQqTkF1MHcY7xya2MBtb7PzYiXMqb9+xnJqhnLYjAT5oAhl+OwhmtvRe68xX19CrbKjUsWOnts24
l+XM9MfpOtF5fC1fEUzZ9Ep1Fd98WGiQYLgKA4V47M0MJleyJR1sJd1kMFxmGoS62anzR1Izs/oi
kk2yoFIalnkjAdKZpJztPeSCQuN5ysG2d379Kfu7u085Dz2+LJ4WA6zPyqnNTUtllvMUWJALHp62
N/+qJtF5PXXSqjMP86Jgiaq3Ki9Mk0o+rM3K8bd2BwBt1kOWgC/NC0Zw8APxWvt9lGrqI/qgY6Ix
azGUe6vc+rfFVMlU53e1NWb/pSeivus3hdPVQlIM1qtjVWBXOogw9HQUk6zq2XHOo/jk1JV5Ey5m
/1PCfzYslcPTRA6zHW5h7illO+cMmz1m1ewSXNt/b+rGHEUQguCP0TUJ8dHeAIw6lTMb4IsSKkp2
CEalBD9t/6wdMajCAaV1flgWjd13qUrNryUvTZXHfHIHzI5K6VvllBWyHpCSch8AOMbsIH1t6UQp
4e8cfdGwecSzgCg1kxjVjgYeIsmX8SvXIOZcyccHq3g2igDwLGzjfFBlBdUFMOhCyIHbuPlLIHps
7nGi2ETBiQi/KKyXvDab2KXvK1O+2Q6MjDvyOQL7NQ6/pize6yQPRyahNSP9CqXeK8nGXD8jah6t
L5sWS9GekQyl7TKFVO7NyGkhT+ebiOitQlAdx3a+aI/wfM2x+Vbt50V2Jqf98WrBWcNQ7kGY5T/8
51US90amZLbpX494lt8TPNJ8ahilHU7Q1z1DeVMTmbhUcrKjhyFGmaID/VgndVaEGLC07wekDchI
A0W55hU6mIRLvjbj6bVg+6Z6OaoXv8L3pIndtbHiqohui1/9B2xC3afEuoOJlaYHcQ20/OfHMPpy
1TtpeczeCgiUN3MEelMbPahx0LYxMnqLmp8i4a7A2GHlSrsB04qFpuHboEp4vULZjdFf8zXeYRjR
lpS94VNUDnMYRpJNtPpKBncfE+HgUuLX+5OMDXTEPdxgXNBIby0ZthBItNOKh/wVaXU2JDV/E6QR
ia6xy9dvEPwORVNG9/O+bL8LUsLThzB7LyFFI9Rvqpi2ofnn13MVrUjaiUo2mF+eeVl8+C8oaEoN
M6wjmPoQDpheIxp/Gd6ap63tbzZmur9QAaogcan0Ud4a7VgwTa4D5kz4tpTe8xxDCaE/GPBATwfF
Yy/S7i0zCoW88c49d538lTx7PI+4j5NgVc6ap2cmIlz3mtCbT0ESKEwpmWEZbkACfYzbWRA6IdnI
MuVigFglQri3pFkFWk2QqxmZboE2DXYAJSU/vFIIEFRrnEWIbaVcNIkbeQRDXkV4lGcYPs7Y9ZV1
5P3VPCyB2HjfbOy1oh/UKlF0iCqdgW5tmTQ61xN7s7Mr/lIlzXBm8xxZtdqEhdXx/s8a0ez2SF/d
F2453fX0WD9U49gir9A9geJlzvQ3zEnHbV1wbfp7n1uUeqcimTBsF6PQZr5dmnPiXkd2DCv6OwLs
jQcBoarRne4CTxCQEuViOdIDVp2UN8qjBFFxpBRYzQOBB2akUccSEVpZTSFT/SLiQmrgnWDYeZ1L
8PAl589PgnlFn/7bRVJ8UsGr8EfbsqTWAQ1Gc1KF+UJYwf6hjizPnfYfaQukgpHQrLjJcbRCxn3t
gawZKzPfQIIcUNKXvgeu12XrDuAPzo7miptDAzzp0H5yPmHFNMWg0dZJF4LewRvZXZLWgqzSaL48
yUxQ1/9HkEnInLwtyoxKHlcLRVXDVSsF76u+1ln5PtdE+l5kO85nvfnT8g4hk9pw4zGhvwz/IyZv
GZWddH+1PYLLsdM0elRB6S2S0rRZODiz469oH81iy5AwhHCSmYgeHuDCsg5Kbqncy8LxnV0p25xr
PfNw2c3dwARc5lgs+9MTREg4TqgHtX7ftUwkE7HBXSdveWaog3rVbS42MDGCZrvOAG8L7RN+wunV
iJy16H7dM1A04JV/nYKTlekFeHPyEoq8djENevITjkeTdZDvVW2CRIC/22kooSGBAJfonwO34FuC
hto0by3bqeLyB5aaE39MKEsKFMtHsokJCGm2e95+ChVsLyd0Yb0DCrsAYPuiED59odvtTXSSGIPk
6u+6Bfvqbr8/kbAP8QnIQRHng1E/2x1qi/1CeiDIbwQy5fC2kgeejDtnH6AF1ZxW/EO4AQMZtTAP
73XZIwXUW0moccMeyRu+s3/HHwY1+KHqJkzLsWln502bVildNwXhlkA7dlLeWI+Mhbyi8wPecEsq
tx1HHP1l23QOWPF/RiNKvS588VVVt700aYezZkKQwNmVoTIb/ltNzBuL8ODe7DexNlxQNOagm3bY
0sI9weJwLlOygOqEMrIIpIA5jvDjf6pCiNwn1fqbrwJUH6bh72d2dQi84IcxVBKXTlnNQDBy8ypK
fTCRXVusZn7FBTfF3ibw0V82VocnGuEna5RVGI3idxwClsP54sKtS3RWJ6O6QHsbxFZlZC31bsOc
xG2zNyTRW6P534Dcm7pgRyk6TME/8hskPpmEcVpuRGBCFY9gaQ19RBlHGDitOZ9ikYlcF8looE2A
PSpeh+xjrmPPAMClkFKJ47eA99slxaTPDSVEaEhkqf+P5UdJW9U9YvTkvPTzUpOnTyYccEFzDCC+
ZL3oMy1PBqwh64pCcPjxiUzfVfHqq+ydGROsy/8ctvAKhRnudgjHeTUUhCXwYeW4hymQ34h5FvQg
N4VnSFZmPdhtpa2z3kEpPyyDEOLFS4/9cuHnetdCWy5gPOqXcxhuFdPS1sbbkXZMJy/ujR0m8fnV
1Ol3OVkT8/PpNhrO62H4yGc+bQzgXpQrMMod+51ltBWOosp2JG39M83E5OJ6zVb0McvLMDQ7g9jy
kEPYD3AKnDM5WDiY11iEoDXxorvdJpjLK5iCNVF8lGUcBfoIAbjs62gacenoA8SGskEvycyWfHYz
Pjza+PTq+Mnn90uXds0YBMyzALp65Ax/SKA7hbj/fTkIYQ8hVXXCo1/zBKezNu5cK/cuGUFoakg1
0b72l7S09DDtrxJt3qVc192IlHQ+YXzvYjySzhTnpve5vivHBXw+BcSYxf+CiNhNpLoxZOylVYEN
vcrS0q13d8xTmcJXlwEUQ2xumtoaUo5tzv1Jp1q4Z8qfu46pDGDulepUkyVEzozWYe+NxfKDaEWP
rTGe2pr12g/45tFEy9TG/GA86of7TvYhg8JGwV3KgElVUNFgAiRfrXODg/LvOGnoLG2RXen2+9TN
4o5xAK2vCj1W+wgHQutBf6ZFsHY4JYQAN+O4igXOrgieRstHaW5R1daSBObXlk7HgxM3oPdUvVz1
rEamddDTkG5WQkOTK5To+Qe1eJ6yPnIxbad8qGZjQqQ115y1FJu4tCNDtrvSstt4YHF1r+hs1fDO
1RHgNdjZ5g/MtiIZOrG6oix6GoIbbGRa+tDLmjw+zvI5+LMXReAqSpwtwoi47+RwQyJLaeBW2LjE
28F7UY3V655F814dHx+l+vcg/n7Jmq6EChiMZkVBf7EFtlyv/hgWuPcCPVLFp2sDoOBb5kmT8n3m
YPVs6K/3z6joWr7fVubCJ0jtYVAlMZGgDqcrkWlF2zmXODSuUJpRZowkzFd4DGnWutHkQdeEDXUc
5bHSceLEs4DXYpsDN+/LxvOeCZaoasS9CaaEvutzlKqIjv+p/aKvjXaO3H0TjyVt4vWlXtAr8Sk8
YSXZE8WIQpzZO3h3UqmRkEso/310oFZ9cdS29IFB5O/MtLLIt1hs873bSpdwPyQKYrDM0ea0MFtp
f2vS6j919zwh1kDi2bhxnNl02KQaXUrGzPGbiDskUW9VcnpLBiF8BBjTKZ1Yer3vjNR+7E9aw2CW
C9xRFNvKgR8WUfWoJ1p3Q7ZeuiReygvW6TFHHFjAgYlRw7PeBUqewJ9ZFb31TfpQx1PU24v5ljgz
Lcq5v9GfLTMNN+Lft3wn+4NJzlCWXXo1av6OjHBH/UQrP0D6tvbJC55s9zoVt9kv92LUrYo3MDZc
pU6Dcx00upMR1nbOzJoyzQMiFPUbnNWJYuQEMVV0P8aKqs5eT20Rx22bj2gv14nLOxzzX3MN6ZnU
5z69FqXNW3A1M8kgGl53WvF+hFXYUyWb4tJZq7psxWeqFjuGDOVRf2Kr5PhbrPuKT301vJjRHr5v
P52r7X8IJOm9Kb5lyOWMhvDmcPlX+q8Fb2ESv2OIzkNgvGz/ApyEzbcA1TSPGhx3KvnShUGWq+MR
1rRUhKy5QlMRUHtKtUIeM756pdPYVPcoj1O6W/g22cQPstpnoL7n9B/zuVAFYyQYdyawDa7/YACd
I3SsWB1bZ1bBmCvLpQvkF5akHuYAIdvGuuNI45D5LkB1UAVbAb7RaGIVb/nsSRDC+kaN1nQh9h1o
ID4E88ymAV/SMCaQDOdM+Cryk6bJ4jWyTmQIGSvxq/H4RPySBImKwi2IorsevUZ4vHUNoWVSs0c0
LZX5noHKF6lmX6VUtc/x45QtJ0WZL7UL3gaibiusw5rMxvhsAKAA3vWqlfGqAhCFtKwwBa4qeiqU
GytU5uSMYTE/gWnAIHwyQ1ukTYPVQjLtY0wxCi3wyCoY2sJK+bQgUuRIpVR1HKeYoc4sgc27CBHL
AQI9gO3u/1X5oLFwD0t6xXCdbEsyygNJcJGbC6wz8DWAGK9vAA9vMCOla/H1QqvECDB3wFCFQSl1
FM2fvZQwkCKITIZ07/taQ4IJxUcV5gGf97VZKGwq/SdEoCYU4uClQxMPKje3lAYmnbrtAI6qQrE4
pjgRCi9PyKfILxV50AmInLEWxqZwrOF9yiL16oVz+8vb811NWK4K4DFo+iaLbjbNRNbqqI+lHxx+
v4D1HPT3eOvAbvDM8ZyF2Gf/cJ31sVoU1R5L+1PmR7wOKUd8r9o8K/S/5jCosrKPcfcd2x1KQcUU
/20HFX4R7jLkiz6oqsDpeEaHQRJ0CBZrJITadAcAxK+c8M1FVHqB43LbF4qHq7AD4kdLfMtd5RWD
4XK84J+Gmf+pCWb3wTy8Zg0jumqX0KEu6sWOlIawxLN9lzE1z6xxFoTzkxIFRdQ77DPcjwV1PV5c
+qClODXOyVGuj1aQF6Hv2Vp+mZ898qAs2KwrtmJIrwkkUr4cTDFFRUOBL24rN/reT67JMjzIy2yf
uBYR5KqC2FG4s54rBMiyXCE95cYGIbStPK7vQEU3w4nQCOHBOtTnHijNV7qevKKj7q+0u51Q6oTm
lsPuSYcNILrdXFBel0wHcrakdtaIrXvj58MG0Dx0hY1nFOlBr9llUcyP94GcqMe7+YraZSMZBBBY
cmVaImIqwgb/wbMd6sRTkrnIXdY6Id6YQ2TZxxPhQln3yWqJkFBfOS5DejHE/Yf6ArA0Z5WUC9/2
tjA1qu8cnLvmtlLyqdTqwkAZYuQYIEmYhpms9R4Uqtk8pt1Yy5k5340/y8+yUl0xuzIgfx/VBVtb
csL4iWupiZ8yAYd8ftQIsK7ZeqIbq2EZUZ61g9aDFvWsxNeQCxCT52gZMGTt+xMPdBrvbVCRDau7
pc9UJ1WM2DYIsPT6LLneDnlzM80B/ViC5H3dn36LF3Sa4xUolXFnsReaGnOvdqBmXL8kUqb7qsEc
bQqTLCp+DC0Yak7FHKj96WQ/EGUW5sOKOwNCt4vAdQOOY89Cu+JJ/oEbMxjH78AKM3DPh4EppOqm
ln1iO1J0m/K+C65SGT78zzte9XWN54bUXtvdpOn9nN0yDNbQxALtXJSrnRbjjno01rgoBj/m55py
LXQTYnvPC6nIzXWNDpWxx2TQl5WT0Wbr/Jg7Qh5917tH1Toh1ozps/EkEips2/+NzCuedpKSt/2t
+cuRgulqXQ/H92oJxLfye/JABQMpqKBOvMgwjLOMzEqVbpbNAPHpBPc/JM+Bd+GoUxMucCXXKwxC
Qlc6/PXzlIyYTowv43VkDZoXegtMbQdOrHbVu7sX6Vty68S60nMs3SgU6gWjKtz9h5jveu9k1qHn
7tHK463pSjSSGd8p9eFiq4ts3FDXCJo9AQ098QikFrjTfxymBooYiUialD7ZxCvo6yXrp2fM3mSS
Xd0W4WhUAWPYSmuGk/SXXugVDmeUHfHjM5+OP4uKcJLESTPj/NLid1pDIWnGX5xyv55pS2DSKJ6B
K3sNW3U13STJQ6rPfhlrkrDHcGm81KTEysFOs6+L1WAlNz391U7MKtIKsU5aHU6saFknpRnplHkO
d1IPtbmu414m/rdgAMvUiOq//GcfTeOBfmSY3+aoVLLoQNcLAfhRPwCTskmQGyQfjgeUlh08naIh
i8Xd6wCsFdhQXESbd9tUpDtml24q/rsT3qEn4t8cIzEAXk3ayPv7YR7W8ElPMlbtpa0XEviGF0va
6TcPbQfF7kkJrKkJ4xr2jkA4AJhjffbJuh8TnZWB5M1a23O5WtUN74yhhs2RLVqrZeo6cZT6MKIu
Lil2OfcrEY3WclCybkM5jd5jVa/7BWRsxujkWKDCRdcibHTqKHKqQqEQNj0mZAkMk2EVz3XWErF3
dfMrOuDHKB67LTrmz3cclOEpzbYEs6dLDEsG/LTb6KBrLyJLD86sQSzCV2JHlw6qKTg1h9hfmc8M
cWzF1wuqgO+YB5pCHkpFFaxAIGoFLHaZ7kuWCCUVF9G+3y6ywQTgbUq4esBveJSXpGkE/jtuyR1i
XWrR0SUUiYmuJ6FPGwzB6u4cUP1aPmTd3RX6xVrxtWl2/a0ZPjzlQAktk4i+ggst/63csN3rnvxZ
mqvaa/Tj526nJyMBDMTZuhN9QC+3rBlSr84h49lTyndAuCeTfr8VrQ1kBqFwUZfaS/u/NdWB7AsK
+cAewW64f7rTiDzk1Bai2T9z1AgDUWYLl2sNqkWwRJk2o8SNjd3QKfSptFy6j53FPE2qF4+6WMz0
FuBkkLiuiHNTaQFvr5vaaeR8KL52CnD+TCngjEklun/mKLKrXpDZmBtWoqGr6X4YA2vw+7seAojc
PF69pOVErDy6KFW9b8n4cspmZUW9vAQ1uWTpwCLiRTsiyveQtAqeD471OLzjmJRzYxu5Mc9IBNtQ
v2QcUSRMM/T7ANsN4bLYEwVs9qms+jJmb5/GFSdxl8ofCUezoUZUm+OlNxGnEh+Tu9V5/dcvjeQX
nRZxwZEELopU6itwlvP1drsNm8nF/lrQOgMIcxlr/UFYKy9KZRWyqUvjMRe85srwHedTopxsmWmq
HHl0XQJzpXd5XnUyU6HDihiFeI9BNYgy4JTc9OydXuaPmB7FEeG4BXI546zSAcdU844txK090EZT
dmnE1UR3CKNKtS8LPZArseRXfqr1A9ZVFbJv9gBSZT/TAi5oR9OeKEENJpEyL2c7PUHmZVp1aAYw
s/ICcbr7fKGalsc6IKL2LJlRt37dVr3zHkjjkRvgRkyT8cBHLNkjoDIq+4ALLmkMtQtjnFrOqWsN
USxc35Oe3whu9FKbHM14HDnEWCFMdDy5fxhOWz3vqm8NOE0vjG56cgRuMgqkYYTMB5wKKtHnUItN
fFzplJkUE94tTRvXy4HP/qHrVvybLytivkJqQbQ5bdkIA1iaUtKS963KqH2j6bZRgIng703tsDft
otjtVALFLAZAiLCEJxJgkuAdvA1MMRbIQtG1YsypSfxmMzeGB4lLBjUnoB86MKLv+Uq/Eaii7SBL
rTJuvf+pH+UFxJZ/hjPaP8icKNbRFN6XlOQM8sG0IpvVJQoLTjFqNvrp+9g4bg1YnaUPsN1uFgOy
kT41HJ9leU55XHI5vCiddaOXhzQUiLxn8uHPjiChMQjC+gq5drxVz51nqvfqxe+fZ0hJEGNRBYlw
0jhzrKqyOmYrY+dsPgd1vhZOyx7Ob5xDnb4ZC0yTEiHJDJxlBmUhAQEcN0rAKQbSUt83WzVaH8ww
3yGEtr/2u63HkGRDriYW+RbDmv4Sj6cTQg11lQpEk33psG8bm7msfnRJLKwUXP4SPSFLja9FVMqM
3ddfYsQudSbP/rLMYOE7NTaWJdosBDtgX+4i62m/Bu5er74CLgsaaweSDAxJEvMEajx/ibprJE2E
8ke2hfeHHEeE2ZAYLzPbyY+QUXYrNTdMyWq6YtUhZ4vOHLko6euCtMCUPkw961kpAEPevzu/LV4O
KrS2S5bx+a5leFJvORpp4fgkhyISjuXxXg3dsNpyImgDcjBKQ5MRoERcM8/eNEOJAS3Q8Vx87b/7
Ipsk1YFXfoDfFAdPSnEwj4MHobga9Jea44F2d4KcM571lrZczvYznG6bpODRBTPTZUCIrIVhyxQf
ad8fxYL3xwl8bTnGiImwdzbax5g2ve0EiC9lHb7RdEJ8bwneMSpH7ttIBRs/deMLLg/Wt+qQvEZs
WvmGkuxo5m4UpyCuJMZ1yQXCFtgsmKhxIn72CgnfUsd5ORGFsjZOx9e4sWqDvQ79OCDsqmvNrLyb
hermsXEj1bjbSshjx+DkKU0ik5VUsTbhIzzCMjrEPiNWCMxNj2sNYgYvqIbt4LBIVPelDJsqhY81
C/qisU3/mHUiX2OXkork7xoOnONRChcE/EMo+XPPpJ+53oCScVVRCRj4xfyrr7BaHL/SH4/TvSmS
zqHZKH5YE8SxoqEqcuFTm/uEqsfWq/lrZZNKqqOQBL56xyjo2Kvqlhc5AMu0OvIftyK5aV++xJpv
ce9FJimLmlXLPdjzlXR+khLz1cp+oeqaqJvZe0VJ2fmIMPh99J+J/LPvxqcn/0w0Sez5DKaJcHq1
jIgAnXULwPkeQFhTndbXqlgl91iBIlIJjhuniTHXnioiE2AHCU4EhbiSkNa2W98UnIctmakA3k9H
pdtkLI1Ylv4oUJSGoeC46o1olKfRjaJls5gL2DCWnn9meb5gPKt4fn5HRdI0nHwLLASlwqT5f5iG
SFc4lhNa01sCS+DLw+54A0ru+1UFkzySYne7qYjdo1cqtmySGB5VaAqkC8CHbn9WTnAkd2kH3JhD
t41sie7bzzJW842DZVh79nXlBoQswVKZdHLgGqIH0018zNmWm4b7xg1os58FN7IPQozOW/2mYIJ1
JXjpFRFoBzUN+lPkbfuKjQy6Li1irnIGzD6MNH/eWlTw/MxGS0T8S1SKVyL2uJYLKEB7uDfxtQ85
YyZdVAUDWrXpRpwdsTo/qkpXNpHh0PzW/WbV/hNGmMHB98IQY4b9yWb6tODVhHlRIBYklXwsXkQP
oENEdHlXQU5A5OVY51LxPVWtKk6c9n6CpdJ2pqzvq6X9lZr5M+3IkeEfACCZbLMWahEIrrGR/QTh
CSuUK59PmArM2D65p3L1HV5U3hJAh751PIRTU2qn9zwql34lQkdE9xBA3JABIm6suRAiXROjikZv
q6mJrlhkPxzHMo4dNFdwXSuTP4R+aZ31ZxsjHiGlStnluFt9HTkG4chvCVNL/d20XdgbEX6gSElN
SR89IgVVKm4tq6WprrhpTh0nMkgKirMavesG+ujhdxf/qz5fjTXRAobzg5VC7H3beYEd/H8MYBGB
Lzm9J5e2c5jt+Z6/fqdVa020hDNIYddz1aSpHagbbPSFsHp6GGWsT5L0b7M3JykB8maIQidxrghR
ktkFLWb+63iZfSRf0T7yEHcuYlvBWIp0d7JHg9TBdJF8+mFOPaRkWft2wLxuZiG45YKQmWm8uF/e
DKWrUx+DDtqiGchhXJPUd1ddLJXlCBRBnENGxZooZ5Ygm3cYt0+LGuEm7QcDRgPxnBVBAkSxvWXE
TNsi07bmPuiTUWW77Eu9Ua7ytC/s/V/sTH8lh2POmQXqK4wPzarahkkRAE5p8C7oPPIOpjjS78IN
vs/lAb85LGV2VQFHKm5rUKp48cvhScQyZCfhG1jxX4LHgJuMWKs3WXOigu/Vpj8xmBGyMwDH+SNX
ogaoMCTCphKolZCCztu4u5+nhaPGQtapgZWNEvRx2FFYl9ME/hfiw4+Y4pYbtXBX5O1IkqSMrkiH
QProZtavZqfANl4nsW6LxfONBYZR8RHBzbE+DnvGhMpYGMYdky0wswoVLW0rkDR735PG4Cfx5BKj
Aam8Ep3fvoJ68p0Zje0sUFMQuDmwjPEAJ18FxlfXeNGoyUUSulmWanMMIxFnWl/aQa9Xd1bsRtwS
ukmK1G4sTJ7t+gFk1eTlgXprUEr4Mup5b5B0oaI7NlTRgtMu34V3kEKaJQJ2Ul3CUhRhbBS734KO
MDwuQsEyIubH2uiSHZn6bxRso7u1vFrfvHhNb7N5yQQSoz7PsxpRMq9QfA1aUNm+5MPdeRVYp6YT
p2lwJgTlRJ9OzGjabXyRt3JlYeLsWfvl4WJn7iBwB8+Uiuh/E9qxkX7WRtu9ApGRkQ2aSAPI5oSn
JYy0PNQtHZ1cfQKlGjBHvbo0xWlWlggnb8mk8/JIFJh8iz5GcSMb4/Zu3t4U1N69EziSRVWHvXjC
CCFGy+sPfs6HEtrOR3XAJD54h0MTSs8ZCe/B+CCc8839lGCO6sjsEQLYxG33fJkUxJKu7yvsc6fp
arn/TmTv+7VnkZXQ09BxJ04F/0uS1EwT0UctWo7omK9zgCMWEm/UflHCYsKvrTB9Br9au0DJrczt
96KX78gVR6tsYpZrvAgLhCpkz2TyZPXErRYIMkG5/kbuBY9UFXnXN9iLYpKia6Ifr7RFVdez/cpp
+rLKqW8HttGM1MgL4PNHG0rXlqrb4teB5il2Eod+0JzzAaKp1puk3o5cDeAarfgfZXf8D0Yf0FVh
1z3QHDk5PadotYWrQHLa5bF0+v9b1+vzBvMoG1jWP6VubTdRflBcje9bkOnp2PowDDjOPaSJ7Tuk
3uQL47fz0VYhPnk9hfP8Gx+0sf5bzUXn9Fijqmy1kIX1ueCPcfOfl5BBvYwyFWYbWVRqF7qkh0C8
IcSKvBfx5HzOw0tZTWEXpxuxVmyBhJkRwjV6uC3v3c1BhCTbSB8HMfp/kLj3fRdSraZ3xfkg3zrD
Wd5DzWcimht65XRIjTWxh2VPX1o8U83Uu1bYRrWQUcMkTuksQgvb5Y25MFyWkWcc58yq/YcDlFlC
rRmTjm/533pdUIxhLVG8Tj4r0p2IyIM1Ow0aS38YgD68JWTFrHx286rTvDg+boEJVIvA9v4VoxxE
UVnXREWN7NcXgZHj6WqtlcSm0jlc+CYlniljIgpIkFI/OVBAHLiwETktMu7jTmcZYG5sqZ+zHm+C
loJQvVMBuPtLrD3lCW/46gW381cPngx/JotAmghQdAh80kereKTE0IGR7C06641IoyXrg3+DLZBQ
w8/i1UqadR4mOxP9T+fxKSiIz5ub4mIIL5FRjuk18VMVmACGZ+SYpV9bocUf2tXZTYUXwy98L6FF
wHBDI1GSUXtBKBCfjzneAmpkqV2LDdQwNBiTxGRaF6cWghLcaaX5LCqN0O/KaFZy+jAP6lOmrTzj
wiLOjOnElmw84AtkRUkyvMYrgBWMhZI4M/PygmBlLiM22gXa8i/86h+H0hUWUEqIgOSH3v+/BJrZ
gsTs7eweUfsrEzjrYh2dbmyqCw9EryYUiP0PsZmII28CK3SSCq4y5wIWelvbu8qsKwn4Kfc9oLKZ
O5BUpFIqYsRXpyDKATo5U0LYGj/UfoxVO5fdSqAFC8FDW1Dubk1bP4iaN9JnK9BOoi6L6+f+o1e4
tbfvr6hRBFF3MQqMTAPSdSJqxPaP2SwtxUXGN/+GH6EQVu9oX5yMAT05KjGGno3qxG0OvLJE+5s2
YRlTbjiiIdoaEzGX5Rbv9kpbbJgft7DcsGwmnDX2sz332Da54srKhFxrMuQKe0RgDlroDDzlkU4k
fLdQ/R8+ewNnvfCXTv2vHOfXmTOpwhkPrlC4eLkL/aXoc0lnWDL7I3qqQdHLP7U6x8eIYy9LxAVw
n75LA/Z9EbF3QXlQla+l61pvD/fIkIJgywvic525udiiS3HEATBhIcZ0KVnszm+Y5a5JaShimuRi
vJs63hs9Ay/RXIGuLtq7P7hfuYyTA2FYTO8z44i9x8TOj5CO4YmNgrAlrw2XzcwE2MQ7YpA+Cryw
cIGsCrGKqiPLZhzPRilGm84FKCD1N47PNbauBXtp4y5PKUjunCswVeQVtkpcEMhxLvtapq6pWwQi
iuXH8Ho6MK2z2fn2IaSCZF6xoCfllCW5OAWIavgTTZipbdys+uos6PPDJIXARnJoo2XjxlOuQBXT
DlUzz2j21li79hNj/y6VGqpV8he187uNxk74FAO3HATT77AxezT+m4ZdIPGCY46UH7HSRKvKyCl8
fEcIcd0vPy5d3JC3FREnLqinHurme0Pchz5lbyxwPUX7hwlyd/1FBhu7boZ1ofNeDZxFIlka2snS
/7FjJxJ7E03lHyXzTajrvh/BS3ljVPLl4cqUsGZYxziDpQ+ig1LLavyE/064KVr15fuqZZIXkqZ/
slvVL/D2mcc0jDTwVr7CS22KezZrcqcGSxoI4X47i2AgXgJH8pgcaU4rFQRCzDv6mKFAJpnRExE/
BklZpu5TO3eKIY+mH43VtHxEBKOXnSGRGAQl4QoUnXcf03BshPsL1F7pGmr8aSaTDBWPGj5KSzbH
/DgEwIW+SB/m66IHB/pOzAaH4/RMcf4XJ9YSumdqjC4OzpfjFLsf255vHmYLByGMADQUYKTO7mpU
PLN98U7wyXTkdH6iwREKE8wBmU8JtwKOSTSPajyvKjMs3gVrjlEkoI2OX+zzS6Wvh7/Y0Vu6myQ7
GLf89hrulH+8Gi+XmtH3Ub3TGmaLrPqj/cLtKl2M5U4QsTcAsXy60QFQaJ6Tz+Gvha4Q9swBkrhW
91aKyIgTm/phuE7/hqYs3DqmHX2paukHAazKWznLp/C4YEjuXK/HSzvSzSFtW6ZsL+4n0FaTROXn
cWQZunYCPVNo4UNP4sbB7Ur95RVr+EUhVpM6/NI4Y2EJyHtpTZOV2RBiqepghCBF686Sb9s3dHt3
yLJedLURDjw/0ddb+R867Qx4mbTtEoVO1gaFbgfNyZKSC6iVwhLk+45L//gAa92OTzqLqMlgWiLF
Nj5SDpQFFKOJ2TQ5UkVW6lNeWToM6LR3juKoTauz/l0GoCqFxRYTBTXebYU7qexAAfFnuxAN5rOW
ZMVFUiaTWOUuAWi9wqsqVRCxhyu4FNh6zoIpE1rP3Ghlq+gc12mkCukYrO2tbYwDrWcn+bZQLjlv
X77vWUiAB5EZ+s0gzjQZuuGiHNlIMs3oiJr2SLj68OkIXd48Rl2SUKsc1QlDKiZ0eZCv5dtD6pQ6
tqean8iAxpjlffB7aygG7o5gXCmoDiKdKolqsvgZmD+FzEvXP1HEyOursefVNC2XKtSu39fytjzM
iWJrB8zQAEFfS2xK8EKz2BzwdWqeODRXukXd6seOiGbHlYT8HLTN/C/LYrTHFSmxp2HF8e1pVn3o
B1G0qU/cikzLgkJQBW8eFa74N6KjRqYaZtbum4xX4OOcHumeNWqyvncFS3Bu5qbgVhuo/ea/C9OB
4K07Rv6xuKL8N4U6PL4h0SlZl3AVaAUBvKevkRhgOqTM2/LDm+uAxEJAInYArCa16KZSNZIdlqe0
765HDaQaTMPb1gIbGde2HEuZwD7ey677RETplD+P2kt74MZbIY+4yI/P09I2h2dZG+VTtHIHoWm0
zbrZ01lxjcm4Xf6QqeiCIcUnqzY/dXTb0xOTL/HaBTeszH7tts3mD4neLXYlbiLI6aMSi+Tm602b
4URVrc50bqPDDFRKe8C5LrwuLawhZjyLnAbhdU2iRGvlTxdbnG12t9fZTnZiuGaywZlfyNei5NT4
UqmygEXR0R+7BaoRLySOS4/biwS7uiuJSOJnrkaw2bmb1NY7JWOox4EjJ3GDTbnAugTRWx1Dg20E
XitAxi40yTWWCH9lhkVvMKVq4HaDQbenibqyTP7NQUFVtxuJFbiXHcL3O0mZXC4CcUEBOGEO+tEm
qW5VEDlEdGIjUhpI7/aW0e5+rXWFhWd4kgbW1EiZW8qKdfzylB9vqGR2ldzePDn9kx4BKqkOrj25
0fDW/ZFkYTwYjvwnDJ3lmcRgsLu5XOWbMG2VyQFs8uwgeCrWOM8d6wSjwdSX0fPG+foQGQbmJJYu
GYE811MMzEJOwZSaZOs+U5VQenSpalRliSicg7OcWVgaZMC1cbz+br/zqrKQuYYMCQi67jqaeiJy
gqF/AXt6rpW1g180u5JeSTexGR0luRi+uzEwetB5xUbvqXmNt7v8vD3C0AbAWQYQ0sHuS636Cj2/
8r6yfT4gcADHYj0qLhiUx7KvlXvVRbCIK57dSRqgEpAcs5ipFkiuiXhRV7M69AOtPHz9U7J3wDkx
QQY4rHQXnsjTdEvHHslIQbmteq7zKCndPJmJPhfmFf38N0h0qQpk/2WeFS10CXoewTaqLqtgIxHH
QO9VuVH/NiMhqGPih1swLkTHg+AyQ+izPYWnlVGnnUufEH5ByzyTutqTVsVxGc8+RVdBAt5eT6Zd
znfd2ze/lyEmzOtnanf815vtfPos+XEW4GZX0fE69dvzO4Hd9/NSACh1prOQwgZ7zZsQ090a2FlR
LlyD6X/m22l7XyDAEd6KZ+LhfeHTV8uMnH51RtgSseq5uhkNRmInic+OxUUI9eescHO9ysRU5WhJ
ZC4+F77NlE4zUi2S4bWlDCof73s5+yQFWd+pFsEXvT7YPzESYGA7MmV4g/Ty+PDlAP0CRxF/bwet
I4BX8H+B/JCd56N7R5w8QzRUglc/hy7XRmNhWVn8bxZcAxjjS7oCX1hNqfEe6VRvF4JkuBr6HKdZ
GOpXZZcFZhtLr8yyZCCUT0OBBWNsDxSlK9BqJoRdWux2BpUAqCTIEzwDqwVCCNw8lppyL4hZD72d
pIXlr3NesqCvPAnkY9Ld7IyyLisZOpF2G+RgJwG+zyFrWcZitbp22+/XhcFFLFHEz6tlvQWzKJgG
DEsoAlR5nei5zBIt50zgokK+jn44qz9tHT/RAIKt02Ouo+eQ8DDJA49BLgxV8in07U7+F/oTIT3Q
prrXKflE0TkCF5b1qbiXLjbvfe47MvH37KvKrIJqT85t7/kfAQ0L3ni8nHad3jo+epwdllW+9Loi
rZs1SaES45igAQ/IvQBx7d6dJZ93dx2f1/Iik/eHTTXxvlEMYRKNdnLxjY3/O4A7fgMaTOpnfYMG
KZ3Bnc+KLawk3TmLspUHJrB+O7ItjnrSwviPYaFy9+VsaItTTKsPC4OvbpnVgverLzCKbEMLeiUm
d1VCfcwnh+WqsYX/R4XzgHrPXTFVrqHcEDMM4q6vo5YUWR/V8jxqDbmnHSKj6In9WYXxZtx7xSjV
F8LSuIZjHmc4MrX8fEGe+BhvjyvZQxFmlyBFucCmhnzdDyBsEJqeKwD3q3+BJ/qEbAN8JMdpdNwR
/zIhMomBWoKZwpqdIgMLFSqvJjSO+bQdSrHR6nOk9ZHSCLjOBU6LfsaF9nqyTxy/3EaYfHy8fQgY
hRngY0AQgVO2sq2sIJkDG1E+rx50XWPxiIMTV91dE5yueMqWpYnCFbbqU1Jk4Ddq7AlVqFU7reSo
MUGGdkM123u9KJq7NUhjk+R7v4IY61JdyZa5cL0wxz4ScK8o4XuR0/4ulYSRaEzbuHBwq6Q3JBNs
xpgXNFth7cnt1GJYCOj2BXJNfWbWGxaNipDF/q0CkbVzfEjRumpXxNpHJqOz93JDd4+moa/waryP
FD2HCN4iUjPaaMvGyzGtYBzEdzwiKpZp9FfnFgZOX9ieDChEFU9nmZK2/0nTfqAmvfgt0SXR3RC6
IcoJfEH/1zHZqZqeNn7i81pBi8OffPIOX8cttd9djsqvhQGJiydGSL/KKuRd46kwHy+Bb+ZOJ35T
BwTpCMVHNYwIxHLd1i5dWzuXXXay8aou1auJPcajTJ6waXloxhxdEl+usXQ4FgHqxvFNukzWtJ7M
7vzO1r06qTNivEhSLsunbE0hI1VZDl+kRFWQlOc1P2zzML/oHQAN9LBurGSmXkBgvY/pdqiR/GS8
uCrln/vKpmokDF7XLfxG8l8OYyjK0PMBO2/HYrTuSkPjAR4YAwZ4bfU3CxkFr6/ejzkeyI4ExU/X
5fD8PB4Drp9kWHmTb64TELw4ibjWM6Z+vHS/kYkuv2cZBOFFym+SXWA5787SP3ARWP2NQh3BQUFz
vABosqHskFYh61nPCxpeUsYWd7fQ4jSPaQcQhSB6SF5c4aNIcNDIic0soTV1SUEglnwhFHUZBgmk
pIXZjq0FBvW56Cd8KWAvBHKYJmmCTWgvYPXlPQFNhYyYIqhUkeRuFtyNPc0DxfA70bGEP8mL8dwV
WqVhjnD0DdcNFX/YsqjddGjijyiEiziq4y4E2x638zMVpisHNRXmROQWkvPcUwoS6D/RzAz5r8pK
XtVJAs9qbAN1lVtcrdsX3GCFr2YFbHUou4k9oeKhJCacLXGpKFno/e0c1l7x7kFxTtgDbY8rNE2w
A1ATAUt9XuAwdOx1zVOyGKD9cs4P747UYoi19usQvkXbq8HlM0UF0zCpblrMW3WHvnLFIJyN6iK5
aH9K0fHDqLq/kY5Chou7tT7OvOXQx6IN/PJiEjntzT6T4oQhwLTymMLzJtpYeOmtf39vgNdrcd/E
wPmz5laRb8cbDeZ7vH8AdyaDjaetk+Oi3SaI928ZR2V1ewvpHtFO0htve1GH+k+HcsOrxw5wHa6h
S0jClCKHiXrGN5CzLzKDf3Jvy1u0rpihXEF11/mjKAuJD3sq9RL/ONAcY8L/Ht9k/sbSv4oqMAxl
oob1I+toV5SBNTNc0KveuF48PXxDglC8kjpydoj9uz9sOtqkabRMCA/NKcw1yFl0v2dbcEN/rySU
n3IF96Hi43bsWfhCD+dDKiuOPTcn4DTeU9CPwRpOcYhgYflw6Jx7vep1njtL1AZiaK0a2ItC084d
mWIg9k9nC9sVcSoRfSrL5oo1ExxFdD20uxNtt9RGotrZXwwqMqYCiHC47/S1gTRbTuz5mLumZjAU
E0wZxKirSrZuGso+kP4B9ZVAeuKVxy8o4zh6AonG+ZBLzHjPEp+zWZyQTjmf/2j9ftjhkl2w0c2c
Lgt6e+ySrWPPbhnSeJwSiIxXV8kmYyToOVH8t7q6mVvL9oxrKt1R/dZjAYvRA8tW+uwP2osVVny8
u7o4qzdhcFYHociAp6Okv4gr6J8DJwysARwhHYpZFP2PkQAR3UgNB5QHMwe7sZ/qIRmnCRt+XBuu
wmmFldRlZjSGrvnPOGKF0IyJujY1+lA5gC2E4zNHr4yYSlXI5TOPjVG7ENmNWsYywEq5JNmcL6c5
VXXc0Kv5HzZA0GXO4wFdaWhzWcZBIx4xjb8BpAvTWO63/MOQTC5aS2LBs4CAOuW5jnKEl7Z6junq
m7cVFGYQScXUHRxCMGPS+6gFL8U6B7Eym1l7nBc8kyfPwalapFjhntsed1FCb+2h/0Tji5XmanVG
geANz26r31+6diZfPTm4wRvUzTKpXJVjblLqqVLdZvH55Wpb1alv/ZUOr1EvzPKWy0HSUwP21kis
KG/SekllJoUF0opZ6Od6n0+A4LxQ8nsI7O78dzDUrDgpJV2346fhVn4BaqufmFzEann6R6HtZLYt
inEKESp3ZHSXsF+yzTtVeC06u8mS7GqrbaDuDcoGCeixGFioZ0hUYeZuYmCU7u77GM/f7clHAhfW
UMRxpMVZC1OT8gWSlDZgQWTrvRFKq2UHqKPYCrHzmKMpck5G5hmazmq03XYfNEJEOhdIyjGiHg1L
+CADOdnpyabAkvqWqDykOzTT76fFc6yIxf2ebMLzCAkAdLsRzi7o9C0K0/dj/Jb5GudmoWVjimJV
xHqt7e+xb93FiBz9A78j6GzstgAoEX2Jjun6bi+fLmesZgiWD1xuEBcwunYvS/3t1exuFFBqnmLl
umgyYqpMBa0gNrM4uD9lBuakq2uJGkj4T5htOM71buUa5lgxxIq1be3w7g/W9y/bTKpfoN0UykuL
dDEVjAUxbjmmZQYqX7woxSbLQKX4pdmILCIFVpdC3cAbq/qGQT5Q25cE1terlL/urg7rhIiYBs/t
Td2iqJRE+2WBtqDTrDn0v05D7reMOLALYRr5xoJRAB3jijih2xElBacZ2Iglw5qM5i1eTeB0yUCj
Pkw5oJ5VSK+SE33XsiERWsB+bhsxyeKrRpdkMriclxByvkt/1kpwF59zEUa3XmSjQudnYKZzAo0W
xp4xJPAQ9EXy2SAVKL9UklwN9xDLJPlGQcKwgDmhm0NJEBFnqZplRfq8TJScufDC/ZCAHWoWpKQn
RypUzMh10DG19m7wiiMLqVlD+NIwIiJQLk9fcRE7WWyW9rEORzpWEeXlenWpczootQC2MdkoKuLK
sm0v3JHyR/oSpiEynmVAztyzTMk9SKUDySxCgKLPjJkZwEfsVJHmwB2O1rntVxoob6sriC0H0N5w
gN3CBEXsXPlJvlJsA/CGDjUhipCEPsQbd73bm75P9ygt9vI8zCei8MsVeJmao4UzZz1RRRuBeMlb
TUR1KpJwxFpPj2xpkZZqTtN80i/1ZYlpB2kqe7i07iSepunFOT6xczCKO9OTlv9z9649fuAJaOd1
d+M7bZiNP+5+1GLRQ3ut2EHSh0KC9gIy/JlhYqQ9AxmM+k1zpn+SxXJUAE/c9EEnCiyDLv0iMiEy
vy5z+WDNt8TRsnnygagqr7X0gwe+7QbJlodUtKWl9EcTYsFPZs9A9sxAesFQQYATEgaDDYszDLio
IQZKhlpthovDwsltcrasY9vIGLWB4EOaegpo92W+Na+Mhd5fG5oQiFHGAIk0NKx4Flv16AsAKdsg
bZ8/EorkeoZVyRoXlfYCvvS+noCEkr+xJ/RqLonWtUD10D6KL+TUd1xZJRURc1pOBnVpYu33gvjY
JxpDTQhY1chcp5V/w7dnyPn8cx2BOi0P/RPltJq4YFw5WOtl36s3x7OsmMrDwqFB8TGoAnU9iZLi
eomnZuCcUxbqnaEDC8DE0QnsApGGWzwyMuhX3srgB/uEDk5IUyKM9j6Wuq3o97CegXYUcP5+jLGA
v8ZNoELA1Q+WtAroNGNEUXjmmw4JgZlUP4/LI1H5FULDfVEys/yiAV3dE1wScwBwGNYpyqWrSoFB
csHCbUOUVobZXE5uhM23D/gFaPcKVaAMX30ui0zzQ0CfgxMR8Ii1LFIRobsZdhSu0FNaMZ7tuazt
aRIzshHncGcqitq4fNo2kKp8Qq0ajIMGkIjhj+qJwUzt2HDuS1VOeW65ZnbQ7LBh7M/ubRUzIit0
IQyFZsZVAwy+gWp9nwNqoTKB6Vc+ZYUg1PCOGtFmacoVtC6X4DancHhjtbCVs/Z1NKcTyfasDeeb
m+tyLw5t22tK10Xk10croFBe2ZvcebTJgCka+WOUqJeP0fbd6A0JGTunJKxz5P1nDYlnlwmdWWum
MdG42HUkfQIOYG6I75FHy/s48qaR7fgmrgvtaxH9k8w+Ej2gapQ1Ec/SnmJ5APXy0OjQC+tsyd2d
tvW3vklmr7f5S+mKoP0z3apvuQa/Qjlsy8kLJc5jEcV5DZ0FuH7v9PodeZJDMrmapd75zncr15w+
XE33Jv9nQNYOyo5LJgaDPwtFGX9tZ92xbiROjdA45LaSQq4op1GIGBzHjWe1iL4XRvCEocBZsRyI
n5CS5oIDHLdGUbcJlrDnJWmEO4rE2t0S18ovNrypkVn6I4mMwnlhUv0uzY0+LwNoOEJ+sVpKhM/Q
u/EtTHX0c10uMqbbhn/Xvr4Bz3cc0e/Zq9iNV/u3Inkpxewk184uYUGsDS909DRamyfxFuEpc+kc
1cd4mmIDotvYnYDFKy7uT6Ktwa30NCeEJy+oCqOQ/Y2c/0aEDboFIcVrYWmr8o2gXdFuTXbdbuJI
PGNPyC9YIcmD0b0cVUFghb9Oggv9eig8XrOY+tX1W4oZgN7fS45jF7QDCr8imjpbvxpAFxoLznrI
IAHUwsgfsFHULyhY2deAtBTVvtftrxG8rt+HEAPQv4XpfzCMUoYCW8my5m122vjS+6PIBbQo1kCV
UGOgux+83Ur3PLrpt7uw49tmgai+2Hi4lffaDTi6RoldCjqOeOkwiQtdgxjpipwWxAQOWeFhIWws
7TszKoyB3s2/P1sM/Hd3HgnzfWYB8mPb0qDiPXjgSR6SWUpz7oMPg+6kPD2QSa9Jij2nIGtIuD3X
mHUGCfVuY0efwZxSIh8Vg+6H2Ji5RBkk9MaBhLbkiT56KvH3uWuAtKv3+H1XdFNwh0pw5p+PXu52
NZQigGwyctSZWD5lWaQ4ThkadGRtKL7azyFQEw8konc7ffUs0d1yV+Akes85dewF5ydoA86xovHy
cyqNqh4wwuLyTuhUc0amOF+9A4MGx1POyb082UJMcb8MvNrTxN7RJZJ4QoWOrzkHpn8Og2NOuNh0
Uf1KUuwv0gGluMrE53gxsPTRe3nEHJEJVUKgx/JEU9Jr1WLp96MCHsB4Zr2qz65tzyOvVqzjMlyA
o7BJSbCnrUag5nLxCvHzvDfb8anDWhUe+mOO4Rsbtd5z3CDfWAbSb+YezKub5xIvNVtIVgggPivo
WLbwe2GihCxh88i1QnMczt9V+7vI3dOEtRGOg4itKQvk2aRHvOAlw4Er1hz9/XX2HRqXX1bVsIJF
ogkgNL1qW9GMFT7Y3lv+Z7BSLjR/aTf1XZeUaxPhPGsBtqw7xiGTAJ7PnQ43MZpi/m8/4ZkicsEQ
eIqV83hwyT6tukYpgjqn+mQf/tRSoJg+ar/+DXqh06YQ8j+fmO5KuKjy+cIqlZeIyBveYdBd+XSx
W26F9gxoEheZigvB7zO3H/dSKW7gyaypV0teS1xSn3HWO+2vd3WGUFyHOB5fwFirC85geFb+hD8q
3A/QskthTsmtqcqt5OUaaTjyKS7ANTQOA1nkLK+tFc6jFwzs80T0dAmio+AVhJqfBPzCL1qC4Cv1
89jkMkPXH4mJZy/7Wrrw/cJukp8qDu5mOA/fhqkfE1ZkR1gaIG/Mo5Fs2pDupsii/C4oP+TfwCem
92s0oAC5VGbMlZX24hJpdQqCKPxLrE20E4a4Ck8iIvZd80J1VLG0fhHUSdbVg1XC7dC3STLtY1vr
NAIqje3L5AT28D60zD4bhCBIiAvl3HXAT0zr9pWXjQBSEYIyLQHS9Ife1H31nacWvuQBcWi13ajN
v3eYM72Sd9TOL+79cZLTo78djzialSuRctiFOt2YXzfxFMpC0ioSRR8O1eNHFI5e1QTTaqLu6ukv
PvAb3oXcSzrU/0PssPrTq6b0zz+9QGUjlATyCobaTzb2C6c8q77rsP6v/ynUEGwrAdX04kirqLwC
lKjY5aQQ3zq9I1cHwfIoi/cNJ21KUFy5C00cQ/6aygM1M6og+MSwe+fgQYUiNLDJxFGjJYfYvumQ
WKBf2Qtn7u6L1eluJI8J7ZJOaxNuBRx/evcrX9MnBFVT9ljV+0d6bFrhT746UUwnOrqRWBIaEirt
mXDXk/puQBH0uBQvOF3IZyNB+XvgJi1OheNED6zkAoq6PJbU2/Np7P8Lu8azq5RI+VMEtjnqEkyi
7RUGAo/YEl2PGtM9bh5BIOp0Rbnwsih37TdQTZ2ThkyeCwr2S2nJVphv6zWGAUnM+8dJ8FWWN0Bv
/y9WKznCGqWwewgEXImtKjmTjc6gZZbMBbLM72/DPCZ/T8RiQ2emSDspP3Jb+TFlhvK35pHIAiia
+OYSisKgZcGOuyBLPVwpSUJRGObYX+flV76Ja+0M3TS+YclZ3ELMogiLmyUfraVowrcuoNKoFqUP
+sT3j/otxo7webBFs3VcmkoWvwKJUjCp1jz+A7xkrmnmGLTxNZAPscHR8hx5zlAEYC9ncEmOQ9fH
ca0xhOEs7bjDJ5YYO/3Coj/SJOaR5mF7wOuFGhuq08ls/cutWmibBR0O+sDjWYNjlWZuByTeNix+
JRcXVIkWMzuqglm+honWQs5YjceLP2Bxfi0mQoV57UhPkTqIufg2bAU1/rpDPOrF+FLRaMU3zsN/
7oWzYjHa0Iv9dJMHvze8jkkUsWzlO9onw7/JoV02EozyehjK1UqgrZTO6RKQqINq7CwU/uZnMpQN
ddMmvCaP52+jAQe87VuBf4ExCOwv88NWevjkpPvi3myWaPjOPL9BM+U8vxxm8895FJiAz+4lyS0e
M6OpX2862wvUk5qD3m2bwaAcUDZGrkNmkfIsD0DNXWyGDQV8U100Kh05VJlX2WPvdGM5I6S3Fxby
fu5TZxX0vz8cearZeZnOhnLNL51FOPqutVFLz3jp+Pxg+gN3VyxZkwf+tQGDyWiErZRf0+uN4AYl
d0zZdBRDvxGQ7/RoDnYXqN9gV5XfrYbmgLhaAfoBYpBNhl78j/uxP8dyt25n0dZmUn9jjpohHNea
zJh8AR0hsirrqACbj+CIvDR/yZLrhbP6vHDvajvbT2b/CixW1tYK3xpRv2+B4Y81fmZSAvvd+Uoj
XRXRXJkzzd45Jfxr+ulHUkJwOvBDzblyPG9HD1dUIHB74wP2SlWWXyN9BUCjaAj0eLtABT+67zhs
xBQ7vz8d9oXHN7VPfjvkwX/FkVsmKE9XXQHx2l/RDYfwYVftCvVS3q6AjYh/y8FxKtKZTpqFC264
XH1ie6SAioM33oEnNY6EKlj8LydRbg+JpiGS0rZiEeWll/HrXsmoxNanaTfvrmGA0xI8bEAP2g6L
iu2XgMlTJHP9PpN41BFX3HkauC9VR+OODprQnstzQBYSO6Fn0SzkSbnj4p2d876K3h1Q0g0b+TOn
FOZRTzYigSwjE/BtXwfy9TsLo35Y/iEEFbNwCE1b72iPQ2wPOtKjKYRxRxXpPUQy5vPuvEY1aKUN
Bjzbl8XKpOW4Hf4BGYzj0xB+iac+fGFGWXWtQRS5ieYACL++DfUwd9oAcMMGoX2HTaaIbgZvuHkA
NCtJLHJqppeRZMIsbXpZB2f/oBvNz6eNsjvO8qezieNxKSiWEc7y3dCDeJhPDXzjR6c65Hm8ziYB
ylWIdiqGap7+WVO47LiRjNnTNENQYpzt3ui7q9oSNGxLDlVTQlQ81z7jlhxEAfd11j2sooAEMaHi
QA2NRA8HVD1rQXjuSaScmB9lLiQlytZs8d6XOBbkekvTISFcwrk1TcBUEHuMbBmI41GZalFw7zTi
r9p8lwomFcGOPBgLaS8fWzcG1SPsvbKC7kg2RF2Gu6YwBJsICRLv/q4asTXQGrqYnvvLNSZ1AMwx
mMkYGVOEErXTZWwpJJRP1nDbP4/fdkTFzJ4oAXRnd2DvkYhpzH0J4zoE8Xc1a+XLc8vgTkFKXMK5
cO7BxLzXGT6tBfGDt9DgC510PQnXAb38muebg0cnaE5uHvBOLh8BYoyi4kfK7UFQHIjoKTSjA7ty
ERaOrJ4MOS1JSRzv1/ARfTRdZV/pISZjZhUt6vP1KTT63QUXAyAXPUvezcnP6GU0vSWIZR8XzDKY
eR/TQxJ2sDNZ5+naYfGlVtwSP3Pxp0X1nB22rWZRzGmjsozNVG80GPDdghsCCajHVGdRpdNQ+e27
gNdlYGg/dfqvSGQKBJm4lYwjLeH9Bf0HHUDeqdW+HZLfiC1mwcx2CPPhP2Pu0ikxtBOLHQBlHgVF
j7SC+aFNn00GwxhCAKgLijfe/60DXOqCW49dJ9e/jqxKnKgwTOWvUj6qcZu9PfXWguz4rsH5t2dL
yQ5DCI0vVSvZYb2Opj76//pidVDuWQni3Lx2c9BSBVZbknGQ0MSQRuCjHaiNCXRFzz0786IR7li7
d+//HMR4cSM52xYych133wQvWVjhhMvWmfTUHgtYADdTG28jjije8m1Ts+Jdl/F84OzwK6I3eCrU
lqEUfCNS8g9kYqLjU7XZP0cavkaH877kJvDVROC1jT+2YF5Llf339BK1Q6W2p9qiOhiuT1grJbiy
nVuPzjjRQ3I/PM1QZN5e7Af46rMSNoEwgKyeCPcIeHRuhGV9L1S/f33tlFHaF+iT7g1NJFXlxlhi
qdKrl7GGx5zN0nrsqzUzsEb7k4clyhUEzQOKd2pI4iE+7vgmB8i+dLItPi75h4gH2z1pFAmAo79K
c7NZkVRiUOqWHkJGSedogj96lRay2EiuVQ4dIA66n6U/f7NeqQkGHCdoW24DZn1zNz4118oF9ZLc
tHuc5NovJp2b4c0d6DT6DbcSAbFTeAcuazmOEcfMgaTyiYqWo0WaV22Mjao1J786pdFM8A9rmJoI
BJsn32b3tgPCTW5zmxmQWUjSD2ovC/SYr8rPGUeW6oqjXmAK2gLhtDk+HW5d4ZWAee8u4CF7JUbc
+6FsWcOzOKOaZaQm3VyIkeXTWTHufDUCMf6cA0pJKGGaQnWK65elT407Jbm2AueBjXECZIDJcunq
hx8FF313ZTbP7FMEip/Urg11/S6O4GyJHYExcFpB8hxO7c/QxltYfGjMwOCEjpyCJds7KM6Oozlo
Z1YZYTw6dJ7N70ivj8tjcj9bit5crzF1Ttc04T3Dls79bSpwHlbQa+RweO/WRV+6zzjRFopKXtFX
MFE98oh/sXb9lF6uCJKIVR2QKRbrWWX65E1O6+W+fENp7SbvmlIVh26H1DZIfnBV/ikqzcJGwC0h
TA0x+IlyqDqUJ7d4k+uRvBX5kIVIMzQ48z0Ii2xlQJUg/q/uyS+xen7X7N/kKpxXMCbt0QZe3p/4
zDt3ZRV/a+2Nys3/NbCAqhlzVtTANLun+KSDbJK68w46sWdbyCcpmo/3jkf0sBLeob5uFEpCw+DS
oPvtm0xLMOv/fmrbKdvBoYsZiyDY48Vq7HMN44Vsvu8vRRhhXwIskQMVxkWbaSod9BVAyeH6SbF8
kB+nEzn7pyAOQk/5r1KL4rWji4gcwc8LIygY6G5cyIjSg9cCzoy8iXIZstZtM9ia82dqWFAiWhVf
SO34yyyz++MvfmnM6yIufOP9Q/GEhiUHP48sjDWePjNG5K/sORG4sWYv15rwjpt4bGVDxWK+Qabc
CJvuj9HiYFbhgU3bC4M2z11WMoXbzZAR9Yz+gpbcA8BGMSX0uxpkbPU0ThGYs18cmr2eWH3IQagG
mPxvSBO4Mn3eDLEZbI30U1io3qx57Aft8bRz2PCT/iHgknfBNn/9gOARAjrULN/b+hBvG9dQV4Sw
n589pT70GxyAhzlHXHcNyP/3Typpiupywj2FEODmw0kjflJos3S09ZRPfUhVnAXnE78TBfTYAkQN
7NYOmish78ZqUCPdGnHScvp2hzR49i+HJMklxZLJjVzJazy99P/xUqb7lTtrIqkTr0/PdRGELVnC
TCphAKNX4RZDPAWKroVjiIeojVZ2CsGgXvIW0NolicrBs4f5zZKGpQ7zrAsyBk4KLLacfFog+XX2
j9D3v6iIZJBrAJRS+h5P0ojijjAKqvHCdET8BdNdPd0+rZu8gDz79s4LuUHvDLWUgeUawZsL5pUv
MCuEOeQUPdN+7AZcU1/1J17M880IWTDcnKSmUUpDrEgS2LfjeUOBzWPAo9h0mZLaK5o5Z1Ctvm8y
qpRm1e8k37mogD+RFRhL3EKIhIReq9etki41Q4FDUw3k5wt2sLolpq8iPk4He68yqTRiAJGtx2yk
qxOgF+omMF3KKE8ukz1BlT7N4ZxjwirPIoDfgTjIeGKxbAfeiG8oIOl+SmezCGhFYWPJ1fev1zrm
22TTQWmXPGqXXDGzASxYiw7AXnOx06OKSgxTlNEx/8mze+4DOOcRycDecoYqKYUEAroXNR/L5xLO
jlwnz5VOvu3unHN/lwDx4hxwicjL5t3D3ch2x/+fseymMNNQxFZXEPWk6AX8dqm+yBg0KSDKokIC
q7LB5zop+U8U0PuBxl2SKv/sTicqH9yAoIAZXhUgyIl2f9VF3+qf7zFbTqXPZ5k2AOZse0PAqJcn
K2gO7ETVe/8QN5gBCSZg2nlGULBCQyMblU4dzUrLEU7lI4t896/g/qeQlQ4/pGFjwnCC/T2PtRjT
ZjxFI6WrhhwGySgXuKdhuUcRS+GCrnZ/Ttvdn13xcvDmOwxo3k0Z4r/1jX7GKso5uJPHA6O8NKXU
cYQGpL0bVKJI55fFrNLQksnvsWjthHs0EiW2wUy5hbhvjbchVPvSWcyFZsvmGlsdg+i9aluZ+hpS
GBYIWyFCaQ06K2D9kwwFWfxB10z5lfA5aabZyb+cP7R3Y3y2bAGtjgRuA8PWe5qXZlU6N/sd+3PC
37T9fhR8OYNtxOgPo8nafXQW2q8zpvHvG3RudVo7t7PwIcRYpCol9abycXyY8X4XWfXqwK8gH+nF
B63m89kLMQNxe3n6Hxx+w5Xapc2nFRF203XKPLnslvlUeAKDqgbZgVwO+AhcHP+mgmfDkZEU9WM9
blf8qzuuVzhvzjyqDb2bwhnt+qFT4m5Jb7SeBYdx+jGX3EOnmpK9Qtj2wRLs0BhbIAekR2LuzrkJ
Eb4cQy40O9U6gRESr08rIQgqgT3wyFYAYBCruQ9RoShEx/4XHWtkRiyNF2K4b/iBfEB3zu9Ie55+
frgjYLzjAuBYMjGpzYeh5pruRpmGqTfuXWjFzti+eCFHRg9AYXISV94bnaJyTvw0BlIAwpyWVBsl
N2YTvR3zspOxAYXt+pqyEeuhvOoZD6sDtx2EJACiC8daECQvolsSZJ9rk9wFlm5eGrqSqRFvn+az
sKtsOFG4PRjf+yxFSWMBRAawC/KTFz/zcILzbE1XG/gjJda9zZUaV/XTJJFXJRebxPMeK5fcTOu2
DZIhYxlpAZgW+rjdg1ZSAXGwGZtBXNtmzq9DsRmnhZQeZUd9uvbPgeQUW2S9yIqaVNvaHuQmQsqt
Y+dZt+J3LlGIofBgx42yasJKtUbCRWT80Ly0IOLwHRg2q/mJxpK6Jaj9eehTdGlZAJcmKRyygStm
4vmQHTJlE+0fz3pOKPV+7WXob7cVjdcS4rr3eXsIpeLQ/O5kWNk/DanxpyH4hzJsDWEO4UCT7moD
zX1Wxo2jhlJu5CFhZom/1XntyTAWKnicTXkaBzRJk38SOFFkKUNn/iLbadNFhMwQCHIwqMEQXHMP
m6EoHttNkAwV8KGeF1fpgYyF7v7GVehymlPYlfcxhQYY5nPCoehQa3Z1JhUEvhMn/ktp+563shkQ
XWLmitRFGAEBfMtnmFzb5in09Dfp/hjIqeX4JgxIogIzSiFEKyl29KUd9R0vStIiSj7cKilMw1EH
DUaSTd/qg/L+0ta4zzZumJ0AVwR7sPKjx4xWFSbZb6xqFSBqecSQLzkd3GkVNaHU7ygmCD5gCd15
gsC27t9zyG4qsmNabFYWpaX5LJ2xm5lRrBgOd60kJcx6PQmQ5wncg4qvvdBs5JgLaK9dmsHd050u
hr14B2rIL8ix57jbNunNCKyXtUjtESypodIJRksUCnR2BhPNDwOA/go0MTSkxtA8PzpYGwTz68Ee
TE8iYTm549mdQ+T7Rh7RXJgRnjEG1ijN+LuMDRhMrL5RdiiZN9uOgA3mJsTkNvuHWzoynmbZVQlu
Dp9mGYe+RpkvnNdPJmXn85cl5Jie4LLkRNQgmbyI566aJmpKQtJX5P3rsJiJcrC2+COpIOfHQfSH
/byOnoZk16LfrFCTkRpZFgvzJl17EPN8B/EcUXw6S7GLZm0ci4wEPiofSNerbMoZDbWQF5uI+YO8
9t6Dr97VaUZ4Q8PWIJgyZ6WwBJ1rIboz7snKwvUK1nlR9npfbr7dWxiyv5IFZVApz8mNRTI/0B1I
5k9Z71oeVGvI1xAk6hAOV/RKr/OizP5diyrd+PQ08tFHa3XWrwc75yXRZhqhLfEL24WU3ah341NK
m4ZNCOeWmrU6EipMgBvYgCQ1u8uodwUroF53RaMUxtmxHFpAe8XRCp7G6OYL2VLiaSK+5krqA199
hBdnD+LR3/VkLxx2iv3OcxhvYvT3MGuN17sKTCojROVPn3/h/NOT90L/Odbxbl7I8MN1X9BmYnRB
Yb1oGwdcx5c2qdMM0wXbQ1TKp+nT1iwCMGxDU2xqU9nNPKz638Rs60ifoJZ9lh8lxpZHht/rnXIn
vhui/vNrUSnJqz1Y4bHI4mKrL+Ihc/pnYbS1uel5e46jewi9PkqFsNH4qxN8u5163SuJKZm2pvJl
g8LPJmwuZ43yHcQErPQF6MlGfOC369NWY9/45am79ABRZhkIxcBOH9V2ri5GxWxbNCyBy/AYknAY
HAXY3Xt3LAKqyDUiYeowzTfBMikSbbP9zkZN84fwy66AOwHaM1UftntiJ75FschW8T0ZOicqqHLv
abqYoiM+f8Z3+Y4BP2MF3J5O2iQYOC9SXIJ36rMMOqvX/u6lzJrjclMcotPTXW9Vl/UogJqbM/DM
yvih0oQc7+flXmeEvwngrOoxSEgD7lzb0VupkuTcDh0NrRICVTDXYZosIOF46nkeXPt+iepCcG5Q
67fBphDmZQ/4Adn1gyhSDKU1HSzSxO4RkaRjpq3/yxcbiLMOwefC7Yt8W/1DqopkhGTw6ilEU2Ff
71ztPtIF7J/K3eExLp7XUZuORKGSsj/hsf4D1n6jiAyF8LmZvxfeQmOBvPQ/4qgzz5lmZHJzWnrS
+teYhNZRy+J0ywGcYFWWeRzGtzSTmWchx/A1paza4eBhHT5h6ClHu/ldW/vO4Bcgin/tIGBwxHE5
SlzlookoYLeNyQp2N3SdxUpxBdubSRMNYGnb2tcrq3/QiVPymjT073tEwkHURvfTeTkE3ILhP6MX
lM8bxuqUdjC9q0TmbDwXRVYboo1P9PS1Hd1IHcwetwFa1SjWZ0SohFDS4vGGUjvGFumEuwgRej7E
QGcsCnQxIqO76l7ahdyQz2ATg/qKU7DXvPuukaTrSkMQrvVCU0biu0xIPQQ+Dmz1DJk4ZDZf7zuL
30JRi5PZxL34KZvsJwxca8s6nLNDH2hPD6A5fngo4RiyfMHqcPpTY0s2q2vF/7IjlahzaiWAXjSo
dxoneQ6AVq6196yPYGO5mlAn0r5Rgde1hZcRImu/lHsLsVfLr0O2oM8yyQZm481WgxUyekoF5jJF
FXdQM7wRd7lARIiL46D4wkGQ2Je69DQpXyxwKMshdrYA81jxyXbE7G0rVQPUDDX+Rp6QN/BA+cnw
qUctJbRR3Lm/27wb7zfoCkHDgXt1bw3OsxLA8C5SGbc5ao+VOQ9L50CTwvcMyRZL9hRw0syA9B8B
S3/96PG5rELJvnnv4jjcyacw7xUZwPDO9F3CxD6XUS+utqqnAkxUU9k5zz3CUKuMrnkX9p4Y18AK
Zi/NplCjvSIprWtoQ7FBbPJnJYkC8+oZbA++KaH1jRME6sY7w2WT5AIdAf+mFuVFN7e3Pac3v9Sb
DldozzpeqkS13/bcEWB+uN4Crt7h76hJfdqWa6Y/5IofxTGr1UcPz2mXbV9J3SpIlgch6oJQWl95
eLir6gh6fWqgDpjV0RBXTUZC+r9XfuzsJrRY8K6XkkrzNLMdTt8vMvoKc6kqvS9KvzpDZNhf8x7F
XXdGL7V6fYf52DMLjmUlfJkmP0WwENlI4hHoXUGW/Pjkr+tY3IMpyeWWtAAO5hduOzaNa+usCN7s
ufiXrkm2HPTtyv9ouW36l008dIXNvPVbJ2TCAfyekgG5+Mr26RAuAprCEMCmNSFOY5ytkUXu+i48
jxYzNwX2B+QlBFshBd/VbzQmJPK/DjhIeVOBtawT0zE6S428AFMOLmmh4ksBE6snX/cJmmUe0TU+
xagfcF5iQnseInVOC5JulCV/YbJiwino7LnE7Q/R3pAPQYfbNljMfTAvJkLkSAucOD6r2gudwLOo
riQFRG4rqGSI3dC/4hDFiFdBF82QpIg0H63aTTbLf+fLEsZP+JxgpAvP/AQul29hAyCjV1Q9+zf3
jcHBqqSwbojFtWdWiQAc4uDbM0dgav6Mxaqyg1tOObArDDfT1Bqu9UWVy5pS/bNxRhdrahMzTerk
ZrLgbF8NRMVykeSjecIv0/1v2qodiWlXEtr9eIbGsLHewGHoZHam+qkkfUZjw646u7tL9raYML7J
0gvylxUMCBWD9jsF2yqXDvhqctrPr/bz3aUKpt8uLOgkg3lC2fLOy21+iyCNEUT89W2bwyemDW/y
vqm+s/7vMwLumDqZ62HV8IdQLXp+CHB6UL9XXagnfHHc+lUV6iFyAS3a/J3lbW4c/Da7L+Sj5DxI
lGJUMc8wcOU5xOVZL1uVdo96PIVdfmWOQPTsIgd2k0pXCkP3DoP1OglmaT8P3jXZ87u6WToQDhV7
eSvF22/SzlBWRt1cgYlkv6SsZ1Y+fzDWQhw//QOd6tVfvc/976b54CZhE2cfPndFcM98EY2Pmg5W
stVvZpBzi5AiqLgPQtkSo16oguWab/HGF6zect8oS8PjucFV4m4aAMYzJt1AhFk8f03MRQXVl65X
wh6fd5h4Jw/OxHjVPsh/+VC0OzFAtg2wiAptc10U3QV49sorYR0viLliIBit9BvOE2o+gJJxeNrt
C+kwKaee5ZMGmD1LexFJ/Wi5BQIBAMNbh+j0HrdsSVyN1yTGh0Ap29oa7BnV3ik8b6qN4OYVsv1y
UPZK8H6nsiUd1m6WZ5I3/aCwqvCWZKr0WzH0/Z1gnN4sDTvSW7UeU3SSZtjHUiuwUHIUBDh71Coc
/FV5FTo4RJpvZbgxr0L2lcaopJ3rGfpXF2eR/sH4MJdyAPpDCtYu8oHQNYpCFaUzz2DS9JMB7j0r
vGupsE+3tgYCMQtb82jUiUcAOBT8pA9J+ED7hH/BnKKpDfsY8pqJOdutizaXRhEvlao9rsK49Pna
JTLAvd2tg3Ac30+mBfQCx3et8sgtamkFNGeBNIBzJevFE4rJwN+U24XGkXV6lPWBmpt30S/NE3OL
ObH/RPoWtQL+a1JZUVDeZ2vpV6owC+nX3pnukbJ3RP9E/2eOwHyiryybpupOGgnclfSlqc2238U5
awR+4YYYoDlmfNv6rkqf02vS+ElMNBvIxtuKgoo1Oco1LOqWM1uEh+CHWN5z5UWbpXixkquJ1Jhf
JUmFIAcwUoBNqk6ZKKwplMcdI/VFlg3g/I+8TRhk2OwxeP6n2ZAy0z1FmNwaf9dZcIetzuAZuMr3
q9qsEFgpE+0RQuId27xnpF1Oq8VYVq6tYy+mivbhuG4yNUA1d9NEJb/GkGOksX85sKTgs55sSdki
qmeYSjAo9I0VzQzGXAjVw2jGG3pDsFplqgL2km+hB/dTJDykU1i42cx1ilSVop4RU8xY+Xt0KZ0D
LbsLD8wz6+8U90Nuk5yK//vfpj7aR4M6yRogZR3d8QB0vh4SEg/Z1NBvRrV4gW1uRqMVtQ+3iwp4
1iwrXB5jmCLMV8dCFQc0ZajLrqhsVgFAVfJQdcuwZVsM5D/p0gmbjL1haJGzYlwUDKE6IXysWbps
uABZQ2nO8Vm5nTN4PY3B8OqWSiQRTpntcOKuRY9aiY7JmcRuE+MkwHio4dQC6KqFGzycmtIblYoU
sHYriGJRHw7p9mGCLBO3G/zmNtBbTqb/lppdR1Z5vkdqn8V7NFgqN1GbLs5CPRHjKRxe7v7khNT8
4K43lRdZdtGQq79N9sSgKNyyMWd6b1n65hMRdmYVhuXB2ZyWMgdyCc7PGTq4cVzdPWU4CBITzrWr
4tDHD7F0mxTNQdqCSkhojeCBe3/KbOdbHXhjBgq20ynxR/fWdz4HfM/C64OQS7RYGsB0gscxNosn
yNe+X7WNIsac1KDFjLC124RS1Mo72DIQpRp2sZSbX7PhJbhGEYcjKw7v3Nx1eRROD8rFdHF+4zF9
WBew+hNN/MTo+UoKR/9q5Li1hUpLLE+VL08r6opue+03shthjm0jeP7xkFpU/4cch3BnNhNbAnA9
6HCfwcHcKKe76YWA0NmSvblOE7ItvpdY91jYvmckZgRXXt8OJqkahkUfDps0mgUKVqSdKS+93q8S
phG4aaE51Af6PWtf5j8Y6CLQMj/AcubM30QS9/BiWh2XRaP6eX43PZwWSWFYPeKuzmyF+a3cdPjm
lp9GiUwBhCFiMrw6MaRtIyJBKkakublgLxhwwMUuYzQtwaUgoFlG1dMH6Xb8qmQVW4TYwBBLi53s
CSM/rDRLpVUmnEKISTXviqStTIrRdoBvhy/1GXlO4+3CV6w0I1BdZ+4Xf4UlPP0IZqShWBw/qMkE
vx6CFPUlujPS2OxWt505LcBpLz4dpMr6r7evuCFbzqXO0lVPx6K4DAt1dVknpPaIecgzVMYqCZdi
yCJqfQFZekXlvWgkx2NXAoJA+9/3l01TZXK3w5j1aj6txFDt7ZwY/k6lV374UM9uKLcszTYN9Kon
G3/YQUqkUAinTAQyjB7p8YTdjd5mJZQ7msn+HNA/EIm1zM0wV26JQDLkrIH9Ct8u3Zz4Ubt12VRQ
DvlVD9B+bX1sQZr6c8NjYjo8a6WY6ZSjsZn4ELbw4d5/B9h+YA4o+fez8khlCMNJgmF4oe31wLd5
LZ2ALbDg8oR22SGwZmzhjDrf23baA5roL90kcTRtpieCFmQkVx1Ic0fkzinzmseF2LS5zLE3SH9J
pgB0Ynrq2eDnWL8dAS6iC2QEOR4s6BgE5kTRuVIlVcCuLs87GVqYKIe6mAma/Ea/IBoU4PenyW2x
tdjAYGkG6JVryg9IzjfTootm5S1YHvHO86B51720EAv/s6jNTU5DGVuPxRYcY80CtDWnQiSXFAyb
yzIdgIE902QHxM+C0PU8AC8mni20EGnUJGwaqppdKlN2YMtyLtXi9nX8VYHz0cRJgIw+5jzFtByW
gYtlPtSYNlWEf9tVmopMy0oHSQI+zvzK2zF1PZbohoI8E4dSIELJMVr44tJjMkchmJ84oh+cBX/K
+cONo+ZKDEuBNn4ElRfxd/aIlxRYl3MdAfWisPeJPQNOkvdt94bKQK8IAwDeSCOof1k9hLHuwHoy
VK8cWsHAbJIH/NTjPqu2F7/xpJ+Nl76bpGzQBrhoenTJZnogO0GLvQZjAkjGlzbXQdtVYxMqiiJl
yZG7fFx/lSA5xrxwL7BXAzWDALmxZ4hdzBGLuFApkw6cl0xbBSmC5pyIiTxj4slDl+PbBB9VmLLH
X9pCmknLfRDaTzMupdYt1Bu+R5zbQ6NYVdBv+Gr4G8ZCWVyX91n8rrOBR/QdeTYUofLvuHRofWDd
a04n5rLtOGxUsIAxYbCXPNHLaYtF1dkRJXfDEKJZ4V+K0PH5A7qnXk7XofnxpeiZ5yA+qcYi40Mu
torXa4aX87xaou6J38C90z3ZUREvM1hm1Ia1WAgt7yq7ZIsA+WaINGr++00g0RUvaAQetMhB8pDk
mOn2opX1m0fZ7Cg2g1TQjVHc2IxgoNzdpvwPTV1BTB2i4qJnBUBN6eJ4EPh4aqJqA+ZyS5RTz69F
qn+CUN7v5ca4m8IV437f9pchxP2et/bu241cNhEEchvk8RFRpaHpbSpmSKPtf3uoh5DQSNaBo2lZ
Rk8GNNreOYIeRxL680aBF5YcHeRFmGS2y33+neqnnotBKJoSxyvHxt8EKDkfsZG7S+oromawK3dg
qmDxzA9Oh+j4QlKWBXigsfgvyxonvCubdrs9N/Is9Tijid1MBjFDaUk5aDvSkkoyiyzV9pSUAI65
ham+2ENcs9TeIzc6/VgGT4FMe9QzsEaYfGP99C3OUjiYoHut5F06zq/mcG87a2ZoDF22Qxhi3kW4
7bDfdhf8l1Z/6qPJ8NlviSiyYGu5ddSXVyuVQcTmJSwD2bQbfjY8PlftIvgwfMZ56YEzh2KwC5AB
clX5UyjJwcC8EcaGXdoD7s8HG6zLIo3nxEbTP+dRe596FmWsgVji4hWHrhse4CRWpFt1VdtnzMMy
aWLUUrbkkoGWUTUGXwhWCBWgLZsn8v6067WP1z5uETeC6yS39nWGZtVqsyyvdEwPbEAj9QG574zU
GjhKDYInJjwtAtIS6AB4fgRU5Mf2lGcmGygxxDeZcU3Qpzke9LBTRKJgt7RIz2dF/KZSvBrRB++H
rVQqWTrwv0zs97VDNzYuxzaoZ+Bcp+ut+qN2kuzJJk384LtwssXMdEbWpuCQMDnzJwVsVdp9bTLI
DCAeQG686sl/74Y0Awv4CDZ0+tOj7mXdhu0Irj+HQOk7S9jD/dOZ1tT77QmYk9L4ANwsinPgUVur
u2c6v3kAbuBV3Ioox2q0cTDIRbP5hsFPekobbDXnxA1IeMz6xwbFKhXYQqIobh8kJgHNUF9lzapA
AmQRdsxEU4DHig0InCevatcvyn347RDlTdBVDtXA0GdF2Qgaq+v921zbNU9rLsrHXDLh2YmYyYxL
StEdnlpVMK0SSoVGoEW7pvLYAJUZyIuJxq0yF3UUZZN/JYRSW0Pl5VOEXbX9MhDywJWAjhO0+A+N
Nio62Ow8YM2ksjO3StHfY9xd4QljEsdo2LhAZb1dEEli6cUzCKlE20/lUb7gXrNzLtzYaKwuG+yI
xD/6i/g5HZsKHDIHitno8i+l3RS/LN59Izz7vgb+BbJhITyP76vhi6LSPu4rmB+lLc83zmdZ9eaq
Vf+WtEbkQYFX+12TslFuChXrnLrDCl+1aSENiwXB1I6aRG/EwuY4FafayAcKNSdM/z1GJ2iExRMQ
uznvwrwF36uJJGDIThUssRmlSQ94wbju6u6kjYJZ6mUhDRIR+fI41ZGa8v46VCrFFvfKuazPGAbi
mFgTfkGHgV0O3Qa4imyyL2mBysDVxt+NNHwsT5JOML3nzMA6SG4bFC6ABDKzP8q5fP/lxC4XYtu5
wiRfCX8jqxsohXnC0ZbY6UUPTH05kSoqn7hVrcg/8wf97UjRKwbUG3IMp1hbknV1GOp2m1qexKlr
1d/Nj+pnXIAnKKkWrXKTw9t5fd0cFAguDVSBtsEROh9GW8HBwXvagnLAdsGVAzyvdZA6IAQ7H4fL
+zd2E9FB4wWmO4A6blwHFO/Sy24lni/btz1yfPsZGacj5EcrhYWJTkmRhCdVTQNNgmRzPK4eWSpM
WQ9K0smuOOqfsZ6Myp5YuAVuW5/mEj057i6/XBf3wwYbktum5QjcMXQ5LHlpdbmbP/zfM4uTFjli
b6d3G9XTCoqEoB5LiFy83xx4hLIf7R/VzPCdBNzz6wPvQ0HVV7NMS9hCP9XoSEN2Qv7hEcoTadJU
0A0NZV+NFeTwQaixGXTyt2ByjGA0JddrjB3iTjnHZ903xRD0+D/gzenRovUQYuhV7UeZlLePpqLT
C4dH7TQNNTpIBlWYlJOjWk1yDzVRNIZO7mRAbps5qwPk27tAIlhsO/2vFaGDPhPtmZ7ro8E3if8a
ZxTIqH2U2FAw9NjNcXfDBp+3o9rUmiHTMc7Y3o+WpGRfqrKhtMnPh2PxTkvbGFaE5V4rQA+irht4
aEqwi/qneEAPVMSeD01qw+1nAKR1C+5fJohAMuYYoRXUS849OCpmwIeccXlKlzQ3EpjY0ec7yYVx
448hyQmVb++PaYk4ZhoSJvLV+/+DD16ZgPtnccxe6xzSrAx23uQ0An+ANr88mnH5riwesgL08wvQ
m7S9W3cFdfgvUs7R2DhXtY8AXRC/pXIsJIOuRfYOH9JgHh/qN6Nqi26/C0ypSoSKyoXhUEYUEvmD
9Nv8/rZzAI6e3LKhLGhKFQNjsg9KduNsXEkvAt6/VDR/2yRVrhOP9WKrZe62WxJ0g77m5rKirkHV
zh83sJd01TYUNtpCTUsRddqBboPA/1pR1OjvbbuHPwz2JWFVokxbiNcEcz/LqVI7eQ8yWm8rYriX
isJLLNh8UZnk4RweaskZA2SuoJmQXjU6vX/UhXoeD//aGFI0YhIsRoWwR+WjAQ0G9aOuLsKMLCo8
Tx3HyQa0Ttr8uAl1Ftu3UKoaBt0n7wNfyuOL3A9jtPhMeGRWEZiUgpjCMp4UMiU9S9sXiaDryvpF
7rI1GAqn18bmGIiczEM1/FL8fSPEovoObgKg8b8nsMQSSs2eGrUDLAUj076MzFzYk20rqJA9exMQ
+rD9bgTPt3ZbMZ4UbaaDAvf6UomO91DG7WmMUcSQi09aM8/Vvy+tzdGYJpXt7YdxtDjWHoAyNs69
+n5JwppX+GqSe4XY5p5upj2/0s8BJHj8Ja3EKTyANcZGadd2Gk7oadP67ZBFm/SP5OtvkN9hydHV
pPaJIX5ndw4lytXgnqdAAqAmtRhYNqx6ykq/i7ML1jGx/YXYfPWwgsISTZPClPDobEU/ECyWrOpq
tjslR9/jfzPqyHftJWGSVSUKuwCpgy8fWA5bscx81d4jwhwSnW263lztPVrRqC5Dysalev9iXGl5
OaTh86JVMytXMkRJQWQL1oT3Eo4jXPY5HOq+ZGW5j4ZiivCpzQRwwDA90mC4jgzK9q4cFodnx4E9
/nX0rf5EEyoZGMB5QCexOUD5KLQRd2ShBhts9OzVDmIVRNayeAMUv8isYN7MtZFu276oGo1UISNH
S/sXaUscq9C7rCxtuZDgnA/oK8iTczX+PB5r7qdP6vxkIXtk2PIEaLwGAOuhb0i7aTTabPEivzmB
wXU7tbNQnDBlSOxRPirzr/tmBv20t22u7ZWe/GoiBYg0cCAvt5TE8ZeFSa+4pHd7N645ByZt+UNi
g2P99xQInMrFyYaJxWjQj9rD5q4f72VcGKfT5YK++vHxGh+w+RomuzF04qKn1490pqDHmngMBlW4
ZZ3C8WZ8bZZ4pyWlyCiZevSEpSBfiG34dhhnGOHA8pHuEW84SfkWk6L2vz2V5WQGqLj84j3hplRW
CDkil+u9sNexdX+dfgeh3TDwJe1T26P+UbNkbKF6XKJ2yQZeEkA1kgvN0U0n8duLkJoyBTghiFdF
mynfYIfimQ6JHN4TEFLvEL+MYLu9W8qVGnMpMPPR+JDjQjyQ4lt9iApi3gLDqN0ypviOpY+kNiGe
4ozazZ4M5XJhmAMNKMxpt9ECMuUJN2kOMSw0YOu5NyKv02j549CyEQvjLJogql2HmeOfaKwZ+751
9FbSco0wwpbE+m8l6azRXrEzZ2bGlzsUy+H5Smec0II6grARJStPlqUXZ8NCTz1x5cl/K4kvkQyb
claCwNCYPcs3cYnef+VSAQ20q1yNmanZfltWBeA1z1PLuqbya/ov3vPzb1gnLA6vBEltPQD49fk3
Akr5SCTMTNulBkEjTKA0yOFrrLqovqkjAj54pacdMZROTGRZUN3X4boXq1mjX5WlQqPoRwt0ceJN
bNpSpyVoGW0CzA7OR8/zyum/KJBlunv4s0UFfoGtdYnUyX48O9dvvJ08yi7SzRHb8DFkTe9AtOg2
6mneTS1jMqKkzBPZ0mhG6jBe5Bu2Wv+y4wowJw0jssTrRM3QMJ8XGdlsrVbuwOgjQ3E4/HK0bHkZ
QkUYqmgxt9pw5dWgXVe3KjpjJ4AMi0d3Mhea0NfBTQlBI+JgNWAYU+0cEDI/5U3xVqiBffDN+DDa
F5C7nldOeRINeRt5x/Ldbpq7UPutNBwJUEa7fsOgrnGBLvubaDLKC3fcuG8/b1o3VzrAoXkCN95h
1WW6eREqsCMhjmBfl2Q30/qvyN+RKacFf55n81eDqRuHyGnw1piyRMw/CC1psh9RR5i1SnL6v5cp
l7pmjB1XK3NWL+ZtJu5OXqxsIM7xOWJ0vYV7HJwmxiwDQwBRTfxiYHDs8lrI1GyMLrQfV8TFlZ4f
E77vFe+yVLi03c0JC84jqwNZnOI3TLimclm6pWMz68muUJKkA/qutR+fsLv4UiPT8xNi7BtFS70x
T3Fax4ya97jN3VhWJrc8GYCdk2BFOJ9LwxzNK+E7U1FD3cyn2XUuFiwwMNTLFeENeCmsxrzr6AZd
X57HO32ExR4B2LGyqm5az1GLVuo7npFM1yXNquh2KK2y87b+nr/yAwA+la4OaxP2iXz5D6sRnZ0/
Y0agk2cLpN8y31luvGrnFKEcTHVIboYUkdXG3MtVcsiu5EPlPTwiEopsG5PY0bBUBdefb1sbEYTM
TqLalC92sAFZ+XKao8WDqkjdIw7jkHx7nrsFb75YHxfEomGDzrOP4l/yZx7nFYJIRkTFYHViZrgL
wtItlhUjbeIk6YvvDzYSGW22l2IrwNg82mv6evM748qPP3AQX7lqaNNX766Xaoloq4qZ/y8zw97h
k0R+Bw4hZYgyJwNDTTDtRh3kZ9t0URcTnI+tx4nTn6i0VnhsEG251TBWMsEm82+irEZinlYA3zvg
OMXKsoz1Y9cN8dApYYZfL8TThbZc65XAkau40PDN55+sGrteUn5XEuORGJJLSvUGQAiicsTurduD
JMJEkh5LGNPhtrzfQbCJ04gANZNNWqZUgayxsHUpXkhtjw23iSz4jXAhUTlYsAi7yJkagYMHgPvo
0iyF1ejseKHtjSaETXSHjpbQ8Nb0Aunko9Imw1vaHrLzIr2FVzVuQc+hyHTfgP5Y2u8KkQ7PbTYz
ScbOnMgWtptxiN8YYp2bwZitwJdAi3ZP2cu1dzgq7rfTuWhOb+N3vwPWM25bqvWVvReaKjlSs5Kl
HIpnr/C50QMARG6pLVf+Jt90GqavLYuKTobZC6Fms2JDn6yrCvBQOQtvQIsUfrzpcynSIrQE7Rx6
jUL2PnlGqDmgfUAnfEIqzJUWAD2RuNBMNuVajN/AFV/vb1TMEJOxSSQlzW8qE5E5uM60COkYp5TO
YzeuBBWf+k2NbdLx/EZUMMLTAKthETpSteV8nQbT5p0Lyx9EiVp8jvqTfiMcNgW/Wc3SXb18xnFe
33CmEzrXvETbqJiqB3XTwVcK1HbFcmq86znYX4Hlc7fPialYburWDzfpE4vZZuNkz0LBThNZZo3k
b/vWlHV1xQQ5Hozwkx3gTzkho7Fqa8Vb19ca460dVnaHDCVvQX/7TCN1tp4QMMfWxlDP9K/Q2Z/3
WkQ+rVYU7jU1jBxVEMbyRFYhHIQ36m2fucV4iG36In2T9XCqQ5HE3o8MZ/J7Ca18hFcDV2w67wWG
pmeqakbNcBa66YzHx1CrsYzaR9Sx3e0Evh/VCHCtrNaJvViKcmOnlZu6BSZLMmzBMAFIKZFWUO9j
1zNgkoKNz3POCw5sRuucZTzwIvb81uKyv/trU36xFdHW4qmWhW+b9K2cEubDtxX6fFO7RRy658X4
jUUoPhsbKwKbL5GVZa+6OhrLzi9kP4nmqRi/Lu0q7WSmdmLebdzUF3g8CQu/OlGHP3Shl36nnRYz
Kzo615e2r4m9vwENyGkB9XAwBBu310G1br5sZuv5m5SUM3CWzqUT2yApEIWXwlspWWbYrpmYFD2C
bB8xqRVgh/IehsjmdlA3FsTYGKHzM3/OmFdJcCVo6afSfMnIkPj7pmzORGui3eVvCb9hZZN9seC5
8mt7T0s12o0c/ObaVD/6d6ChhZMfKYZayRlNaBNnIBFSzLRnE3luwXNh0C27Dr2tyLec17lPe1CF
eA/zm6E7/zCJ1+t27PY4jxKUvDg1ZE1FPtTrVSFCsmEcuo/Cs48jtI6eu7A0l16iePXAE7++1dyj
7ia6OfIr+cvNdrOE42jkXNKrrUPqL3RD3gs+g0volrtFHCvr++m5cQLoUivuUFrcZrkuu+yHdT4/
Xy0ECVRFRKuoP2AlvgJPyiVv58ncgCRAI7C5LpoPc4qND72wQbuKjDdwyNxI7WpvSx3HKMXS7l2H
Gb/b8yKU4YjoeGDnk2151mggd8oF9tZKWaymAX1OTqnA14FTu50Ucz7R+Ek40s/lXpuYp0j/Jwhw
zcpQv5O15Iat25NZ9t0VJ9TX6d9OaHX5IB98Jd2ybMV1V0aaHOjfO2HcJ91IDGL3Au8TubM+d2OP
5w4uyPRFukSIDAskBoVcVLVfzgDGjTjh0gSdCbfrcsa1zKZkScOODEc8nZR18qJBdF6Ji1N1J9Tu
u5c6wRbKy9BpZl2SIM1IzNr1lqp4oUaA0+T08A7Wa3bXtga1mNKgF3K5AIAMflF8VL3tRjcaW4hD
Wt31wK+QaWMTIUw74F3buGrADd0a3ZJNHa21v9QZAvUmWudZ4ZovTmyglXOh76G6Aqa6Phf8aCuq
IPNtJ8r7oPz6gEFBQ01DYLLV8kkWk81nxYhh1Frapmi7P0Aga7L8QmiohNbxnS2aXiFvZ6O8G+n6
3+kEwQKqWAK3DYAVEpZLO9mVp4t3WjzPftM1Nga03SrsxQeQE+jUBIW7ArkPS9BmHVN93hrrJcZT
+/EkpFV4lRVuC6IMhtmyaQv1Z3Vxenh1py58UkVt3ACJxvCzsMJSI165VBKvcii5x/XwmSIJ0UD1
T9yd0iT85VUaJanbB0u5ov4XVLqV0V96ASdQcg+Of7CoEyodZe8LtcI5WguSVdcPwh/lwUp8UldX
1TD9WS1A9cNB6sALey7GNMlqMk12fqjVcekCCzMYk1MIoRR56X8moqNBqrJqAaGHXl/IrNDKEazG
0PCyQe94DwagBtGiyWi68TJSe6NJWvWXRy2Y55tmz+YsdB9wa4rKO48HdYphQRG9CrB5C6ZJdVk4
GnhWURLIlKIuocyPXh9Ml0g2kDJritVEt4htnHk4vXml1jkp2cJ2srm8q4z6tdLX8lZTWgVSYHu8
+jo+6JFGy/smpnMC7F5CiESUpKo7EKC1THv0oKSKppNQvzaaRjNGITw87H4z6QRukiu3afVA6XpT
tHborqlbDxQ1xpBkzUhFbnKYq58baElu+080QVocx2D19fL/bq5N56aSoEuD0ClZzLztVuDBDyV2
s2tMIzmmtwdvU/1LFTgmYqFomBHHzR2eIJs2H4k9L6uwBhBhy5w7LN47Y32DJlcdPvJowWCouADf
IBSSV98W7B/jibKDcxaSC7LB4PDtogJEinF2pkcxyyvlqtjXDfBCcNQuUsLik2OaE/tlR8TKU+kt
uWgKICwD04lWHGppFX9dmbd6YBczsW+zjGDdadF5kYxIYgq1/saE6WibxekoCuaiTW2cOCv4HR5C
7DWYDeHHB0KoocbdzH1/+cIK1hKC7PxlAJoQQ8E8s+4tZbi1N2UUZZywMPB5eG0ptbvXB8xEN+lq
jJe0sxhdjzC/UOrU7D4Ar8j1QfcsKXgobb2k1QcSaDtYH3v9oeqwEyiO/jgbvBYmxt5v30drv5PB
eIRX/WI6Xfj57/JCKtbYyDUFWribhGskDoV5IFm7W2s7Mh34siYzqfNMpyR+uxukIwPy/3b8hheR
+e7dBXaRggXH4i71LLgVR4biSmHAtDTlsVYBcfhDCluaq5Oi9rz6q2W5SJD1s1CRj62P1ljX1kst
euXljx6FjUwq48/NIh1uCqrIUu6KJ7tdcnd7BLN6mvD+tEpVwvxuHrvsoD5ydBb/4sSMQtsSDd81
QqSbEMzsfNA4/4WExSPOURXX3/kWPbsfMi4Di/T/GN1bP5fBBbwt2AP2HcxlxbpTgCsElPfUESfd
hjT1UTTjOpICAqcoaRE5yuRjBN8NlE0dmjGbmkBhsV6koS0y1YijgBG40aPWjBs/yHFPdDjc8QyV
bSF2HQt+VTpruHGbymrhb3eTJJq8XNDo5+5m1/R9FHgqGTUrDnTMe/ll+eesGPUA8ly/7HOo158/
9JuQunxJmkEUfo4Tsq01LkJtLmGpmSX3T3I3lmPujh4FH7wHiZonvMhA+DNUT/8r2Ko0mMHEamMG
HDOTSz+Wlo+UBQttA0QsmkrOfuQnEeYxNLBsES81Pf4yfiVKs/7mxH55fmQ6ywmAFwpADvuQ64bG
q6VWO2Y2fpEVUrXcpfhEqIZ5Shk3bX8q69tOlG+E5pQAZ8OOJswxiILHJ40eRzLYfOo5tbqIhC4M
Dq2ge5Lc5fUWbLSrczigyWhYvF41b51Q76BbmekYmFsosACsv/kRtda91GC4JySl/6mLzOwM1cMk
L+xbzzL2y8ZtmODAX4+rc7nyQsldNizekKuC9uIoWxsoEtokEZBri7OOcJ6BuKYYf16ZIcHhXqie
cCGEqegQTz0boL2Zy0Ji6+eUQL3W8mGui0kYMhyBmkWxs5h4UID7hW7TCso7g089yTmhx42NoEl2
zdoCLtM0QB+tt0FTcbA+gUNoFacMkv8LgfzlzVEecsrKJvw+9t2Gk0QNIZ7A4ZzZ02vZnyGOCP0D
W873wyW09i4Jj3gApZP1rX8XmwTDOt9wbXtpgFmPqNSnG6cRHVgedQt1v9P0LH84a/crIG0pP0WH
raHTjx3eBcValzSQ0AFoCWtyD2AsV+UVpWjpfQvtqqLjvMBMkP5U6MaAX+n6VKxMy+BIiISA4doj
MB1/lR15LTIXp4tOtGwPXz4oP29cSAuqMypfqw96hPDzeCYKk3QDJs1o0T+Csi2uAT7gg1iUUwph
5nyAPZOKgy5Hq+RQnbLJtJDNi1MIPb4UKhbHlAN5XkOECS0mKdkLi4JMv15q7Pg+0AKqdoltSu1w
MEBigB01oKq3Ua/yYvD5s3zIfCbhCLE1BzXvV9MbQA/tkYP2sana8mGZKQamLr1p0Ll3Vwm9d0jN
ZXy7XSfNwlhd4Cw+sBZYvb9nrBYsX6esQ8iEY9BAaK5ryo3WTsm2hwGc2dmK49CavmREcncGQbMU
z08gEExq9jbI6Ud975REMQ4kvd/RiPPPGzg9TOEpXoRVZnB5sNladCuWI8iLmSrDv/u0tJpuQCJX
k8JbPaYVLoUIkK96GWt+8k3xFcXtBcTQrWqpJyw1BAQ7kSyWVsWl1v95M+XvsUo5Q4bttk/iqvcQ
WHj5umHqeAzcGyh/sUVI0uCYucab3tJOOdJtLbukwa9YipjDI0V7VXlIhl/40FsnPC4qKMaAwbt/
CPW7UEXNW/77YY5P2bdwKAIe7OyuMnHqWgfxuRxKAZoxieVogzEIc42exUCyqh+Ot/hza7L53RQQ
Ac4AtH9UEL9IEyV2ZEqm9WBGkwjKSGoClc4/PRezwLHtSh2YQYw5l8vgS9JbjlxAZWO0TC0zpVYn
yICSE7lmTCEw/u85hUQY1BJExWKUbZ2UDZMdWnCiSasY11WJ93Rs04LO2/f2ZiEfiWVRTmgTHG/L
E4puNDT/SND1yegMxrqBOHLFvjN45MMqZ2cpQChIMWrhHLayc2mcjwX2KVGl3g2ifh024OX6mzQB
WuqpsmzmA9QSUBCWEbyajKjop/jmfgaX7ZxsZjznHQ/UCE8EwUo28pdXa/7gzOpOkMqcN0jkpHk1
FoYL7YWBzZJ/RXabvwu7HnX8WSwJTWrL3+D8uebdF1hdqRbwdkIDjdgbLj5fnxILvZ1FVFyZT8Om
GJX9FGoHJBZX8RfAkXOa8mbhf6A/GLB9CIzNJ+SiBkbKG12yZrTqsZBZuSRg0OtiITzezEESPYFE
UAmrHdv5QcfU0ZkWpQlPkIiu0Za3qANfiV5eQU+34y/Xul1C4/K2ZbhgtapCkpnYvTTxeLVrtuS+
6el9POgBE6xDr+asgNSKyQpZa2Ki07rQlGSyrtDgGzt6jJTnY1ao5MUWwUpn+gv56/FPK/aJrjrs
ajAxds/uXOAQDGdbfFllsIEbPRV0O0yRgr4S9sbKmcTPWG4GBodPQYKPQfH9BElnu8w5MSagqz5d
vYh0QbIMiXz82hVfjWhO03XdpeB1h6cTwN4f1UDjweXgYnGYHPwkwxK6i8A9v4OzSmu1LVWbBZYD
WZ9xYoaYnYq+srdLasdLzzjXfjgcKV9q8rRERVZ4zQVpl/lWN2zlow16GhJhCbcyWUa9/JpqZH8p
3Ql0DeSMaczAnzW2vVdo1AtKe0Ngzs/5kkEb6SvxzgOLNWUl7SOHdx/HiadhQxaJZgbLFFfHsTqO
Qi88f9tLWQXBpBARQaO5vZq2l9xuDhZd1GG+2Tkx5aQANyVHr5cRbFSFtif+RbYvuRjPux91ZSjM
n3bA2SMDZfnUMlqcReFBDgIAjpXPN9c+QcC5wn6ya7/nQpIITeI/kUj230lbcqGhtzBZ6HJ7PCbV
KBbU6BAYrndrbh7sYdhQfpWz3tG+hdys0S6rxToJ8GfMK6n8R7X1+WsoCam0WE4PYLKP6kiDXKFF
INUDUuKAo9kTtYqEu0JNfn69NSVRlU/D/mhr6IpCUYOouwvkKxOkprK3soLlIgR78V3Ziw5+k/xN
ZzcLtGLAgeKv+ky8bIsmk2mQk2GvFq0Fprz2s0kbkDn6Ns5FKwz+7qFgz7bMn3vYfzYi+XZsXpgq
NJPk+P/DrqvymtsV45fYrP2+mGbSIc5yzN+gpLtK30QvJousf4nVG4Ppn0ZbK4GQslImApDqut7P
h3VY6KteB9gLYZSrcdKWqAyIL9ZWj9Vndifn77c4a0h4dLMTHnd+PcwJsCR9jzpqBN9eBHVKNC3w
0e01gcDJQN5H2/FEkvm7XGuVC4gW7z2QddJnDe1B0OWCx2hAG4xwEOCA7P/H6tG0vbXwTXBIPRwn
lz4Y1zs9sEz6WFqhdlhDU6fFJZNl8uBTfsagidaDt0tFhuql31xgnzovni6HtuNCC2fiBA6sGRFj
Px0A2a7T+Rfg6IWHugZLBS4QdeUiaebF2/kcAA483br46qk6YmEhqDUciljV2vm3+6HTQdhA88O8
IlCIG4iGUMdIMl3F78AA7hYyx2k8t4jLv0MLfNR1vZ34RvNLG4LivFH7mBaEMUBsNcCXCwer1+q6
Rasjns+llmb5yunA/KZ9QOlFfie+m3qjcZUe7E4FdSy78Cmw60A64SDcckzojQfWxvwY9UgJUlbc
PsftIGrHCURG46udPESyPOraQ1m3sMH/F3EQHdRHVj5Qnu9XxYDd5MfktwHbjPHO2MXmXKaB36SV
f/L0BHV/gvwwMlQNwdELh5UeFmcOMHglYLZssYGCCeEsmPRJ1l2JHFGoNSMiIcrLEeu3U3vD7MJ2
qZe9KfpV8yDsMU3qc8lo5A0nIx7gPyBVIFOwM1KaiKu0OOJGT4a0fgKd3yUXJhhBlxSVz00sK1m8
tZn1FtpPsaD7ay9owUApTjS9s606udW6FO2R9//iJBcg8KB8wVprr7wId225vVS3QASL25VO7LtW
aP9q/XkPQCmw2ozXTengG4HIDoah/m6Li9tLEfJiaqktAnJ1/nrdeyeDttRdJnnsXHBxky5osga2
2+43o0Tt2/NBuHspO9aaKBi7O6DwBRzbKeEgZTYgme+GYRFB5A2r4YMT9E0UGjtybu+CoVwDemmZ
YGcANLPHyTBYio8IpppN7h9kWrG3PGkAvrMsW5CmVZxfpJbcsrwUj0Go/DHpDV1kTiENGkeLTKTq
RwgcPMEXz9C7gsGgRnd2OjlZcpitHOWa2w7ITK5O1noWQzX/iQ+zPGb14gtk2MTRYBN90MnvDNBt
et5bAfJHhtcLsEcEUm3FUYdFn5gRKzfTBremG4vob/b7RaYQx+x+pEAGWYSUvetVG2ujotKpouK7
9teK682KRaQd/dbwF/QiyiotRmMdvIfiW75/nMc47b5GsS3C6cO6gDD5L8+wjJBpkljlhcuj35Us
7VRMpcNbr39Od4TxrVlQh0rWMVFV9iRZpHskfjEaS3ivHdlrHVEeZhZA0et+Wm+g/Zp1F7ZbM6W/
VX3vTfT2ytjIXLSuUd0plM9MuMlcHtNgB0zzOv8spsFATBmg6f1GqWRx0Bmo++oO6U8dnwnuWRbH
cHcMsOVbM433Ol3+G0uG+pxsuNgztUlhx5z4I3HndD4QifqryQHlwRrq/QTLgL7Y9P4xNQdjFG2K
rniPjXlGSLzjvmwlobIGZKAYJpw0GQb3If+J/G30m4frqSn1WjgvKd07h67LljAqjXNBpo9EjPcm
xwRe1cbPxhHZsTVxctDRyBTfytVsy3DnUrkU0iTn745omsTP++M0j2dKm6sQaiY8YRZoIR3FcmmP
ZtH4K5E0l484rNv5O7SF8MHCuAhXPN8t40tbwcyZttMjBM0aEQTSm48+roMB3GdilAb3FKNrUC/G
2BeZgxnG1UQwhXub32CUeltK5BK49jHgXrxE79hp3jj9+1N2LLEQ75CraDNtZyaROoph92MWhomC
Hj0PIuVMkjeVxUshdSaoEZZeXecMRD1zKXov8lUFyEgCplbRKkDReAfMpLVUBUkk5uvUPNLTXp1v
pyux52rxk114ZlB5lP6G5HSAcDYBbuSO9Tb7J/qdMPHpS0f3wzhl43J6MPS9QpC5413gAypXuiO/
uVUIECDnDvLxTCFosAPF7GxjL23KM1I7Fb71u3/RWb3WMi0GzI525sZ09L+flbdOgsqR6zb3A6EA
Ho4iRFv0/zYOebGbAD5i3rjkKKr/yA+m48lS2MymcLD4j1yPRa5QCuvMUWVIsE8zGBrKHC4sgUUT
uHXXH+7uM3HGhaPRdfkqgXtVgXoUA294OFBJ4BQ8Zg8CtsHk7+bBhSAXyWCGe+M6sQDRKr8Kl3MC
Sxpzkbq7cZGUFyuRyVzzktvz7L50gIW5JcQxPptm9lOlXDgvDHqvdcCMnrzopGjyK7Rdm2xs3hkQ
G1+g5w6yFW2lmpVdAgHIwvOg88sJnN2OvUPKR70Yd1Ikxm3VlivQlEklwim8R/LNPL81KvzYGhlv
gVmQ0ikfvSIu9qvMxHmR+ks4yDym9Pove9GzaGvk+HqNDGqWuxBQskodZMg0sQJEdCd0h+H9iPnw
HjYt+OOkN2G+KkQbUZLEip85Kkz6/rLBUU1kok/Ds94t7kVRNHlVF/tBW8aQfSKbzZhWinN55876
9tERj72dqkAFxDgRwyt25sDo5tQ5llWixn+P7AxJKPmmizodf8CPSHM8Id+8MvwxcUITFpLT/YqD
zLTxMRlT8334G1w3oidELE382vsw6LViACAbGbm7rSRmgRHn8+XWjXssRpNHrjj4XMGDr3gypzmC
2v9+fSLAdhCKfCCh4AcRq3H7DJDIzKcjmzspdiEYRUpV7+LOFnEKdSF9NsFpt6WTnSAh5nziZgPV
lgdIQEW5Lrsk44EAAygGUOncVmDiYIDYrNU2+dxfheGwYk+wi6Hey5tAw98tkbkOBLptdpeDEu+T
/CgDxLX1EjxiJ/fedrF2c9oQSUTDXfz0Sbrjq28l/jeHdZikPIwJA+MntGVZ43p+nPDNbt5GM2z7
DaI2mI12TFIWytUh6zdUtTE4j8qOOi1M9I8N3gBNxpglrDOtamsiWbhE+bSgz0MuXh3NAopejvxk
I3b+165o67Wy3YiZhlYM0DoP1yoFg55/2Lyd+vMtaEgkcvAuBe4Z3XQAU2hBDia/IjKC48c/dhyn
7KJPCT2IQ5IWxAXdmbyOfAh/y/iDEVaDsNccUmmlxdgMLBU+i/Nnh2rJp8S8XBj8CBdd1hSoU7MD
wrBgjbD0HsG9ucziTsXvL2q1bsfI/WTzv0y4+49guW1UotRxHv4pxetSZet/3aLy+mo40miHy2kG
XZ+Ij+xvb2FSfKtg1qB8WCKOY1Wu76+M2FJ/XAmegMJM7GGV6cg9FLhm09zobYkxUaRABHJSIswK
B5mZXUfTUxFdSy/Ysx7kMhe7SYMN05NoOLnfqOKJQgu+ShBEq74deEzTI2ETl15DvwsvqziYl/rk
4sG1ZUaiWgCgLptIkCaaIQVm+BAH0B1nUCT2KPYAcQV730k2Dl+8y+lM1YuL+20+nteO5/wFzNmz
A9W6op4dX4L33lVO+XOGiqgvOMvJWpMwBXtdXMxjshaEn+iPUy5e+U5HlqSOfDqpLuIlQNwWw+tN
dNAb1jtXZii0v+pKz4m2L06xIgzNp6h2h+43yjmzXHYt8bP1ab8vafHkFX7fRYyPJwbz5sqwi5K3
G7rDq8/VSO9eueEeF8Y+iCU2O3FLALsugUGVE8paukvaK9JVaPXDmbjkAHKSHDbM9ne2Ej1mtb0v
Oxf1g9KZ1oPwitTEnygqd1gw/a8mhacOtYbtS1tqOtKw7CLM29FTF4jTGJ1zGH5NolKQ42ZryV+d
rZHN4Ca5laHiRdO2c+nsT3KT9OhR3LZfRHtdGQwF6GvwmUbg/A4J7hWuRknrC3dwmKYBgo217EEr
TKcmyPLihUyjj6WLHptOCj71yDdipTNg/LzGHTyHcAlnJSf746K//juSKIoaTX3YR/uk4U+SYINi
6wD/9qSWDDgY6oO/aGEG+zAW+1ivnrXjS7r4ibppx6n0ipww6YEZ1BE3A7lReZRy1UYRy2UseKYv
zZVCepRA89FzMA8Wys/RMMSqbhrJMs8/P2z+jcIU5rG9BRskvzCp2H83fj7fUBVxe1oXhhTpKvhX
rdyHLspIVifaQ0x0N+GsD51kJat7Ml/3GMXTyFmjyenowMDvUHVbMu3V7RAzfU3G9v8umlwLqmno
btWFGTBhVL+PnWf6ru8WeB1gVzCnsrvuXnzmr33fpLP7pl9Ahog8KJpvnTi846HK5XNb43VSHpjF
gVVccCt6TWrq1pMbITUirN2g8izFUEVW4RtVg6Kw/H22xBrcaekfE4Op2pUtkWNi/kWBHLqGxlQ7
wSiwaf+mi1VLWbHov/HAlgHwVH3M/4ldcT5y9eOSqz8e1LrhfJmwi18Lq744bTnin3JPoy7MamOa
P9mD8N8uAk57/VZAY7Gy9KsSxLDntOh7OLUpJ70d+W0x3MX4fjAr0D7Hawvb86tYvlwLnfLrUTVv
5QhC1M5Rqms9gf1EllxqX9VQ1CuOpjikMfap44VZlujPwFbd5KQD+DviHrpNVzQUNMpmPMwCHuon
7/RkzjdbAzSo3zZYr6emDvSldaiM1htGcM1WA81O999OgigTwfRoMTHuvhPnYWCp1VawUTZYQlVk
i8xw7P0YZwajqE4X83RpOwKghc9k/F6C1XNhLRdfnOWNiGCUyZb+ZQxlfL40c1t4frxbnxBHU5SI
ztGqX6xEKuodlB1oSvQEFem6Q5FLBN+b3nEsqj5lX9IBAcBwkLGF99Dd9JAohWkRlZaNeK8+B30y
DuG1ZJBgLAZe825YR6Hx/bE5TV0H7hwEcmCLwvoWwmpST0nmsjjzRyiujyt/VqYw6E6U0GM981Va
R/dhgjfYoDgO9nIgrwQEGtyC1cfcWix6XEa4jdDQMBBNAubNBYKYJbJFETV4Vw2CsfFJ0RSJOUMv
/7WbxJTvbDXauFWuko7/UWWmZKMVyrxnbpMrMsy90CzCjpr1xngMKg7gdkSpq4dREcOrO7TZafxD
8elL+28Lyx1Pjvqdt4sid65SpTHSxtkq95kx1LwTX3BQjdyGwPJlRJX9egwDzpO0XaAFr9R25MqG
5Gs5eJS6w+qqwq8QpT7AIfwgN1UiUgMR1cp8xOCT+ldLwMfyN/jSEQCgA5coj043HEFzjgLohUyJ
li94LXgB8L/yN7NNuyRtn7oC5hJ9dwDnyd4AU5HSDKmrwJzkMjrtb7TCiqnXMMRHsLDemzgpOWjz
gneugGsTlOJIrbWpZirlr0FgaOgI18mVstrT2Q9EjFz9vLAeVDzv8qugJahylqBT/PN7Z8pZr/0/
/nksDN0K16/3vTOQ2gGh1IqxdUlvlaZAfOU/dUdtIOqcBs0X/Wy/tme73u9jwdjrA4os6e1RGcYH
qQtcgHiifnLi4tq8yfoGRaQ2KDHBCEEgfiBl/VF49TQXSTVgH7n64JjRHuDGU6uBDZPBEYHAuStA
HMDUaV+9nahzhHufWLzkNLG2HszDEZox2HYnoFW0ROQvfl+mPhlqYu0K4cKdY0h6pJiMX9vfeaoo
g/i0HDNOD7HAS4qkJkfHcaHku5RfEH1lnojWfMZjZYnSRvCyuF4WzcSxb9t7cOttjzzpIlCgGlmi
cTzTRPj87p57bM1usgolW53pMpehSRmytq0npa9cxjZO5Ge59uildOrKVfN5MwfzESJa1v6LZk3M
wX5s5XMxWetS3JeMJpu2dyxDCOqSxPPHJ3COln/hR8d72lz8m6mPcm4nOvTqC7HNShQXsNEDfNwv
iu+Yn4h47UJGAhtZRmluC3sbEoB8HyttrWLiZcesQK2JvXOrPBylo+IMI5gKo2hHWQAGVHwJscgq
+loIVv3rICnHdYQrHNae6Xa5J41ELUBEPgXh7B50THBEbALRK8ibQWB3GuoHfcMcuNCeCF8KQtCj
ll7iLwVfgJbc7zMQ8+2Rq35XlQNrwLNI2KzYGlqebotvoaZPvq/C1vmtgA177S01z5z0gXTTE68T
Dop5sg8+qA2R6EbT79xyDf0uPwJ8dhNB01Y6ygPvCoHx14NOQHNOipNgga+TN/TbIubHNrJMjvZu
1KsjkIrVCTWaCSuGU2kTiB/7cVNWvvx87J3JigBfrFGbaye31zvvqEw7ULHcl4MeF1IN5ssAufk7
eNPy5pYmxwjOUT3vWN72SFd4qO2KCKUKYL67ytnA1cXaE6Jv1+TmaGHfBGkJx5n7I/1TkWBAzCFo
NIIebLQ3p8zT2PffZz74pWbF8peNfJrIZbrDr4qFIUKIwYFRQOAJNZb2ZCh2bPtcn+2Eo5yjWCOJ
MMTDiAFWvjXzu3yC39TCz3m4uwf3fH+6i69MvMniWHZduS1E/IbZELFB9JZXx1e3McQQ1JgadMa6
HdvsEaElkUWT1c8Kx37aaJN0rFURIPj0e8WrBc8unOVbyXGTJC/9LuF1eRt/sPv4sX8uolO8Fqn2
iJYRYJ25hMw63++Eqd5qpuMG5k+9ICNtG2sWcuKSN3P5Q6PigM4yyQmeUk4zUVg1LFfc+bFfvUml
iPWZOrPVrHZ4V3PG+pXJkxi04yUNHYiL5ctn+cuJwMsxBjBiczHN5IbNOfy6Kv5ZUO1N5Fpk6W3z
D6CuIwTzGM0D3GxU+Eg6n4iyijyrU/9q9IxFdn68M/yTboJWJQVFxj1FSNDPVxW8Kk02h+xP3H16
Ce3055m3nSTEGtXLBB3UnmBWK90pcyv1NSdI3rhyXOm1gmvpcR7uTBxKKOkiEvtkdHy0sxPpkmIm
ubQncDIwDY7051iHAywEDQAWhkAmNGQl5qpu5x1vKeoreaym/mziBIb27NQ7pguuLobBJLw+rS+Q
+q7E39JIlsTEQSi54+YeZpWsuU9ezts9opnW0tW6w08jz4H8ntA/Z7iAZFnzbvMVeaGS+wfTwGI1
LCmtN0J1dayQXYJKfVMFBGLnA96qI9v+pcZxVPgObIhFz82FKFA5K2G8bE0K7gnQhhkEWnGoW+zk
VHPT0PXQStJS/g/B27xArMBPgPW0uqOOFVh0GGldpfb53T6FwjZSbA1nYKUx0Rbkltyb6vvUHqv/
I0qLEpwv7Su5NOlGMGBTYgFeDq284EzpgqQHFbkSg1xn2eDdqaRNCLf/kvAjOoNHhrZafNBEQgEa
zgeG8eDVCvChmqvUw48vKvnHI0zYsiH8Yl7SFXESn1gyKNXmozTZw0eLuCHk/V01I1K8QAlG8JIH
ADlGpQdztLv1YJMuQnmSsW/MptrkLy1nvv3vGhlj6DyNz0ecZDx2sMt1DvfJC1wBDfCR/LRvBbHT
95gN/WMBINf4S5z2Rzbm4cvORshTcDI8IbhjTytMpjdaPxTy0boZJOiK7ByXZ3+voAZW9RTBm3SC
omAja9ZmUMX47fbcloxSt+dINb9zbpss8MqjZ9dJFKnieZraEGckizyxEUDdsbmR+G4Kvo7CjPrL
GTPRZaqS5pD5SqgcQ3cDetnpLydyxiVPehXi3c8LdSxWlfPsIQrsMvmbjr0+pgu1BFcKO/MnTas4
cTuWvRu0dSSE/w/Vsc7xw8rJGIdUwz4kNZUI95QB8Tlr/pcWUlH7FGzzAJ0be8effAYYKdr0UbYK
AXX3nk+uo0KC/Z3Nh2Ty5xzqjxtvzHnF5jyYNVKQurgpR7oGxqyU2CfpbNUiDk8GcPMnx8mUz0sX
+OVjtLk411lTi2ydIab+kcoA0NFHOXfKlnD8+zwjAL8gKDbLoJBnxfXq5qf0azdeGG+eQjSVItvM
0hNpHLRBabOjHI0/uJjOteEQ7/MJgGCB1EuD3tlS+0EiqmVYi8TqPYjxbEuI8P5WrdlsXKDXrt2K
odL/R+7gPoJbfQu9lPI3IstA2PEpI2VHx92lBSt4bGQOOyK65fjQzMXLjIXf9gAVYD+Ir1+yWf4S
Lx5fzzIVuvIxO9fK6CGQCCzTbhoMYsFlPO1zb2ijlbirjb//wEDwpGGjJwkQHNQEeABAd7SlwzG3
6IwBxGSE2fGOZXZYEIIuK74t3EW5xWKJ3asA+vdS+asjZ9YxkZJjsfbjiCKeiYosjqzTUucQnO1A
PdGiLl2KS9vUJju3r6QQkpHgYjC618EDV2exG5wxai1sBepM86/5Efi5GLYU+do6tueCVmets+Zr
wZUEkUxbBnmpA8go2SDyzBkaKgUQzId+wU9Cb/G1ZpVlmcCvr670Dev5bhUKPNpaVOeap9+vqUmE
r/lU2LmmuudbWe+cE6oEM2vgUIF8j9dR3w9bkpJEJbpjg201Z/A7QHgUD1AEE5E8ne8XrGHo6BTc
OVZ+dANfDOr7Ct7+VRUx6JSP7qRDCa+S2jjrZLpB/mVPiJJl9GFqYHcb2Aab2Z3aqC9dxZ4ZOYgD
WYVdOlFLq+PE2h4b4c3bfDxgenw96XmYLjTCPFPkUBVs3p1qPG5M0UtcsP5/UIQ3JGmkGqKqYKo+
RABCeEAGbGfUhsiop+ywzI4hmGdWoD8Cl5CG14F3HgQHvxG9KQn+VqoiLIXYwUH9J9Z32mfxYY/u
euPuUl9MNEcBON1L7G3+eXOJYtsC9Ra6oBu32lfXnns/25PEXQ8Dyv18XiLeimni28ITM9HrmA8X
TJInjHhBEmtf1wlOxEgRQLEe/K5E0ouDOJDXDavrjb2m9lA/0QQLg9nkgg89pk9q1qKKJtlJx4s1
1gaJN6/NLXXUy4OmZqVM/azYfp4tQFQx79l+3bTqrfSp4UwJbNHo0gEbAFnDNUMsiseNGjJlzSTm
UKLcfQRKyU8ut64sq9423bGbZSzXbbhyNg2SwK2IznbynU3AwMbyh0k/AMxf/r+otc6MOjSAOnAy
acMOjl1NZDHftaI75lcMWw37nH/MsGqm3vpAwF8ZFKbYQYb4Cx8wmU7B+EPs0EVyFHEyug7R0rEa
zFptNxo4cmlNNduSv3XMs7z2fxGSKZ0CCberuSSHRm+lta5wXm0eY3x/L+3hhjoznm8SSZnWiT5r
OjqQwYwo7FynQmxwvX2eYA/Am3nUjnjEJr1qgG0MBCMZd7dw1CDR65o7HXYdto8X/L5l4wNGJ5Zy
Gb+zHn2j6lku2dxWmLSH12vw7/XZ/j1KasjBKuzmJ1A0rMyzZ+P0O8EdznhjVc3Gal16+E8Ur3Xn
ma0irutlVsriQkqUYwQNlRmljWs2NEjhZPbQcMdbwm/oxb3Jcs/FRMNOKZ11tfOerQGWPQ4WLQbC
DJVArvw+J5XfIysl9qYN2aND026zRtjR4fJ7W/ELfnzRoXzXQyEvSDxQLmCcqF7i6wOzDB/c2l1u
hGD9bgEo7+sm2XcKkm1mreqYRWL2yG3+BEMNkkWbZR7+DIKmdnP045fiRxG7u2V3OLPkM8/5ULd3
3iOxvr5xFiFHSx+ZwB9UAZKfNt34vG7GrUy/ZFAZkn9/DZuZ/GoDiljxJBLKGY739fITOt+UW7XL
TwZFW2jSJ+rvURA/CJk1nQ5tnHqebW2VwIRC5DAuK6d66aEFIhXpHEsxRFSsN1bkQ7S4FWcIT2Av
JT1MdYRk8yPp7XVD+h4XAAetTzu2BX8RI6H0sn4k9qiDUfjfBMHEQ09WkofM8k4HN72P8VvLnc1z
ANvf5Pt73nmSpjIFda9378cxPyrNsIxg9BmpS9yrYnLYd/dmqm0qqa7+6Bq9gWJzbR1FIJGDEpDl
+WZXDcKWPGHSV5fBXXQL8KgFfT1Gij4wMaE0NBRE8HKfuOXfqdOjByBH++FZ69lyJVEzf4sHwk6s
vOt3PQzYmwPgiF3s2P1CABwq+oMkpjLcsw4XAkEmMUrx13oThkHC3abF/ebywt0Nnhonzirih3PR
mYu5bupZ9UpJcmWsa/MfXpqmNCZ7FmFnMHnEQ28YGBh7WkB3c7KMDxY8XsBCANZUEF2iH1upTXBx
N/n0Nz43IegWxugGh7U3knT0MIhk197MszVHJAi/CohRDsEplFncWHd4u8SQL5Pkef89UIS4U/F7
UwACZNywOwnZwMj091+KDXQ+ABIMqprOe2GRCNExJgMbOiu2qe4q01t2CJaUxy/Y1EELYGJqShDX
0ZltJDauPc2kWxSuHgIjk0sk77khUt4+2JAFa7wlfWARCQ9gUx659ZpMHVPNL2TkfRVWOAqVLcjU
DNJAviq5eclY7EVOV9sdMLMx01XYARh0aElWrzVxVGGArp6E/pdoIxB6ZWqc31iTD+DUhA4Mgi79
7k+KeEmWLnSKZ0pByN6o0si1kUeXx6VoVluzo1FiGbafAspnm3o8TGpsctalterosLW824U0nERb
pyuMCTHAAvobdjtKHQaMnQMWd8y8n0+BUt8c53J4aJJurTO9ls6ziCXdrpgpO2bmwegESBnVtTun
6H5ZgXQm6QgYNGBYAcqi5CgXi87kdDzwHyHtVAGbTb6+7dLdxpFtfKUqqdHpavtj87/HR4tIhYzB
1BREZZKXkiWVAPOTnB8Sp5rcuYZpMQVJCYmaef5o1qKGCfiuHn0ShuZsSOlzij9bFGjIUzpz4eLc
v0Rk5tgnQuf1BMwJIi3wuPxa1CYVvFm7Fp9UbBI5gSYNFzi3f1GkQUoN5dF5j6yR9QCM/VVnodjm
s9HesFvCnKxvRt3f+lc2F9Er4rMI8aa2mz+VYbymjkrQJAURpA5gyB711k9HwLDXgwvk9LyGulLt
2vFiUh/V8y7ftq0r3g+JP7Ir1rCWcvvRiX0kzHc7guJiQ8CeAjYrarLQmX2PYe49p9Hx1TrsWPdW
7pA/ycrwbzAxNGzeVJZ0Vi5KAOt2vckXyclV4xWrEWmihav8cGmby99q5vsaNoLzCQldUNVqmJVz
Z2bdH3UwcEf4vx0ALctfz/ypJ4pW7Oic426aN5GY5Fvs2Anc6hz8ljifki+cy4PL7hsMDkXquUun
kao+wj0wSeN8LpYYGi8FB48BdjDpyb8XY+bIJGd/AcACtccMfWUNNLT0kP9o2F+zh56F7dv0Jpmv
A6RAMOIXYQm2otEGtiqIRis+ldt713EhIiMj52np+7vWywYsU86CCeztk/2IAhavuygDs2RFtshh
mbz2ZSHed7ZYWZrVGl1TZ6E2wEBJjaERaJ92YWT0jJzjhGgz/frWQGHqkGjojjnCoi2glUAfvbuU
f/fNt4A+ca698+UElwFrKWQC3GvKHFnTeaiC2wHUbWF5ea5JwDD4nOKsGuOXXZETLYN2vLp1ULjs
16LWThH4I+rukmpbau88U2nLcz9gExpnlDlRwdo6tF0Sm/w4+Bc/VREpprRolZ//M1MwansQ5dWT
Pqp2Jnn9ZSjTztCXs9Bum4XYO/pxbKJP9xEROGK/qVd92aKrqSJauwf6G1tXnbmK4teJDOo0AQo4
22x1NJ1+KszUZhylPtP+ifVh2l4zjTTdbXaopDq6y6KjKLE2F20rXjEOFwmgzOsEH9oDmNZFnGVw
NTPnnDZGmuwUxdBu1j9uuxZe5M5Ewz980CpOfvKKyNYC3KwfSbacW4lYgUHPjdt/cfPYI6y5CbWd
bYBIeOPPLWAWWkT2yBBSMH7+iKtf1gWD/d+Q4YwurrjOGvI+LvRcu1xoWKqM/dZqTTSCQqfYs/2Y
BmRmmVlDUNM0Sm+uFOObHX/wMio6XcPH2V4UDtXTgfr2DW816hjd5wQIrFfxTtbPpuYcnygS7852
3OYPJ8UuFvC4CFLvBi5sPraTAAH/uxOsfhFvEOlriDsSA3d+VMzu4E1c0K7v2Sm51S4GZP0q7UfS
pDpuckw2dphnPFlGkaAduMpV9QqOvSs/iJnXNxZcrcD1seGJAXSgtmk4wfonVWzFr3G1EqU6ZT5r
slu/diHQydSMp83h7hxjNc5Sn9USnFn/IUm+Gd26ooOiFNWp+7FiPf/VZL5UR1Awn9k2rDydWi7R
vpZ7dLtcd7xTMG/dWlFwP4B/vLrNq1Xl0c17oIybyhK2vNiTvtN4n3EMcpXosYIUK1M7I5uY8600
vjJNLLXc8LYSGCbar6WrapaEm7BmJPd/9y7ttLGLP+3T8rqH1XGlLR8Myv+FZpeJ4RUm/HOeeS1C
0yyUQgx7GGDfn6u3FGyqZrObnIwMQR9+zdyhBJZGW6il79g6W+A7GwbgtYPSvy/tH+Jqp7qGkOWo
WZqDQAgJh5KuYPBL3xlKQJzpb8BrVTRVXarQT0qqe6XKblcCckKQknVIovyeurstbJX11GkoIhdf
i+tBgJt2CcW60WtVe65xeYUnA9akC44Vf66FYG2GW+a0/DoqaAiqpA8b9yvuS4rEcWj4LoikqygA
fbFNkIFO3HM/scIZ5WsoXsbilD88OmGFjJ8gvnvzNpKbvh6zNFYiVrQqLmr8/p3XRzUO47zIrWIx
0B7tx2TgO28J07xmkbqkAUuVjqtkkjJV66il9Bsgnj/KECTOA2Vex7IjFEvH7PuIQ/r7b1ErHdzl
lx/49mRrs68UD/+9Iy05Z/8oTfzOY7z80v6o7XbiYZE6WmD9/1/zOiPO+yWVeeDRtk67bQ/zk2AX
r6JBqdpdbK5WoousGHDlWGrdZIn8UFMWwl+vjC+V/+CJGnrAcEloehtV4nd/DqDl9LGxduMUDJXr
0vxTo2xRRnJ255QUymQ3y8y/LBvuaStmlpdbKAlUFEFvsg83jBMH9r5OTCxKs9TEj62n+YZECDcl
LrLHO49DksppwTsbzrcBhZ8+kC5/n9vqB5WPirxkm4Ji8KCMWmfk4kOY1wGJ5UrCrr9+r3QbLy9J
Y7uRJJceR2pWd7FSXRvBmeRpLUCccD0T/HSzt3SyRYASfnNz+TIcTMi/ZXFFNTSEdbCGaJkwyv/P
EgTmLxtqZjrCsfmoFpLSZ3i/UcRVg69/+YAVR5C29MTcdt8aP5J4UwmqId3V9p+zhtXEz1o3mdqc
E7/iZQXaiJi/wybRE7aEDpvhvm/CKvtvIqXY0ka3UpX+tnLe3K6INv8Xlsq4AbPSJFlnN+hJkjRP
dQpdLD9Be+OJCi5u0XWGzOOZNAR41YuZEXynZJ2788sOax4H9bEDmM9oNsXHOUW6/kBZQGRk5h/L
VSf+4LrFfIM0e3vkqBrBi18cu1zSkNtpTfPNjjbcFRj6QrYCKaLLvc12hSHQXFEaKsieDwGb9gZR
H43XS6mSLjo85lB3qAZtewPj6EzLy1l+p+E23SDm/UKX5hGY7dleZ4GadBMXQtuph30AAnNPSnla
ZR4O55b/vzmiuYoY0qJu+WCvYcPBnrdU7oEhKcoxrkzf2caPB3PLGeWFTK8kXo/5mzp4EC8reRde
Fr60/GMTsjw/TnlbhzSUoKOCCrJU9F1LSWbx0lnbqqca4w418OXskQlwLUysQzpcnUWrxQXNvKhH
yfgw8AbYa1wRyZfuYb3+vuSgk/snKaeOE/oWfSj5uhw8zRlcxh9NwYujeySEUJ/iQyzY7TlVsfiy
C9YkQE+X2T34VMRSl5nwrTgPprkoXimuGVI7CbkGsioyDiXr+x+49FM3nssABCtQ4F80i1xFnOXa
AQ6il6Y5dBS5J6mbJG4TXdEwNbXyk6iKZqxa/0msaZOD3nsPQkNyXpHYJzhrQ2CFEm/u54DnQizC
nNj0HLKgSI4ETGV3XA9wf2hkZcYmETk3LQC/+YJJP/n6nOvqJwQlSRO3703SUqP2V8O561kMFmz9
/UIKk7nbcufufRtfAe/6usJRCVP2axpr8fxoiX+ECwCMnI+2Jx4olPu9O8ZNRjrtZDYhZzvCFARW
EHd0m9W6WxUG8Gwn3UtSNfqsHsFOI5FQuKcSM2e3RHslqKeWosig+L0uwoE6rx0AYpI44Y+XkACD
KNtkhuHZgsAYJM5mFwWbqrqBQMhql8a8z3LckoWBaZfuCd41TuCKFlgL4mt2BN7xZ63TiOudITui
oKA/W6Cx9rG2vIPQ9bvcNgiiCMtO/XAFiGj6bu6RvnDjQGV3rx46mRt3b85LEx3ezht0LGCMaDeg
hwFjO84fVUJad4owdkvpAePiIMG8xmDzWAgX2itIXwl/yb+MgZ45IeIWnVljD4OpcD41TCacilE6
4WxuWYj5yxiizEy1d4rFOIjdSm1KeD1shXi+TGxUj0LU8laq+/Ulzyjsqdbg2/yNFEh9mw0kPitr
VXgmAblPN0NtXdt50yAgkL87CNzGdafejXTds9nnmzAGxjDgSfnPZlhiBZUxXYpGwQBpJIJ5lbqh
7XIkfouAqdE6f72uJadzSx97dml/b/gt2KGpFImTnnuY8A3pS8SrvKe3S54HW+zVJnhZqnDOZ+kI
306kxcs08ZnapBx4sGSYsOfH+V1sphBQOhjCZjiBEG7gi1jRCRQ9d6Rr9ddlsSGT7Iodt+h0nlvZ
pXY/ysQV2n3TwQzmR6Sl1JMlZ+sH3WcdYzQKsGC8+CjDUM0CMm0YPtUgER7JGgiDeo/oclXWPKci
BbZWppZA5Ymzuwd6ojIk4a92MNyncA7X6VLmy2Lpq5MoZm0dapQwxpOhjAWrE0+ccEn2ARJ21n/k
uadqQQHbNxVaH066pfnOD3MBk+uZLMZ9feTO3GJVRISIsH7m7QEP+rsr+Skf7IVw8rZAZngJb7Gk
m2UJoPxLa0UqerWhNdoMuy8wbzZeprIBb0njB+Px9IgIOAdnl+nrofQtEgUtMM3CfAExl7J/4zls
7kSwzCNEdJ74FajHyiboHGu9IPsFP/xl3SHwOIaMQb+YacmF+1HGOwMJjjQdD0jk05uTEu7qO7Aq
xlRV80sSJVm558sW+6MKuTh25krDIUzE+yFu/Xd36BA02MToN6340N0EyESyPnAyyRboSiW5opPk
FzVoFfJsfRfCr25TkJ7v2jwqt6CD0gYv2YeNGBzTrLL9EK9tB1lAu6eQ4jTSf1ozVfyQEu2VVPUf
fCT+0WJvNwE60dw+kmSBTh+PY5Iow+gp6XcwXzGQVb/K7HjWPC2+RIWgsyox6GR8N/8z638rxXTZ
8CK7+r6vYv89QLESJnSAmrNiNu69w8tPrGbzWxh2OfV1C9UOIsrGdIFFB4uF8B5eDpSFXxGJtYpK
2ANIXbBLhd55tWl8e88iUppEpf0tLJeNcJ2gdAI4lsOkFsBIoEO4nA/nWoUyouk6FSBGY+D09FqX
jLj2d3MWLG7DOVSfUsFUQDVfAdqlXcWXjKh3KjI9MuDK66TOmF8snwGOdZc951s07ethIfLXezI8
Jmu/cpphUgSGeMFGY/uGgvqLVtMBKywdcmOCwbvDcod1vtZPS90p2C4huO9E+za9fP4XAna3j1R/
U7/z1efQ0RTpq1N7cXu+GBkPJAYyKEN87PYqoTmWtNN17eqPH+5aXgyo0w4FeTM7bWkpIr090CX7
n0qZLV4C1ozAU/OMr82MDTRmU+bxmmXNvZlnwzkg+Xek8/T7tev/96UOKqrV/pMjhdlV2DSERczx
c1J4AWka+PwkswYOkTMB83BtTmrwc7RLRXpz53VkF/xNXSgnYInmWuvrpmkKWS2kOjSeHuR0JZ5l
I/bLQ0AlMbz2SfZ1/kHyGFybIipJQggfWi7aGrqgBKc+IGmOfGkMze5sjYWnLEsPURYAP1GnOMHd
n6c+MKXdpzsVni/ExWVlH+ObyHURqWn1SLgNkY54WAnWgs/jGxcElvmsO8OVLODIZtCW9jdl+QAE
nWah4hrpMa/Et1aCT3dOfFLNSZE70ezOzGueLKwz2yu+iOrWuw3/LHaUR0U1xRuxhCiMevNiQtOU
jBvmk0mF2Umy+2GZ9DayoeBbfN3ZjXOtvpw+i8IvIsqzKmjLEyffcVB0gWVPoE1Ablk8+Eve3Hl9
3zGXGwNUoMLZ4REx/qdF1VGqrs4WEWe3yBs/Ik2fl8ULIQVh+fB07pcoUOuhDgp2V9b8BgsH/nCU
CLdOalQfB5NKbhRxbQ/SVlFUERZ8XESPtR5ZSH3VEo6tbhMUrmJIxreueujkqK4HYtnc/pW7X6Vm
p70OVhIPLpQJtVTTa7W/BhCl4a5d29Jz6lQyUv6HlEjmq4Gk+iisLwV/5q1jWBnzQzYBeFOVRQ/6
6lbms02cWnxQS6/6dZtLnDbDlrhZDcF0JWdltbFxaMsHluw7a8LbTlMMrlXhxvlckM+BHG62Lz8J
f1BIlTTZmg6NAoa/UsemejjJB3MuiZWAQ/aSc3yulnqejwk/bWa60PA3Re4kEkbunQ9MrUNh4FFu
KarhHmzwPOtGsjUIDKHNAAbzGpuGNGXzhRBy1jSb3zNUzm1H2Ogwkh1Dbp95ua9RH40Se/GKx9lk
hK1TSbhp2X+uzH95RijT3bKrsd+RsVGemJQog22G9S06f9K5BQH0mb+1/qzgkNigO9111FzgJ+uM
u8Wowe64qu1LkU/7YRBPwamA3d2KLkbrq0O0unipyjhyk/BR7nCtfFV7EuTpBqgvgdlaSb+CAyGy
2HFQTTy/Z1NUgS8MIm6lITomkCnIyJX6K3EYyleXopRMfKWzA1IPGn/hyzZGu4Gh5KX3MJiI7Y42
sbVy7iKjaWZ2c4jfx9t6djjjZzlwvX8NIOQdazYv29Y35JCLnREpRpQJTfz+/NmcCzSCn4z53HuA
frqMSqUYtMsik+nQjidN8qSJo3UqPgcY9nrJbesG+/p4QNHLTkyKT8JHJE9VbK9OnxRwxMPXobA7
Rq2tmjHIW7uh5XT+vknAbPxiECsnArLjJ/e2PRKQqPshdnwjZprjSjmNLvBHR1qZuoniJOwWs24D
txhHCKaLYWC4Mvdb0mYEEP3exGlS/nikwaklJb3bpwcoDK1GKu+iGWnz0yYx5PjjXBX2N90ErxlW
N7vkIc4X3gEkVHLpm4QrNW/IgTE/nSrgdMA8C88h+RPEkvNtx0B6TKOyBxykmDdb2y9jWjJ46L7C
Oufj7PQRsno1tr5WqasSOPeYMZ1VJzR8kiJmTYfAgNeq4pgvZSa8JS2ef80Nzd7+EtDBh70monKb
BC6cdqccffLXed9oBiICSIjf1fWr8Fkyflry3Mdao7qb6svN3TZtCxyODQE3h+EGsw7TFa4r6Sni
RxLX/z61ikplG7JOtj90uzWDUriZq+1TySNACtEGSyXvwoU32nu/e6uzS2LvY6ohVQjMi2uzbkHM
Fu0YEPSiodMDlmRmImwpxYUkIDLsp7zFNrETYa/3qBM4c1Kb3RYKcPTv5iyUN1l0Biv7i/zr9bBT
1Xu1SfA1QZyPbWs5Wv/5GHE0Dh779T46tmVCyj3TSNAcrtEPzutd0xJTNrsuAhsfWqmg5U6y68hU
0gATI/EoBOpjp0NcUTYdtu8QTLeiTb50eTtmHr7iYl3OsHWUlnBCMO/puugseVE+fhQxWuiEKnQh
OTUNe+4NKnSV+4OkOJ9iB+QjXSDLTgj6CpRmZT7BkXzhQGJQCYqvarv7v7Vq7uvvDI8An5SRrLya
sfZqqMsgBY2LOTDFP00oy+qJxZ0AHMzkQWYpQHxKymZ5fa7GBT48SadjNv5QQegP0dyX0bOx85OT
tkXSsZQn+KFIdM5yEVo4Ji2T/h6DhD1Z8bl9uf0G4XEsRcFaVERLwfFJCi9wI4Q3d680KUIhh6aZ
MaNJFbhwotJgPAQiBMWkY4KwWZxnZ2nFL2rqpEVD65bN3zd3sPS1iQQvbmLV/Au9c0DEMEgrCLwN
TuJkds315nS2+WaCSTxV+UY8IV8dddAhgQVeh3PJLGv6b9uw8o054Rpx/WB8+n10PInLNOhwEsXT
xE/mutWtdAAbL98mi9SplavUIdlBNlqEuNdxvqgmmeVFqHe2KXscRP09M3hyjNgo/axQMowDAjRX
SdEHXUcNo91DM5VVb2QAdrxJBn2cpdXWOIyXdZT+G21HypBL3HH+bF/EKGle05nQxENaoFQPvteK
D3ObhqkU0Hj08WjqnGAtXtAkX3D0RPoD35Ei+GBHbna0fIH5utm/2BRPKgGiqp1vsoBKQqclEHoM
rQ6cM+42kg6qrgCqRKX1i5DMKIC7+MEYJSjINiJIIPzozDbo982EwLzxTNnfQw6hBydVZ5n/l/+E
2SWGAKfjGzhD53WfzbcTx7FUcwVwH5huWb+GFAVnu6qfy51nvMOewlXwEtZH3ZPZ8Ci3rx4cTo0H
dqfFxEGhyUbMJJo2RDAjdnSf1pLHFyCQwQnyhW4/W9IQwcap3zWak9hoQHidE5A6oWKF4YiUezMV
F8uOui2slWlYv5B5UAEW7Olj/riG6K1rJesdT1vTK1IdTDfAuosXUcWZ3Kjmo5KbHuoYxvbOnOQG
9pAnub6bu3yDBvNSMXoIW6UDwozKRlWC20Z+1rJvFGC7Y5c8i7Sop8gNZSNdQpzIXu+Kcf4RiSxD
foDRJZDNZq/MfLSrENQbyF0GGhKPtjt0VIXgR5GEQ7c8LPkzwuaHx7NQ0brEE9iP6owuDO5uQ5wu
cUEjS+uo+bPeUtpHSx8+QQhR5P/O+7/zYczr/Zanf0udHv/RNx6TGiCEkPuZGQ703NNe0ILwOTPK
EF+pCVg9YVBl16OMQxznV2ZvCtsLBNjj8Mhd+zJxUKl0Ml2LNyK4EYcRYEg/mpTApNHNzQ+CSV7o
r6tVZd7WzTgLb3EE/j8+e1UhpkazdSk1w9uuttD1TL+Vw0K0GC+EpI55L7wMzU6M3KXj1uBuqVpE
B+chZSMqI4gjfiWky5VAbsumypCTMCKO0bpJjDMhQvWpCpZHUkhctHOm2jklJZTIRGXsz7jpSK5B
OIB3OOGh+kLqLD2LUXLbaOEOWnBsGh4+Iq1OI9LjC+HBCGYZd9rioe9EXidncxfJ6Icv0z6hCf0H
MUaixuuaBcgf2527caZGKWRcKHuupCKzPcXzu9oluk0cLptpauKGvrTd99BAsrXixVfcDNviyv0f
EVxoLRQg37oR2qfyQ9+BVzaSBosHubIVnBdmrGmgPhna76fHjaOHQ2SFPE74cXn89M5HsjghyWTv
acDE1uwadVDDDXAB8SkS9RFP+PfCSEaKoE/eb9Lb4Ye2s2ym1uhIHtCBkd24AAGZB94ncsGBXAQ8
S2RucPQu6vJdK4R9pAQDq0tDrd/PIxb1RSgREFa+dx0jDdA97MCrvb3j3CkSCCB4Bf5HVCXFa/bX
Tf/beFlIVw/IpFia4yiqwIAx/4yJUeKd7WD7UqPKxemSTEj1zLQFYuw8o541l8rXdeT9QYgEfj/9
pqEbiakSpkU1yVoHJ3Urq0X7jrWZrlfU0M1SApniC6tKjfJcivmYtDRhsaaDsgtVY+pDvttXZn6E
fAPmoI3+gZTH+p2/UNcx8rgW3NDWmlmJ5JqKcswfocm/SdIfNRBYY3o4Z91Mg9GAsnTa/uae3eAJ
y5+8Fr0NIqrq7xuZ7DoSmZkNca4nMKb0Gv2YpvZrz9A9SvYVoNIo9vj0FvsFMyjOezZAJufc8mhH
v5okU07FeG4EA2mASjVO+OwQRxB7yO9IW/7W9Bz79P0tEuWb5FVnXuy8ofgsjHOaeXZK8UHewBJD
tyE1XVaBP9farP6+7cdJhlaCx8jQ8YM27gLlf/2Yie7RjHmesHyJSpyO/Fk9bek0lA/w7SzEemCf
dmQcHhnQRhM/KpPKhMLKX8qZYqLGrXkB/sGXSjceCysWI/pH0iKlXT9nzvxEcTsQG08QW+tLyzfT
kqLnMXqP42BKcQcY1myySTgVc3Zv6LVktWvzXcHfr3+jDZaUoELxbHF6T7ph3ky+SVx00PezvSLo
DU/4ra5wMpN7XHaKB9M+Omm7dSF3uJN6aNSgaq+trqLIqtb3fWBM6TtWOLaG4FmslPLnAdPAquSa
zuer6pmuvYclYfLWRTyfo2510j/AlFoVpMdHeoByENtgj+CUaIL6fOqRSl/3SFssS9BKvFw1coKl
G0Y9CBjEWyXsG6vhcM0LfdS+x2aGFR6x2Hkf+pgV9n2u7eAYnAUYONJOuqGaxl1BojjobPaAWsgr
XySS4TqLfTWcABjARa0vHKlPwJsmBPSHxf0cEmamGDO/xMBa85+W0Vj01R3wqdASYh47QowZ5c/8
6cOc1GtH2bTUVoO+1HombHMR6thmuzdUtgEGKRYTT+q7etCVmV1s/dTYGaNj9hIp8eLrdS015WfR
gzsHAHfH17liZFj5+7PRyBFoG8u5g1DYBRuhL2WPn0ErZEP0i0HwYzmLeB/6jPePVJmJjalJYJNB
z0X5R+u+YXZtrF72r9n/wYDLNv3mKxq37t/B/+1bP75LDmRwq9iqrQDOp6DQOL84qzrFUT2vkqFg
yjmkPtAzFsNTozyC6lpxk2nE75PmFXL/NrWlG1lO/rD46OmHKkGi5eHtSESSRrNFooLBMro8FGMl
CJF/tTkMEeVvjLW3lq6Y0vhfGxtv3McDwwxf+DyDkx6W8XTflxz5CS++YxbAgcxm5u+N+/FM8n5g
70hraJalzbgPlAChCln7MOYL0vJbX0gU7VrT/Hqew6WCfxTrysQ6Bsr+SqxKt+s/Svemt+FFSnkd
zA8yMr6l1CLU5kKlhoXlRfZYEth5r7ZnmrWEthbqpg/yAgSkxIarkWxvfr3UZgCsYaBcWWAvYUVF
6NhqncwHJ1fwsSQv0YJ5b3AOsKfegTDEVsnqg0je4b0aSh6BeR0MNOnzxGj2pNtlQdn4X7Ibqnx4
KZD5wh4qg7JIMMivk++fKfxuPgE+IZj/HqGyHF2rBMV+J8+KyO1Tjzv+hg2qOpa9rP48w3DTkYE5
kroGl7EzkXyHx0osrslOS5kRTb1/RFxv5Sj7lHtfA23b4zbHOJFx6JzTnnWpiAcXUFk0iH4siWl+
mbj6jlmS3/OCydVz0aKufVT0pqXEaOTyW6asCzqaafLkrBeHSaR8NFbyvdhB0773U1vBl1QlgZBu
wg5xGrGv5nUMKjZIClkwHm8eGXNZPJ8EMKS4h0lb2nsBxgVMceD2jjS0ZS+PkdUy5Lj6LxB2GORQ
YQQcJrfkHQL07YWBpqVRv/tDbputKhVs547X/G9XSLkc8bd1b92UxWc1JzEyhTujldtHLBJW/nK7
BhXi+6Vllarutv0P9r/VKdykY9rTp2Qfs8ZLo0t0r5HHTNIuBiwTS5RBjTgUaW8QTNR2HyjEKi3o
Li+v8uel30mI5xjytSZI54IGPwInLUq6YBTcyXlXB9jLcCu5zh5p0hWOaTkGnPbUYz5CgJI8H7+x
OaJ7FExweS7EQ5oEfkhNUSEePR7k3twGaZbvjCItUhcMaQ4H1km4PD3BzgiLb5IBybduACQjWUPH
tANiwnP18TI07jphMDc4NbnGpFfrbLG2YPM9eYo6AAKeB9vKIxXvFB38yyjhyd9F03bN7QmbTbLH
j2vU/zq5yD+ZpbPuTKTlljZyGZM2+96TUuYfYA/M388J5VMegy3JbOKE6SfXE+euegy4hFBwGEi8
stlPxCytM+ZBIEaW9FQrLa/X2DtgstrOaAEeqM5v1ydCK5WUu8gaEJwHXXlzdLmPU1s2Bq9WKa0c
G2XVIVBeTxY3RtmV0lLo32RnZtKJk7qD8Vu0u4Ysdd5qEWDVXDq2YHSzzwrW7+IiUk8caP0nVHWk
pxvcfRLuBAMtxdTlOoZemPXTlQMZtYjmpmWCkpF+uTk84v9XgM4sQWkD5wedCbWmjIzlfl/Civx4
E6sMrHear+Zc3PsCYn5e0IXllhsktNVJmd9BN4sLaI4Cf0G1EjhfZJpa0guyH6AF9Ew27D8il3v9
3TIhPI5ob/KlpzVEt3NCRlGnsJQZ9ds8Chyd1X5vnPRLTT/mlCUXM0k4EyF/Fzu0l/P83JFU/qa3
SoQ0DSMVEa+mjLP17GLFBcRFTsVCaDHBodJqQ8uZJi/6/+uUsv+uYWnAlPzGJ3+pP4AUaRhar5bz
9OD3+0DXaRZlQ/FZBae9tmvQZOnfGx0BKzP8HNCTIntWdg+1Bqki5lWEFFaGTu2Q/nAinW5jHiwO
G4LjDnycJi4r2MuKMgc7og3U0r02yYzDeQ9N5TbKyszkUksIVvI+NoWIZVSqK57D1ZbLzkXjGQlQ
96KV333siYR7jvTc2FTYtQojO/XtVI28tc478NhguHoOUoR+QmQj0O3emhlVWZhvzL6K6ZgaANY5
WmvXf70YeJqsof3y0D9vDWFM7DIYWo0IAdZAf0ReM126LmaNbtZohXIdj6FJqmICxhcx0YWYiQt6
QJGrXDaUJ4/GpyR2vdEOcB4FcBctPMrTVKjynGB9ffQnPf8tWVOj/SfoAt/KPC+IJAxV1VpAqI/8
aOukrY7E64tAPk71LCLiX5VzWbg1sFlIEkRVAzmaD9eex+4tifhN4QvLX9thmOiQXVazG4qYv3uW
iQBRAhCzuL3gwmMFOgh2CA+swcBhay1B1ACGMPPZapNui0jOMqOB/m6kuqY4dBG+Un1GlshdsOXV
vi67SiWag+z2M8o5gXImVrXa6W7ZDlmGU+gdyseqpuPfyVrJJNwtc9vOGJMoM0T7JKitwQ1uFpdP
0TCRdysHKt7YANSFcoFHxshIDOFFa/1UZeXkRn+A+wF9akcrmPn0MNVQC/3StjGDJEsqn4DZw3J5
KRd8fYxC52AZ6fyH2VvlDRusL3zDMEJ6morX8eOn7om0XqlAQMrkLysVY+/F595Ewx/zrJFTVgD9
g9pHmyNJuhlXaBtWLnVAHVsNfSZvEpSBCJCAJwfTv9CsKphD4di5zbvtUuF7mrbEeWUgMDiINrbP
py3i8cm4zmbDmilgZiI/JRoyHNF1Ooq0NPbxO/s+d9/vkcByne+yKMR5Rhq7ZN/cuS/XoISKB2/5
NNFAr8DjfkpYFqkXfduAtwZ65dkWfW8rGnGPVe8Wpoy4/mPV1kaj16ue6hfN5VsvfwG1JAO5kvLC
DcvqhdPMtUjD2nrHsqO/ATB6de8FzwOUGgkiPJAWywQr8EQ//dOwhxZLOX+sjAmJhj+GIjHL9fkB
XKzgazogvqSyWARBmqqHHdWs4/+XyY0NJQJlly16f4BamZrNRCubx3l+TNjThVDYjAoj8tOG2eeX
rG1lcvMfO8bEWViUnhnvdLWHMpgQ98y8vmwjZ3Zsm5ZS21dnIabloN63djdIjzqzeo12MsybI8sG
O77pYMX0tTxfuzWvcOq1rISJwyLDYiPLURd3MfnfaYq87npfR4CjodM9MGtfNETOJWp65VaM3qz0
5wfSOgbHRG/HsifvB5xkmuvPSUwlAha7ysS/wkPcSBSrXNGIGe2/s0NVjH2qR6eslOI8kDyXBgJ2
zaYxAx0Ulz8b5ze9iWJx7/xOJVa4J0QKv28IFZqYsIEk+/lGyKzdc2BHi336PKdppvtpml89I77g
2Ly20kkfeufIIF2vGPDIyBFZbhOLfMAH1nKYSyVjilupq/xxW7umSIJUs4uCVilk28/OI6ewPUao
8Qe8zlTA1tZ/N+cpqMZ7s5Xe8SZfHf+yZNDLrQkxV0RVN+dxj9/UC1aB5/q+zDwNsiz4jP44Gf9h
LM0mINs225pNugP7HeRbSprWzbUrFql2f5uF5th3fMCfvU/LZa6dtFTE611ps7+mXhEV8tOMg7Qp
Qmca0laO347vUhldjv5K1AN4PcinQIz9fuNmwjU5kLJlyL8CGLTGlYLbZt6cXkgiLVevHShxb+dm
jufz3xrO0gdEfEjns4Qx/m840wN+/q9MIC2VP8cujRSEK/kLpD2HKe51Lj7zAYHLoZ56jyKzknfW
ZJPZi35GEDKyxc38tbcbtc8g0kQq/YEwXuLuF5XLf3UwRopwetfRZp3eAn70q2y0aSXS8U3wdb75
4AGeo83IPWsRPEZtiiH+dMS5chRhbd6sHy/WOHOs2l1CdT/+HXKEwIGqim/dm0vyn5+WtFxnFuJY
U18XlvIvbKK1oOUKLLJcnNJ3GmrtaHPiU9SRVP87f7VXHcZoOPj2BVdvR0IBxfGgtrfrrcfcb3Ru
p6MsL4CWWyiUAbfK7MoeEPb/pa32ThM3kBSGqycFAoONVJFs7vGZtaLJZyQHVRtQ8AC8fZ2CMgoc
PSv4GrsdJvwHN8lNwUldVee7KifDmwc5Tv3nOFSPgEWIrmXyO7v3tAXIAYN/jxGwfSyC5jG8p/5V
iTx32RTqcF05CS0FTPHC/Eo/O7D9rLcxi1uWuL/vfWocVaQq2LAE3MnNG/9aPn16sBgVt3/CEHHP
fkezd2ba4gjDCy5zflY0fyXzgCfzuudkwRuepWs0PKo0sL4couoOdxwSSU6X2yQPTeXgvbaU/9do
LcC5Mk0jWxj/yOByE92d9q4P1NQ3Gg/l6oRg45dgSQC7nxZeJJeKnd2p0R96nSyGjMoZRjCF7PjQ
loifsTzXo6KV4fhWUmXpQZT/2EURt6Tj2qfcA3iz3XJKFXXWUbaSogDFUgOykv6d2/Bi/5h9XTH/
KX7fAD2fsQmbkQPuS3rTp/T0hwz1IRGmExj5bAivefPE7ExYy7+Lv3R+P6MUFvvrizwE5Oynclu2
woFepV6f74jL6/XBdRgTNtsm+OyKqOJOLZKIQmg6lSJ+lsDrRWDKi81r+l+vb7aNV+JQr67wqHF8
qjuI9UoHi3ADZ1UUw7FPROdo31xrJmIHLgvqGHxAFmgqTZ3Qye0cwqvXqBlMaR2w1yAkhT+uJWS7
DMniBs2oG8pkWE456VMHHw4pQ99jSKwhTmdApQ7o8Ys1O3FgWEEVdf+KAvLsLcwAKNbhyjmnKXsC
0X9S4GCBCZGWLKboXRmxVt9KO7QMQt6yc8PCHa8yhLe7yNXgYTyPnIJAhchvDhkHSOkhLDeW0aXc
YmRIkMLE9/+ajUcJ5soN/Nh9iBhri1/gE5xx4jwF1CM5LrVSg+DnksLWwDTq1ZKK4OJ5VVFml5qV
xzHJyvAhPpa/C+jB2+jHc8BHbBhe8YEwikcVnss9WYua0naRCNej4XuG3hg6Fg4krEX00+e9u4cG
ogPeMJzuAdgiTk9KiOHHFtgrOZY7dz3yWl7Nh8PiWo+Tr3Jsan0gGShOPLlEi7ZwLyHWIapy9a0g
GbtsxFqOGODX/65UIgqmLODj1DOm1bX4wtKo6YYNh4EjWeo1omMjw61+Ek+FI7lKmS7cK1bqTTFM
x6McW5pQmFGw4qTfbjF83zkXOYk5yAtgjKJP3m/ZX88VeaytWxLcMWCSyfeGkVo9cT8U0wfJG97i
9g3sYlACLXJvSb0spOP4C8wynyDBDi0IVfOANV6hat0OKCxm93vwkcWbIVL+YOljGw83FHjtFLrV
Fmi8IsF4Y+qUblWDs2ynfw5JA9vM8wrLn6UGiIeRaaHfUqAROVJO418cndWIyFSXbMB6FCM3/kz1
R9x/mpN3t2y57n3ZfUbrXbAhtfpLCxcWt1w5izoKMcJaGrbTuoCtnLedecTTTgC91FkUUA9XZcII
tO+Mfo+wRjV7gK0XeCAb98JiN4SeCwTl3ecKad3hs7ULS2tWX0czq5cA8C6qODPCvzyHfI4fyIpL
/DLg0BddiWsv8jJ9KHXd6ngBfw4Tnxbkh2nRAvtqafiCvHb/l/VD38ybJVEao3yrdGb4vkWJCwCA
IHb2upobbJiAlpEmIxIxSJLAzi6tfoIYVX8h5COjNqn/tB2fhl2RZ2t9jk+MPo3nIazteFDvDnTa
1Mt/y4ZBB4UkjLd94FMnzfgmXmoSn0QPabX6lRtV+LPA5jhvl7wsbsY3uQL4WFVt1u6D7WQV95Zi
kxT+CDKQ7L/QCsdEJ1mQA0dYaSo/e6qLC66uBAUbr7t3ubdWwNKjjNeTnf2D5pgAUMAguIuYHOW5
lFcqyH54dghBRqDBnS3xrYZDbNqtYX4wYFOD1D+jCHx2RMeVF3HJKZkb91vVgP/lbMuHR6y/6pxk
AxV+IscKfLyb0Yh3DdIGWy2+k0TMA7ESIheoV6HyZKVMcSANeBKHVylimsegxArS2I7xl39rtycB
r0oYIjhvw23P5gkvowjHOkD3+Oglu1wdSNte1CfC6tFCRnccAM8Oz2U8QOZAUX5z293FWun9/zC1
daxKcYosgg5NuMEpArrGbjup5itXUlZ068Al5oAJlmV3aWBQUHio76PzAjN1AVRZsmg7REEyPLSA
E1hvkhCBJQaM44pQH9lwWTlY4S6exR+VzoMX3GA1GtTiOYh0eMRjDaLFMsuOYM2A6Rg4rccPk/4K
EJV/fBW40ZjDFeqeyk4pZ2xaOqefutSQ3JdyMtA2JhNqmI6U7fWROb140qTbXFrh+lp33JRfswCT
6izrjp980mbPXVw2a12PDZAVXWm5DLtOi06JVQGBWFHh+efD3MbO6Pi8PGFGJ1+eiSFslZvXdUvv
gfuXnzYJVAheAc25faZEfiljEg4enn7JvUWcDlvNuwUPdZ9dB2P7oi2ujnyG+qA9GanGoJUFibNv
+TBmfwp3P1lrdaFxqddlyEs0chvIWLqWZBKU5+Yel+MHl3Kh3xRfwRwwwIc8A3D/C3D7r3cYDFyL
08epUHYOcs/FaeWc5b4ursJXsbTDCBMsGdkapHJr9wb/UJdK1RLDWYgIA0dq4F7boHkfkdYjXRr/
6yaTNOCgosi2MUgyTk+1fhcPk9ghn6DZvEoFcGdYGFMhLUnZePRTQ6ak+DQ8dRIIlKly86PlXk76
Sv37PGLqHtswGKwUy3N3mwk6aKIDNkNER0RcVbvd5PxG83wEdFeHz/2+oGzwUBFqcGFSZfVSqElk
kuxgxfdPYXFh8mdD6h5fklvKwWlB7Rde4trevVAL6+tL36w4YsLh8Dz7OdvdhFPoj2lqF5P7Vg5q
uAqaM3YebTYpoNjsIDmfcwGpPWmisTvaXYyAi5lEm5ahe7EjiBczK8N7T/tysJuazBNBV+u4rM7o
aqI8BwyyWnn2atHxWklMSJjD/nOx0tmznfX52g4fr7dFn0Oi8bhuh3vf+UTChd7LPGW/lZe5DTWG
7KV80nLSWOMZ3tJQjUJRZFudY9Q4IMrEE2ihF3QM9wo8ki/DLKiEL1pst+b/g3TXzAtGudLeCC5s
Sd4xlW8/pz9q2QY2q1iSXlEmHMjN/LnZruj4YravK9JugvEzD9sqLyq4R0meth8lqdZkkFyI6qG+
GPs3Y2o9E3OeWYZJQGhE37nJPv4tWmZu+ximRZdiieYt2A+Cm2C7KK/WVZUyEOtbNn4sD2FjG5Dr
tug7ccRgdxtC3T4GQEUZ1Tr3b+zIf4xMDy40Fem+YllKR3Csx+6EA0JecRPSdEG8rjWrmiiwD0Bd
7EVKPa0A3O50WN70bPf3BAd+fupNUkzKyibfsaklk/HMBz1hLAxyFzcFH5XYeazigtUDzzlHrAIj
nEI400P+cnjqWtAqIiCl/ONHaCsZI27xXl5kqFAZVYuYgh9QR23AfeRTk/9xe8cbsgMLu2bCrDzf
RCKaDN7Q72WIGJxQJvCGzx5zgw7U5GmvPJY46de0/Yz1knD106yHXx1waUcNhV5CinYTfs0h9gld
yOYxWu9Qd+q82yZOCgRAHK2ibd/napGfYHG7GvVay8HBq/iZI9oTT6TM8RTb1orPNi+CxKt53JPf
Dab15ZhatM7WumipLRtt510Yx8voaVmhCYVZQtnZRGPwpSIy3wZoxYJw9hyisLc2GzvKgHCJgwD4
KFAsmbQ2eJ35SSFE/swWBOFWNkkA7MZyHV+yH4g48lSgPk5cptKMlHCfgDcggW/FwgxRJzx6KYiF
s/NE8toipPrGKAJ3siopDNuIYcsTF/XoFOX120CWK0IHqg4qgpoNjcvfecmaDT20FjEONqCvc+bD
TPQaQihF3fLdu405IFaPFFUYV4fHweqsHari2rk9t0YsqyP2eCWvb+wzSV6T4pVFNOGfVp59zLHT
E3ef5pnSecxL482pELlFp9R9oyG95cEWV3329Lp5nmmVqqSRIIoc1qahM+uzwYpxmyJNZrYPVfpC
8IeYiR1Lm8O9tSwFbxfms8Qx/6LxKhstSiGGo76E0gBYgytTIqQCz0TluFAuxQVFFCRg5izHJi+Y
bok9iivpCC86Imw5MEcxceufuGr1uUSz/xGiJSxd+9TDkz82Gw/bw8gbfEMYDNyk8NO03Yj7q9Ra
DZyHbAnhCT36D0WZYHEi+oS/9d57F1EjNhozpxuQSga0t421VkEqf/DQkGHbCSDq7UuC2Fh8Rxds
VcdgmO0CXcK62HZiVpzKVa9DmTOjvLNp1xYpQwUXMJJH7/telGuLIC5i4Cx570dfKI+hPhAORa+j
CPMV9YDCoiDQ1AhWgP89o7Y+LISaByGoso8mSL7Gx7VsINNZdGkasSK61og3NzfPmvmgCUhBdMfT
5f/SrqkromzPQKuJCIbwSDeZy0YIa/mo53IjVlQaHNPhx5Ge2RT9yBZod7s0nssVEt97AZhbVMr/
atlrDAyPSpCYE2Fn+bceD9ZhODxnBIusUF/pG5RhAGDL5ZsT+5NEZa0tfiqAxFPLV8Zlv5C2q6af
cbRjrjsWoN4pEMnzzzaG+KMAg4TaFnzBjIU0uOEinfYHTL5/gZFVRUt1Od6Z5B2RZnP1DPNASS7E
u4yKNrfQVZ9wyDSyChy1uhLOD9ZL6SnkknqHRqseYFN7/GeRY/fVp5YFuWgS2wYsu3YwB3K2F68o
aYH2lUenGqOHaLhxwm1Z8Z/rwCdQTrLBMMO57Xs3eTgxfDbBzI8BPUjX8f5D8zboPco6BDtLMRB/
lmxJIG8sTKgpbJpV+wvGfseH72JMMPCnisOAo6XZ7j+i3e9Jn15UAW7M4SsHBqXw+1RSI4ewBoFW
ymbnKl6GAp2lTPc756aaRi1vzG/swisVxJXysTLjaFpejDGScxSlbkwSBxbBEiUUbK72Kfh6SeHp
/fM4lAIeSFaoi8apr7ik9ZSOwgE/kvljDSjW74XC42RxW93ja3LfbSMlJaShqPIWOaRIu/+EuycY
IBP5/6gI69FJs4ehiXpzenDufiqDsd736esFUYJrAvN5OQbFLGalhI6xqFz22LT6/ir6QXNB/d7n
avtBm7Ob6uKBN+b3WFxYbjf9VAX+1mHofW4poAdb+rPVIHT+vVEWU535Y6W7Apj1Xb84/wkfEsIi
oEKRIdEmAJIXImR1b36vIXdnpXXhAoFCdL8VWA/czRq5cvM4QXSbWybuPvzCndVSmyAIeYQwIWQP
6c4vgHdcdmXlciN4bfVH+hXvfZSQmfQYpOBqW06XOhpvrD/lJOLAMTUXHx7w9+uzMf2gVWdDUrI7
xiyAO9pfI4wHJ2P6DKH5az/ahSYo76xNhsb+rFelLDMGPD/Q5sUIWBA3g/O/cxidtDeIIwZj3cXW
xEMRy9EAtVCPsZfF8xWhGW6nvEFqnNuslm0E9ZUWsNie1+Jz30LGoDMDKexUj+XVNVFJDwQr6ila
4AxPvWPn9MEkyuKLPqd7OGhNQT0G3c+62HMeg07LhZHzFpTgXeT41Ea/ZbLJSiyO41EY3aNJA+/r
INd8PmFY1tfWEl2lLUmuprpc7jRcR1QdrP1cevfFsLG4HEeiMIymHechR8pdKPUW0U44s3vlvAne
uNxzMLU7HoXl6tKx8QFZ8Wh3SMRXp7dCGVpUXkV350ZleO2gD424oDI+t7MRa7E9ze/Q9xw50vaz
hZGLDwx21zdH6TY/TArBq8Wbkdxy1hWTuh1gzp6YoABahCAHiaPJ7VN+SFHbxgeVsFm5wDeEE2dU
0T+TlAk8/i5sNpECpkb2+EKWldQAbQnXXObtQ9+8d4ptiK36AUpUyU0mC9MvsYZtpOEwmBAFoiVZ
9PRTxXjRfR2PZFQphk/ylnAVbWWoAqjkU9++AOsgeH89juQm0o5igt2aMDR1wRm8IEnK7KoPA/07
pODKL9oRr3xMnGHAXdvfAfYbOuxyV41Hwf9u0dv9co7/zKXCvxheGNrGBaw1u1FqB52waq1V2/ek
5fx9jZ1GLvnnP+xSV7K/r+edY/R80IS1qgMlhhKgOYHVwmnq++tRHc42FeH2JRgksAwyZjzqt9ho
gfDbAeNs5wFniUcjdJ1LNgc3l5asFBqXF0/GKU5oKFnD9HOV7rzU1nsE0UuiWysWK61YCVGyP/nm
EwxK6MFmSEbaXY0IgWe2KZR1ApEpbyr53Xvtsc1yc8Il3sSgOVwLBmdilqM/5ibJFA8ngMfUGQb6
S2RehgptKDz7jTWIigXmJFGhz+Wdo4A+FObqyTQH4f+hOJdfSbVGz4HuQkNENRccyxjBp+EivEK7
+9+Om0+B7iXq3juHnpYR8AP9sU0Lb2R95/+2feMFJKyWzi6rtDyysLBMtG0O1hyCR2Qncj/7SccQ
68ndN0e5Nmw3pqXEXWLteUEmCP/ra4ThKRwaqgU7zxqF4qEPAjHBk5J1GH2E1jf5nK6oAXmHW3RH
cCLF4SY9IARO/sSMaxVDon7HexiA4Le/WW7CWpg5GmmWTuziYNL+eUOM/0az73ufY1WQr6jgTg5p
7M1skA6o+G8Tc0jcxB7h2BnI2PX0OG2TBlZqRg6bhK1GP0dzXgr+7LvtMyug/cz9s5z5vIWGg9NE
p8ZT0rKwe+BxMt0XvPl8im0CxkinTrT3TFJGJz4ovkilaFHu0YSUG7wktJ8pwmc5zDKtjEVn+fqz
j2rGeR/OrMGxRFALnQyBPLEjT1gof8+Ap2rZcuPH+69y4w6gXlxX4EBWY19KUFvqZt70CyIddd3i
gmJX5sURL1tVw+rvEh6uc2parJqCHKT7gEotgrNvNl+o1Ff6xI3R9cEFh3IFehZ/w2d+6Smk7nzs
Pf0zPcjEqB2cGGQmiVFqRil4APBgWlfobRADxImG4jdI+z7W+UtR+tKLgEyQNrVeBzmGwyI0COAN
BigzHO394LEhm3GBGO2CyMttP3Lmdl+KmDz2PEMVhmYw+ve+nQDA3FnIJM/KxPaabaLpWMnb5I8z
n7OQiiAvcUaaXgHuehL+t87pqEKoCC/8LL7YPiur4jhs3tco+gg2xl6gd/DABtpmLDr2qFKiMN5M
2oFD834ZUEtoh8B4x6MKwiqkZ1tgvANeEhpKw/jGyEizLugO4d+YLapa/1Vq6fsFvBGHkQ82qx7Y
XuiLjH8NBHWQOc6psyrC1unGDsE4fWFySK3s1C/ErMfFUPOyjp4Jou6rm2/sr4M0yOoj2Z5H92Kr
o7ROitwBathUN6Qz6XH59jZh5qhZIUvSBJ87K0Yi7KZGsajw+d8A1iGlg7XYM4Pm1n8OboqRtfW5
1Bwsl6XNDD3ljhDgfFoJwSNons/YW0pnF1SCG0LLcqE+G/Q7yUzvmwa88HF2ru0u5HHWyJRl84Gf
F37MN6+/gtukyCfTHnep5JCNCcFsT+ndB79896Snp3OO66FqMmDv97o8cskAI9lj3ZsTrrEGqHCT
ibaRuRH14oehHmF4C/5KTYfshWkTSeKNOELBIB7AIIYjM3LJ9/SV7lpj86yNdFcdUZGJH2/+rxSQ
HPwuqwKj0bPtPIk0KRhI9+39CtpVl69DKy4jztFJ0kQw+4+OP8QMlIbsSCDP5q10Do040ksBhgPg
UpWrIwFtIq3vQejsrw5ttilEUX/MSGV9WTjKONTeqIgg1w4v6Sb9P0ToT8srngYYyLHkGRl5/+f9
J/OfCVUJe4ezR9k02kK1AHX/3RzQ0TU0gUTRKM+CyrH7MDMoID/u6zd6TSb4IT+cD0jO9lrwq/b6
wIJ3T2fpIklom7ScAnlwk7ObdPya4TTRXm63LK62+mhDTnV5VQ0ygTNKnwDdeMEb05dseK+hpuAi
6PLJ0D+iUj9iLdTeCT6eEVpFFD7+N1Mbi9jPk31vfifB/RDMuwQ7M5ZoQUasvh8Nvbf8d2XW3MAD
mDgYT9DQj2JEQCgcfwspmiUlegT3YwcyP/2t6jQ4v94vrjHL+4iSMyU7ZXQHvN93WagV2WwW3bmp
rybX/IBLCLNzcQgAkGNAHwfRk4iOduGLwPPgSzfCAPP1/Yq0iQVNHIQj+p+z463WiGpopIHrQK/o
NH008jHA/yz019pH5wKCiIw7wVdhJ8Ft1pj9/TCZgMt9ZqGXLoUhoOfgTR7G3bnGKvNQ+igpSG8f
aunzbAyeJw/Q25jbGXU2KycNwWWRM0TWXdePdxZ1SdAe0OIb2YUfB/HJLoD04/NCT1we3eYg+nAD
8HvL75ajt5esBeJQi38S1Yu46mSgojp9aMB6wOQD7X6CXUx2Tuvo/IzZjyne2ffsRCm25PLHgo8B
/yxIqDPrQ14bU5znxzFxCH7NqcRdecjIZo069L4qb0n7/BQ+azD/PEesJBOOg1oCqLjkxlOQc7ZK
3URLIhzeRcTwt9WlvoXiKLIVuChG+b2g37M8L5gWBW9vdNExdAl/8dcprx91pD8ZPUm4XeTeJD71
cxfRs5ZQWD8aHf1xIdCG4G6Y/HYB86OcIBPXQ6Y+EQGxHX28SRGL7I1kZQGhkOiiEUqfUUg/ACI3
094rjJdh3xX/2aZepE6MiRXK+O6YHVNNxRnDYYA9GRwpdb6YiI9QCHw0cg21D0Wq+dErp4mu3U2U
Mb8B86eshqTvH9k/ejGQfKeE4Q/inb8ZqdLlkd5KAoJLeqe0UKZaVcog4OQ8+ZDf4Hh0yyRP3+i+
xSNsu/i4mB/FOmnGnGN5UdnfEFcIZ+vZci9qkyPXGmUI21pE0iLh3b9c7OfuxzYAf61kIJZY1WvL
HQyZCIDTNyqxCXbdgm/QpEW2f4NXSy4gxPZl08GUoAnNnd29YeRmPSvdiL6wDZfqK5cFYOcCDcCQ
lDweiJ/qAlQ7FMx+c6RM7GjmJ772uWdJfdCgTpIOmnO7zJriKibNZgFx2v7MIznIVvO5Ghekzomu
5GsvQgBmrcgp0L+HaFcTS4QxUjV0jt/QOtm4Ye9gqlt31D8tubY81Ud7IvBCWwRuukwY7BhMwWqN
7Q6LNeJcoRil9302x4iQkfjCf1EYVAvqY5SGeqsnxsSG1CEIeYyOF23tDAe7/PCUA5TNh96DBcPY
w235zLvbUd3AtkoxNIo/L7OOEOKWUKnpN/4GAGuXe2bd+KsFfRfqvjAGXDDFvl3WBuaIHgyL0ily
bHAlzWfaw2WduH8CxGRlMrAti7fmV9U07pOuUUts0YDlhs2qqy8VvuUMNaSJSiT02i90Aw65Fh0k
5KG8Ji54dMCmSn/5zJ90bqobuJ6oCpvBFHzSsCfpMsw7CT/FRn9LGm3MJLtX4wxlkBzEOPpej0ma
MWwkmYEuXQrv7J6MESgCiUivxaaEJlwmrc6eYXs91XIqqcDOqhOXj+lfOK6aX4bezlDtdcnbOZhG
SU1JBVVxbOtLytZCvB+4RNGv3kyhwSzWalGIvJpjl98PGBP0SQKwVIWoHV+0GzyTFLjUUrJRdkAv
RAWFJvliUNBTFL1U3pX3wFij/ViPiRqmSrGmBEtvdsDOzbwOXgd+xacJjM7pbxoDvRzwn6T/BFbD
kuz9gRCc4fL9FbZBvEnqMQm2HU9FA4+2p7J45kKTWZ7D0bAmDUC4NsBkqPcV6DIow87pHHQuP3h8
qKsbro+/xdVY6wRCZqXB1gbWNZ3Dxm8D5BhdqLKsL5zoc/1x+ZemL7mDUnmBCW2g0FvZ/yi5eBoI
mjBzzh+RhHYp2F5xjAWPLtY34C6HBSfrH5mL3yvqAiBjjTOFLBoyzx794TllmoBVFt75rgPFpd1J
7oe45WmUZntUbPSWXaFCEBmEiFwF0U3zwjg2dV6WIA+K9p4STTNBY59rxh4LqMsa2GBxWJXzzIEU
c1Tou6w/Hg8mi8dSezWz6tGUKukFt8PdwTFHF7A+kPNHpIX+UbxtKrJsodY4mKwc3ckwRBqgr4/F
BAMgMkLklWs3AnW3HBGbR5MS5D1fCuk+siC1HiqAJBHojC/jfPi7dC0hCA31LqfjeyuECLUgB9nH
OK1dw+wxIBJakGYmfm17nAsLklooX33vgBZPZOJ+GXzTRsNse5igOoWPR2JRRQPRgDJHcnx5lGSN
lxpdOEAEHmcd0gIwbCbTifqlyHl5JiQ5IwE2UH1Og56BjKuLSFVtzbvNTe773XX6ctx7sgyNrO1T
OVofovJHebYf1Tr7MZV/xJaPdeLXhO7weJMNfrx0IAdIyHITa9j//lqIJUZjE6Ez8os7KbeC5V62
5AzcGHNb5EIQAifFJrjU4CwKMf86BpxXsWfAgdkgfNLR13cNSBgDwoUe8ITQ++Gx2m3y23dIxSzf
KD+oewTWHCIJ7lkTFpi/njeeffpQa4rAk3Fn+/3OwofPqHbOqFJ7/uuz9XUPr7S07pxr20oq6IhO
3nrgMHtTT2FTutpQNYp+5oITnthnlXZc3ZyC3OQeZywYn+W0NXTmjVhsbUKykC3xyyf9q/X5Kgz6
tyfaO1D3c7JrHmcAIeMeSI0NRo6YoRAJULRi5a/ChV95e3tocg+tl0m/9BqMWmE21km8J6CR5WSA
enBafcGJYX+RmMFzV8aURi6/H6qAqAZn97n6CbNcNtzFHB3doakjECXsmDOCRDLM/tk8aP/gyHIg
9zBBY43nWRYI/UDJZzF7oEBIyaKPSOYMYcrkWP8eNJGnBEg9kZEA7sEgMFegFq5Kw+CaXVU7tlGC
MaxWfd6+Tu0ZCYoJqDjN2Ha59cFA+i8Oz/c5e7TMtRbwoERB4b253lQc2iX4ZlhVLA+zxSXVJiQs
VGkETe0AKsQMW0CPLJtsBjd2+P5BfUJAvYedT8YRUnB20U9eSJTfWc4LMj4BhzR+L+0LDlcES9AD
fVH92ByHARIkoEU8swCvsL2QjFX5POOhW99B3LXJjQa8WeSxA7PIvyRNTD1y1DYlcyWYaoYmsc5q
v/WY74UeDF4SID8Zz7XDtV6Zf2lTBvzrQ5VXJ+esVwBOoF7fynH2mZ3nPl4bmWXfUNvj4Wdk9dIe
xkGUzrOqbr6PpVfjwbUSyy0BzfEh/8YOrb+TJqCR6nCC7ceB90PU2NLmtmdM2YiUpOAm5j6790rJ
+gca0XYWmcW4+VDvC18EVHyURhUBK/93YXYkxAuWE/TI0vee3gBnzBLyHRtVeoWoF7HFRTsobzab
VFvpB/isaq+ncX0x6xPNggJClbJH6zRRmDZ7Qz6P7HnAF1RnF2gwRXbxc93rWvHs7mdjosHQG9LT
MoaujHY0kZa4u74LYqWNaYt+mE/pmUrY9pZyDnVLLLBNOVzjMymMaj/VVI68XlDMiM342jUR6w7x
0czy7xZRZJROIuaooxl6KcOfXSNaWrgsrt2g7Fn/cZPSBSLafqmeQUWqyo9sRKVb66U9TfmdNiuS
vtJ8DKBSj0+Q4ldtYduAGHRDeK8kMWymqIpQ1DmHmIkTCrOZgtRgg82OLukauKQ3RNqFuGIgjwG5
kd5IjxpyRt0+QDcXjUV3PF6XPb/VYVeioQ3bHsoZuv/ajHqYJcVh3UE8KirkIKkqMC8f8vi23Mio
lW6TyVAXqmjgxZlT6+cMMDbztFYEESzwWr44bTzZQFOSmm1jL9eStGdEKF77YOMyvyN/W0xPXqfC
AGWHg9g6HgeBMzR92/a9I8uPvahpq7scARQm8tqX7mVPK001FPUVEH3a0YWGpR8geE4RT3zSxkIf
93Xo/IBc7r/gpm26l2/h/r7nWve4kd00VVg03b9b6rtKVLJpZVj2FTAgW/ooRFHCytFXCQeGVNCy
hIoBER841izH4zt4LbTqcNKKCIxprF1BTOrZUr9erCctYdolOHEGdDDZTaQ/bHJ9JuD7a/MzZL42
/EbUnGGGeOVEyZAIhBIWvmhc8LgqTJUv0CesL5coLWgVbb0dJ3Rr0bGh5ZMay8DgY7+BjmFjgNL1
sjWx792nLOx1BQx/nSbhX4MzK2xG//EtAYkWFptw2i40r+qhvYCrvR5xTiXNMTXEX7VySH6Wj0xU
rA5q4/uSS8nLIQo/nTBYgZtA9cYGHyOqzCMcaZBnYTAvCj4MQtF8SUgs0APHbGJ6QXZ0nnHBMqI/
6mwXn/um2A4Rjmv/o4Y0kLlyFIGtSxqgcmBE3iOg18n27WxmjvteqdjlazZvMgwTFj4PjxclbH8Z
uDYw9BfYLtG55DnSjxWIBXe3J7C2zlPGKi2h2jd650QKYo8vsd+YVvl0cy+kQ1z9pkVurbIj9vG4
ZgbEC5Ftt/wu/ykQ1SKXsaejNF/BQwLWm6CR8a0Yx3oxk0o0EvhgxWisLJSDb5Pp5d88aomsMjTf
JfxgSyh8deDGnQ7OIa92OoS0JJllnp3hESf4UezfigAOWhr4XUK4tIsUDZj2vQv3/L7TQH95oKsO
8THE+VKzJgmVgf/heW08LwQlsaHTIu8lDZpYandfGb4aZAN6OR3KCoCzLdbyFKjo+VVyAYu6Jx9W
mKdrl7Qz15LZQBhOeolcHvZmq8UblcfrNQCYsJqhdHvFvfz16rIQ0BQ15c4qKU/ZoEJvprMkCJ/E
2VW2EKNYusI0bDbGmRVgBXfSYf3bVecM9KiORXfH1g92g3uUpCW5HudRVI3++i6hS698lF3qdCAs
C1fHleYQj0FsM9sV+1V6/01IS7QE260aV9uInc7VO84H5CpY6osi0NIeAdGBQSSvbJ6aof3iqpPX
0Aq8r6bcoQu3TxyHifyF4rglI9DGmP81rW3estAL8+ffabS5sLidg+xISbQuhjkP6+0uRYRINocA
9eZJUJJNslfr3cQ1nf/BX1FKDRYTYvCHigAUph2DAIG08fFOZJITMulE4LO68avw+HG5FQ0/0k3J
9SPFUsJXg4huOTqnH0B9mE+JxUrzXXCeaUpJCOYcK/IGV+4/HebgR1TBRxmXAOEOv1pF1xZHS92b
itNuiyhHy1LDdPprG2b6lLJIY9MEWgzjDl1nHOyoYcrcakw1ubLbMpVq1KFcYtTjTYbVrlmlrPS0
Eb47SkJXH7jUx0JfLHv2iTQrdWBGuA2iHIVDctKbpkJAYWtLnrQuJmShEZi8bMnH5cgxZc5FMefK
lmDp5Q7ceK4lblv7OZoctWXdZP04cS8LUV7aIj+0+shd30CsD1V51GTWQvo2MOgCn+QnSTiBJbaw
8sZw8ufnQSEU043NwmjP2oh6+CJkiRFjoMNGqRMqElc2y00xzPUQH8qJbhRjoePSLxAx5Jw4rbPo
mnkuxQ6QtQWH3ShZMaR3aZpiXOQlqsSEWexlWHvjJ3ozROiU3/0696DRo/KBwJXNH++ExFCZYyEB
3s1qMqZiGfC02u/lRxBvo7pV2b5brHQKGElJvDl51I+MkE8BnIDVT8ZZ0dscTaW91XZ6HU++VR1G
8MK6rT1geKIHwPTW52tPDmVwyhCF/UVTmTq/gojsZjbJPF77qwK+SoKays6G9xXzglkJJ1XNGUu3
aXkVtnmIpRoUu+ocAuhF1939ulnPhN+/ilpIUGqLUNkA5ux3BYr3cAHszzVTjsQHSyOLDEwfA4+c
4ax7Us/eN4rWze7z0WKXP2cODExOA3551Ljtcvtaua/tK6UZzuaT+uamUjmMb75GMlLpwTciCNXK
q9O8hVETmH5Je1yQAY4op6uoC2u0uu0UAhHWXGMwvshX3g7NdLS5zKdNg817Olr5ZATnXbgtSlJ9
gNfX7Q3Kq6W8MuocY365RRu2yjYd3Te9bFl0Kr9kbBjvE6WUxiYqGa5nQjeUEtOahjHE2mZ1pgdy
8Cyt3WIgk0UGUMTu1iHBUXeedRbo2HlrFCYwPcIWHDov4tF1SdYCth0VnYXybXg7QOpwrW086R/y
V03+quwUjP/NdUcaXg7X155x8Z98swzkD9/zjmrjAo0KLofcpGja7ecJKqUAEYk1UpsfpSLXj+/5
vxey6XO5jYot17iH5SRNP9BCpofmgbRdnu+1X5MKSNuGIWa8EoDRutW1r9hOeEf7gCU2vPZ+UBza
WoMPMaF3CtKfMKiIuygkm6g4ATTbCuVcvpb/u21z+mAASg/8AjwpNrOyd2QDg03yiJMM+UZ/Kb1T
h/Iq5SgDDCLf6CLUVL78TxmEiRgFrJapHBE6uZxMyN6k8S+eryJiphLbvqj3nTA12Vx7ll5PY1jO
Ao+wzAn8ZgZ7K8PLIjVXMlEMx9j4dx1qBCkXzFk3CnYGPI38ggu6pj4hf7hj3PWq63L/Da3W6Oov
Q2I0WTpvMskBmEyqFSnFe9onT+wpaJ61KteW7ClaOHfcUcrNFC758X71YPsxCCFy9OTjDHoDEW2b
ypdUcxNJCwUquoxXz2xvbXR4QAq9zj9Agr+DDc2A7h+fZ33FLOH4oOHEl3c03C3RxidoYPKlGxrA
ccGRbL9wZgt5i6cWzsVAu/y3jO/a8kkJnq2EXDbTpLna6kG3+H72XNHxfsyNwCoRVCFrDvzwm4cG
7XUlssZeK2980JqWgLmNtCtrWDt36owZywS/NVdorvZW61wKCM215Yc3h2qqAE/ZPEJNTKHxo6L5
zczlrlsXh/lOfczwyz2ib8+jp5U0SgYHMDRKlImRUys5a1aF1XA3OoOyadKEJ1bVrd/VP2F01BEn
aJXVK8nKN1cF4zB2UN8sJhWzqc1G28edytcx3R3r/CshX9jpg6HjUFczYi2HKUAYQEWk9M+Gj1A/
sP+II8+t6+BKD7BInQBxMDw7+Y8nyPEXsAW+2pnHhxTwQXr5+YqGMyveDOk9rOy8iJndEs6IQ13I
vOIspLDaHVOqhyq22MDPujU7u5C+ZB4ZLr+FLwO9IqM+oxe+bPp9RuD9S2ZVUI9+yZK8bHz/kPPM
shXwsF9+2cdkdI07jlipMBTZ1rgAUyvfKaN6fFyGPhB3VeMh96zUqBGDhcF1SrPeGpSAVDvaA/OD
fJ6MMOsRtZxV7kR6bgfvRVWYCvhU0ppeEkRzeuPcGFu2f3lSwwVbNm+cbm16wCBKu8ipMyDfLWcg
LWXM/rUGwxH/Qx1f0dRyhlKRBtNDkAgxWKzQWIromraOBpe4Dgph64B7+aVsuWYJa6Z5eWv2Th61
dOXY+2X4CHueLVrn9qvkP6s9ULVgx3wPDkKqlp+SfVqeWM59V013iJEHrPzL94d4UAX7NCTeJ+4O
0wS/9Qnf5t3OPlCe8o3FrnZQ4HhV7/cL4BNmZ0rANuXp1spVOFDzzGtc8DyHcoClaYgWiPWVWvIN
KzPtT3b3+8CMk7Bjtog45a62+HIBulBk6cuoCpDCgUGsUDDFV30Zmv21PkJ9F5mk6slCI3bSJXwS
OnQ7VpcKULeabiFk/G6dNMiBLbvo27aJlxzf7LduEuPXFNYtCtsx2zaZgP/wDOA4aVoVS7KidtLt
rJ5MKlQJZcS9EfVtAvVbdMLG37a2Xv5CePzKjJdBuU/5DKGRqcCFf7X8CtrEi0OG8vQTmrBMKUMU
+BbvfRywWccLxmakgLOXjGNNUdyTuF0jt+DEn2ANiqZj4XaFPctqT/z8+XB6dZEhS9Zd+4gkM6OR
hV+OH+T9wn4AJKR1t9s4QfGMBG0SbCMa4934g1Rzq/pKE2vAkf9jwpkU1T+ZW+R1VBrdpd4KK+BC
ii8D8sK9T7iUYN0lnmCp6IHndSHp9MsL9C/dO6M4Fa44oX5fY8pr5wT6+pugOVCrsSeOX4fM9vFt
noJJLB6mIvguCwg1/00dPhSej+yCxdxmB3lofFX4C3EjS2/dCDmH4MeYLsGPYIc0eHgwHuEY/Teo
PGCtqVoPyS9EYbCZ/NvjkEx/l34Cwuy6b0exmAw9wj2PWv372nQf3Rc+kMAP9k2G/sUmjMtNk6NC
11VN7Y3veEaPnF5eZUWPmx3mbdZq6cKPhwKrax9S+LlOxfqA9kMzr+RUewxW2JisFsLQ48bWHtOA
Cx3EBafr+ozBAk3+SPZw7x1qE5Ngf6Z80QBMvGRPGhBU8qkCZpCkvQd2hXE46CPEnrhBNBgWuxLD
fVC+dXZMzc8oyWxDc5oMNf4o/AO3B2Vk5FVJzxTNu0nI5EhvRVReG+8TRgPZIP07OOqkvjRzbt6C
3trpHfhvoRwUMfk5EUevscIJp+L0SCDT+5uZ8HrZhFIs/h/SAOXYMNPoYvIQ0QHjl/CvAcN5m5qx
W7p/xn7xaWsab5ggq/vg6rwMSX4FuMAbhYWbgVlTQjAzTzK5zm+VcBppddSpfPJtGVflKTR5EJn/
PUgoFMSi+i+/DHtbreDnFWtNui46SoFB+r6pno2VN2rxV2x5ps+W11kQATFyhmaYxzmc4Nhle3nK
DSS/WHvJsKBBOgn2pyu2bdkXryvjrKHMByoVaxF1tIAo4TyPYXmF3cHT4BCUK3hUYz+A3Ds3POzP
hEfHdKkUcJrwZXpf2jbiwB1NuoQvfivJl+t6uyzI05dMZNRG6qVaGeygW7K5X1ak6cFX2MJaDBn3
Lm5nfRvw3vpS28P0MnkNPSm5OJzv+r0NEfdQEfG8fyOwYEtWgQUoHT4cE7wxt4byJu0PrrYUewiz
Qf9BxIaVz16FNIJeq0m+GC6w96miCVfYm8duMotb6DHtlF+M7O7jPJpYKhQA8A5Mg/qxQ+RIUSvM
+zWgu0E44jfO4qL9mZ88W0AY2LO4zo5tWTU+4HHlYyAMZr0MBA+yML1tJJeAgc0S71NjLw05sa35
iKmBZ3X1QioBCtDTOVxe46wifTKqMW0SDgEg2KGg0lHDMBAhy24vv2y+cB7Qh9KhekwMj9cSbKKu
vOOOr6wRcyhqdBaZ/S6e4GiT+guRuqUwF3CNBYNrjwv71say7DVvxZInh1wlLNF/azIKUqGHxPLp
HC2ENwaH5IqAX4YeHCgx6keYdcgR7HtTqO+6zxRsisD1DN5lsgVYX3yBlxdLu2xzKtbWh6AKPlOi
DMylVP52xqEqyO9phvI/w5h6HgJKwhzwyRnkYpQSw5mCAWZD6OtyftuCdY+gtJET226OprMzy693
KKedl4Fe4JVtochOEI8NsoGR85wka7bVtHhDgk3xxABZ0/RRWKHw8/VdMlHfRg1zPKHejjjhWC6N
ZjP4Zt6f5wf9bZUwqO6aW6PJ1Y7NpvKITwLHDE55nkuZIXa531Pp7oLg9FkZPzZoEdN2IdgpSs/4
YinrgCtkmHpnnIR3FeFxSvk52lBLTdgHoWVx6tIRuWacwv69jWipWt8YuB2n9O1YMcnUVKCFRYis
WbhTxr/4FxmIxtfKbMlfX8pUvjGho8SARRt7z1W1V5IenCiSQ0lj++mcJ+TD+EdDPk+FDq3//Puj
rQb6k2hXVWhkgBZME5W566+EfhVlzr2ay8UXPsMuBMwf6vOCjToOCgs+My6mklt7X88JZZJ9RBC6
EWTtuuMoQIRhAB4mycQ+S5R1C/JaMLbMny2X4Relqtux4ytPhKRLxfahpknAQrz4cCrKQMUqxtC1
MqKs7p+LU6aMsirx2xe0UPm82ZwIZvZLtHZ6O+Ad5frVeHZnriTsma3pmKoar/i3HgHDHMDbp4vH
9AanZE93s+Hz4TCchVQOT9jgKxTO277Mz1TGESi+d56q2PvKlc8xGza7MsDBX2GS3cfbN2NgNAxq
qNnNX5a8n82qfBZP2ha3SH6QmmOWiZJsyEakkTmzjatyHOX5l4YRY3z+Uo0F/V5uL7ruiDe7CRFD
YLCEGMwoSAWMPwi7SuWOVVSR/KCKTkGthxIXLq5Ip7G3CJwmePACHSYn3KMMi8Y8+h19s4FPYGk9
mBIb6lZ+tEoT/EQU2nqFQOZUgWgjvcflpYWpmM7ny/0kGvL/QI5fwTwwsNmRW33vbLCmwshld/pl
0Eg84EM5iWUuprI9oLIbAX4fKLZ4OmXsSXprXR1Pz7Zljvr3I8D6SkUFbm71k/KNysPC+cWk2CZr
9jBKcJPwYnX+l/iw+YPPqBpJsJBBkCAfUnEIlmPj6lbUB7bezdype5Kw2d8+joH7Fx4tuhRQft3a
m0CGZ4Z+TP/756yByDuSpLF/URdteLMtvEsPYL5jVbr18hf6U2i81ggDhuWIJGEjaHGml3bzm+JJ
Jr0yA1WBU+eiCSLiXY18aNCmaGsur4/2DMC0XAs5uAMJgH6O49vpXdB3OKL2P69fysyHuZ46Qwg6
MPu4qflexck9jmd6pnO9TfLzrXsQM6ezKvsLIVLJAbId7CC6FMjGFPWZOgr1DZXeEBD6pym2lb1Q
0rbhRtOjgsPS4ah2fh1PxmbPpC1fKMyVLJ8/TvYE18Be8x5Jexw8I6kqQXfOANKlR4bU12vn6yB3
nJTACLrQkiC65fKp/HrQPVmYFmUAUwCgns7lCzzrx5K5uyPCrth0LdsdhpDBIlkMPEuwAg5I7Cc5
IoLtyqFxDAKetv4aaWKIl4AxtX2S81w4NcMrj6bhR7elptPQTrr4BX367Q8kV0ovN5VvM+pffkpu
oCMxg00lxmX24y5tXCHo5Ibtj1hqauMBOUcqfsZcvqOnd9f8vuayLM7eGniFXDquiRxy5/MVhigo
JOgFudQB6PoFN02s5ZORb9AHaw/Sq8VUE5QhVph5e5tPdxgtJWjYBUoKjpPrJ9N0K5hQfrdPgNjQ
lLEsoKZQLF2wLLk1yDujmpu9MGBISTTUtiyjhunax8vEWaq3QIFrBafJKFncKidjFdvUYwL5zto5
vcya6XhJWpvk3YQL+2Ch8CGSVOvbU7a8U5VVa4XiPKmn7nYw+ZRw50uOrai9xp7eZG10VA39GmI0
jxwXjFdg/4WI70mwSgEjuEPKttznxFdH2+Fr4IPTDOCinEXfI6q3a8HXytzRWPMPjMPMSi0WpdVn
PsS71knid4LeC5FhEy6ILUDI68D7nR5s2rU4DYkKYg9KS9ZXXlYv/QNVtM51+0VkooO1krXrXKm2
gM41vCpauKvYvrSCk910epM2zbJyELgjkOxld5LF2Pmf0WpVxmNiZvtHm8zrs6whlGomcsD4NL+4
eyx6VI7Jy+kdHMRiBUFMna8mgEVEB1QqMw5mJAs2fz77oHnWR9VzetrX/xfUcl+HxKeIBl1ZbUuc
IodMZbGXho43F9Ixt7E1mihL2cxr9A684iai1XC3An28EFcJAXNCz+6hYJ5biyyQvCrSO6IuHp/a
DTC4j2SSfvCaLA5fCMVAzUcM9NXgXx1f+L+9cepR8w6atjuO0RAG/V1wd88/cVtLwDq3IQleJYfJ
wu3cUx0ldvVa7wYjWhTZqfPIO4E3/GxRXvrq8fZn6zhDqK6l+Cz9yJmsRttQ5w3yRWn7JH1yGw2V
5FS4beNEyyTlQSQytxHqwyyfu3Gqs0CLBBlKGswsvDqqOd9M+jrlA5A6Pl4V3pI+lygMWZuuPr8L
rJObaJqb1oetEI4BrQlNjciZdASPhPILgGTWLQn00ZD/JCvNgwZJzgSqu8pSLrF3bJd7TyfGfQbi
XDiA4okG1ux+Oq3FSLx25+ZV4viy4zBWHZ9zodZGtiYr5fhCponQZ+aGThY7IX2FWVWsPvUZ7DEf
YI+P+P9PlL29Md4azMVdSKxonVuRkB8xYSX5nsShQ5d/UdQRtEgmJZzaFLP88GjJynkCv/Y7tZFi
zC80rPoLwjEMqHwR2UpuE7xyontGbXIu1DKFmkxxALAOhuhdNy65P6RpgquglCNxNQaPJz7m9HTY
e5yWoIHE1hbiIPVBsx+QFqyZvI2PFa/RmFnQ3tqKjRduOwEqDJEpFj9b6Rb5GccVotBn5XeJ88cp
Hjys1uE2zNdodLeNzT75r1qo15lxlMylS4U9LIqOQLYNrcjqBYafFgT+Hzkc8OOmQobeTx6e4x68
jbT4XhBhgjb4mknagpcfZihlTWNTk7HDAdmQgXzg8ec9EGyPAV/DqeJ8xKjLxWwrfCocaE/S0XTb
662UAZJVF8EmiUr6l3o8wXxncVMMxl1UHxjtQ6iCR7skbhvSa+WAfjW39URQPL2M3g7ogJ/fAUAV
NiM2Ar1iIZ9395rHn2MzQetuQ6i0yqzgIQiErwhasNDZtFAEEenxzpxsDv0JvUJk5DU97QNAvNiY
zx/b19nYvjyWq+b6ksprRfihBE5msqdDcdVF077K312A5cUxt0WbK3R+gDuGj5vrp9RdLZFpnW5V
uSaDr1RFeHIVoE1fWyTzTzmGZ790Vvfy4VlbIuA9N5cY3sXSPXO+S0+wodx5IpxaMYFXssROBoyR
3ePPLhuz9f6NJQPMX0pW0xEckEprfcMPZNyID1vXlXxWaYsFlAZhoQGo55D834qFTxKC9TyMFb0Q
m0lO5Xmd6od/aoKCBzz1Za+Jngh9FOjgmxx0EEeuwhr/UV/duZb9BUZc32etkHcUJ8lMiYHj6TdI
oz6y9cdF7qduBPbUWUbpEWZzLTROzgQpsNLEfD1fPiu+QyiZ+7E6pM80ofW8pXhKpAmX1kt+SbZl
TQXQ5v4RK3LMfBvI5s7OgS5lPK7lrtYz6UDulwmeYha/EHIrJwYiCT8at/+3EUBrmSYAOz3G/Q+o
aydiEmnHLa1NXFw0X/EgT+m74MGWtzfW3Q3ZqJZLRGPcW+ru8MlLaconGpbUsqvl7+ezMy1pgFKT
ttXyFSYP/e/Iw2tBrbGrgi6dlvBZvCpr62ULhRcD/E66MOc5OoiSNJuthO7X/MahSdFkztB/YJ7/
zcKvfP3ggh3TpJSF0JLIuHBEm0AzjlwQ9tb8hxNOVo/90Lymz099JiEZZ9CEho1TOt+876NQij9A
mWH+3bs7fNeKgGwfaWxalRedx58xf7RsrOiF2SJkEOPhrRqYV5hGTvz3K6RyKMsloaiUEPEBDckt
tbG6cUuOQjVyIJjK9GQffB3uqftQMOrunjb4RfQevC0Vn1LE+fyUq2pcMhk7cOJI9ORTEX6Shqre
Df190T6KPv6g7PD4qY5RDL0IT2J8Y7ReK1zLbAITOtP5j9mNvmXZy7piNunhaO4HTiemxUpL9/Q0
oB9fRqBi96QeKdk3A2BFkngxMjkXQUuyupbK2vipq4VczhVvpJIv2qzh9mlrw/067drNaVtQKone
jEmTiKBoaH9LI8iRBpz1zQ1PAuocR8gWvXoZvAPSsS/EsK37oQ69DuLFBvG4NkAOJzCEr9uc6pKI
mRKo6fq+viWSaxZcVh/3k+iHMGjdyvC9zyyRmj5w//qFTXEg25y266t4dYyWIfBCmRvP51WVDf7i
iWsPKEcx5AWe1kLwOYVSKuHrT0S7x2qaDSJOHMMgtQl94mN2zUmYZaVQQM5MQjXMGITKNUVInsOw
P91I1SaZzivtu+wKopDKORUtcTiKPWhaPI0t9VQ27i7cmqGqwVK2NFyciUIkhdL2QFIzNCQ6WdCi
8hE+9r4Hnex1ywLZhHFOxKJ5hl8ruAlZUjqFrvGiZtEAudeizoFtfE+oT0IK7BNx69JHQ7ip6/SR
CIK8geuuRfCbwaIStT8m0bB+MYcRMNi8d23xmTJ+ZX+kc6VnQOQkt4VMNDtfN7KPGT7dDugpqMla
mGngx4L4cv/jB9CnL3uaZiYFGSROWKej9O4CZewFkmW7XXf5yoziS5vyu1WKkwZuEE1zR55LBe+3
Wfr8peI4ckOU9ZuhIeujkP7gcTlhkfGFA6tKZ+2VNyiJeXZxNeoH3TJEg+FYRtrEZ9Njt9PQ/+a6
4VYvf6ZU/IAscDMUm9Tq8HJ2X49fu91KTzVzsGm0Mg0DtA24YEJIScykVo05B9ox80FSEuXQevhR
aji4HGZpKspRyggJADqNuf/5VMrAbEvGHFn9AJohgXKXECNt0NelLsqo3aMmVss8nkBFrjaWd4ql
pS8bDRDLDaoUsVKMg6K3JfEhrRYC5S2aEDE24pBx1BweRWn3lsBsJtFik5/RrhJIhaqYxHsrAyuz
q4GtHnwLfe5LlaKqq6/Ykw7AJr8JaBFMYgB6D1cPVWubQ0Nfec9TKW5pGjZVH8kG9tctEzAzHZnM
ZZxgu0TPwkQdp5EKVvJ24IV341PfyDXwEF+DU3za5RYNX6VB1Y6Wr3nujXk3BOfcsCp3/pkFHtWg
1X891AVkpPJawUG9ZIggbis98bw9OsYllRNDYQM5RjtRFAgZVBfxTMA2dh3eHsnlKzSqwFT8Iaci
snET6ocTm2KObtmKNbazGcyvurnXo3+A6OasQPqHSAvDA3upQrkCvCXUYVNkokWRfENHpQZwzOfD
An3V5Ht39L1GyrmuFoupDIIXh81avHVFqyYY7rZfuxN/elQZK7+tNNiZaIJby2vey2zOCEZsAgX4
DFFHAioJ6vE7qltCgV2AYrQNiyx8lU77pxlAk7BwShCc26DQ2szstD8RSWunIUzDjYpf05qi6myy
azt8tcn6YZEpsBApU9w83t39lxzP5uLQqn8vv0P8u6KHD/SHMnGTO9bGxHows1I1kjiH8yd6xdK3
LQfj6r4YIyrlVKwg5m3KLpWFhUYy4CKE8uWajycKWlxNu4V8Ysxu87GVR+faQWBpiGDGyKyAuAgF
GcI0gbz9csN9g2aYaAscQLh2WmYlxB82ZLxIZlWGk17SDTiyjikZdop6wJhjxQDR2ePZNBOrBZ2b
CwK1/X7OyolwJWqZcfNzMYAtzUYJ8nCbt+1NFF+9V6/2QgFR3dhwQlIOlNh4WaVtTbb5mMIRGSUd
dxjFdWOw/ZtI367r0IuIrqE7MJun9CEBfrsptdkhhhD1B3rehFi1yIp/n2ELlpqMJ5lHRLyUnPqh
ARv6o3mhWILRjJ/9VbbCu8Ly9Q9EY7NnMKyxxXiA8KwMpqOOJmbNimFHbPcJiOrfAy5NU+nqr1Se
o0fgjC1/Kq+1nomvuLf9YxMZPz9qeKZ2tNZNycxeynN5ojT9LUV73ZUMQfidqI8Vj0cpiwC1Ij5t
BlkZb3w3hBz1sFgaxgO0eN/Bj/zgInUN4kF1fhOJo378RQxRb/t65W5tQ8vI9DCYR1uCnrMRJK7N
DNVeZ13O8vrNRwe2AnBmc6F4rtmeyroitwCICkNVFwbo5A04FZ2BLlw3I9oxVKA+0Vt3Mc5lBKel
CSgxL3NvBX6SKcCasGOZN3G1apwBMf9Um5cRfgRPR+e7Tawbw2HK37GAOgSZSFL+PuFZaP2N6PwT
Dsms41gJgXFoiGOKsBdhlqmxUnHm450JpLheO5CQVJqcuJ3noAHc72AavfolmKEKo2mV7kz/f/Hi
xJ/KKHf53rhdGTwz5Qn+q9dDvOpkkL8JPMr5BPIx3heHqALALAqgXmSXry7Ngykjo8hsWIZ26zSt
5TPivLccbK9Dlc4MgGSmZx+0fx+c3/hUUjMyePD6xc9uwOzPTC8ei6EqhZhoFwbFr27uaWN0Mv5T
YMtIJ03ndWym+PnCM71UdSv+hpFmtPvG1rsUtwdcJBNDdQU18OW9pO7KbhbReWrzj96qQ3sQM25i
DwIkcnirGbZjIo5WJHuzxAA2I6kTvuWKjtuVnfyEvJFB7RKgshfaLcxmWG8dW4SQkOChaFRNJjDq
lik0K6knxXbPLdpsmp96Enjtu8kpDwPeoD1CzyESp7UOKBMzxON+7426XYoiOvhYLHgWOZ9/4wiT
TskEF2i593JRN99uhvUlBL0WiDJ06ZLwjHZ7VUjVdJSSP7KaDH7wkidjAjcHmChSE8v/siMTKRDw
h3MFG7iI6jbUevz3LL6KH99Vt92Ox/DKiZpGZU7sQC/NfYgQj15NXLyHwFZarrIsdQ+AfAaN5rQi
S0gp0LKjUXincFsXJ/SFiPWvkic9poD++f6vm2j9iBYAGDbO91mDf3CRAtOBQn2/r09kzbmP9OfM
M3EN62wG00ZsS7d4H4pN5wGT8Jlron2PEIGNcSHiLZQbt9z2WPXdviGTrdhdW5em56Fkcy4KPI6f
elD/mYsUsII+96DQVsdg7ADf+snb3wZkMEDFuAhRxRceRLzxs3DiMFM7arM5nVyjzAr41POlxF1N
jyewGPdLsgOQsQdJguVApKFmHoCI4XgovaxzF+AjqSNaNeclr1fWBBE0lEDxvu3s0CDbJy4P27eP
TlpXbfyaDMlGW8oKPJMd8jCPeLf4wNnJ7tsKhL6gMPc0al6/wAdb/RQ8J17GhrGWvYX5L+eW6N0R
x+WXA2dQORzxvxftWm88olIqRpB0AaYmFSggy4kZ2U10bV/7J5vQ/6OYJV+3XUhocqQ9FlaZPcua
1H+C8fZR2YEVM1hErsW2oGlUQey4OZ9KrhAbBFHZUPQU6535MqEjuJEdLyoYP8Rxapt1by0Yu+Qf
iY/qlyzHjqCuge3JxX5kaGBM/GswIiIit6hRmIIe0X0KkN2BjObIaEn8DEKPaVZgMrlJBa2tD8EG
ZrBNHUnJcxb7/7htykN7YdpOqTyKv3ENN/xD1eoEd5uOa2yw63XHxRFQRikLrCGdguSrAz0KSx/l
tw8ySD5Df5UtBV7NaQWOIocxSEEqB5VaJSchVtkdk0h8wWtEuxJl3Nz27xvJ+Wwpm3QAtgOkiuao
CohM6SsZ6tun6C8f8EUwwbWu5P8lmrHoDzuA4xAztrAgQdmrOI2Ngzcb6F8dSwBAB6WuPCDm9qGQ
RKml7eV8cze2PQGFn/WvRKPqsfXTQxG75dznl9+Z5BS0jkW1Q/pZR0clCKuWCu434wAd5a+4b+3r
goluNkcyqmNl3eVFq65eeTlGJdBFT9BGR+jnixtLU243hVRtPO0CgF96iB6sargNRfnXWmgGhOhV
2F5BlT3S40mY48yqJk6HP0jYj2SLI61XmDU7KdfESPWcZBAwbQJNMJrrX8L2sBbJLzS5qUHCi1t6
fRzXa1/Qe5qcPQqx+g31lBuZ6u3PirIU31Q63SWBj/JwSonGVnWxy9ro50TXbYU5NdJsLLcCp5Be
vazcnud+1pbpDLsymDBo8dN4bBNNB3mA1+FIvB2D7TrfzrJK/8EJQkWdjdFOLQIaJXdlNO5drQYZ
CHVd2EH5a6L16XWNuNgkTXzfqgCGyaRzJ7SfcVOqw12NO+XGEJG9ArHeaJW64R/CndWjugNkr4ko
fIFXcZDoLwtDTgd3wSrLjvX93eCqXC0d+zyi9BUUiWtXuaCZHJ3NCGdhE8XKy1XyXNvt6YAoaHLl
Ck97NMR8Nq9haljSkaYPbtMCygPT16RT4jrFwLq341HScSRocAypeRJ+6sgJ3YZ18fz/WlxNB6n1
D9yO9jGW8MxY1WtQKEav4n9SgmwNsXG7hjK7G3Yx3kSwwvF3Nm/o1L5/TiV6iP3J6Lh1lj3BTWjs
KxhLEq1dLyzVcvXgOyMIQDoWjS/unAsEnCeBA8uigFpdD08O83jJjVsM3QbvzrrGTzu6TR3fwWFO
F2AWRdgaNd0fAMKSte8+gCcUomH+p7U5Eb8r5cdqppddDYiy/CTx05BKuHE1kI8JzaGcdjPxoKsG
R9M0clnIFaCxrxejoFl5N6sERVI0jzTDMbO1QWrwAyfbPCCrSaYbFi3JreSAgU7Md3F2sjYEI+cU
0EFQJxRDFQhjdqThvNp93YndI74wkCDIf9ZWdsMmWYnUtBxb/V/CkAi4UOnnsYCjJ5JVmQvoeXyy
Mv3+USG2r9nJZhwz3mC3NVu5JrytLcumFsDNDWTap/7UxheanPUjlZ1FfLKCmZB2JSeMndW8ZSGv
/zWJ8notrTIgrmIjwEs4xA2EK0LDxG94W50nzM76fJasxsFnBJtQm2wcSnYqOQvn5xNATm1rYf/0
ISaZxFwZ+X+8aUDt9EoIgGyAqJOm8f4SRWaGL7SeN01ovjEqWLsmzTVj6GxMll+98ui7aWQnDCJC
LV7HvK5hPUZjJWKkHuvJxEFOLiEOoVjDgjZkGCqO8R2qWviRGIxHV0WfpwPAeCaHbxAFE8d9wPlU
qWGSWM80uXkeQb1RHdMagLuOeabD9xG2e8LVap8pEW1LrdcBvWKEQPjX/tGslHZb6DEtohVIgsuN
oxSvO48GPNeEJuWp8cfnbINtrulYQRL3NzXHg+eOO6dEyYnZLlH7d1V/fO/OudZkUGSPt0UJ80h2
nTXTBwfF/F9HqKDbbRAMcbtmveNolNJMQ6JR6Zellx4mm5nxMuVgHXTD4c3k/Bu/UM30lu9/SZck
6Y1qhbWE0CAzNBl/qaCh2SQBZLyEOleaMQfIjKi0+3FBsjRgA4dEk1MDFnOkyoVCX/IEDP38zMqj
HzEqYlawHS+yMPWuHOWlUioWtnOsyWOZGxXi8KZaioF309bNCRmMBaQQlsQZS+Qakdrmm4Ay5Ul5
m1Im3R+fP6XbF5lZo+nF1CQ4/RQD0udPS/1r4JSoVBxzpQyQHATSDWQ41Uc+nOggjY0/PFtVYhVB
LoQJGLwm2JiYVteqZPVJxMyKWJpjbdmn9yk3yp+YeDpNbEStKgyN8Wg6eLzuqsSKqTOgk8J/qisM
b62RlpyvsiQdFKhlGspeIEDtXIB2DjFPlp5qC/BGOZJR5v1F7/CjxPH23xWqquwPNvLULpV8aB9y
kM8cGnotnTft8ZqU1z/TNKO1UZIXxU2QBnsgZJDXN3Ehmwm2RZRgycp5XoN3/Xtwus5QnYQwmuCX
C+d4EjpfzCnVydPAIOYKfIoDbQXHYQr1ML5uMqf9Mn09aDCuBs+bcpUJp4hWM6EKOJbdiBDFmfLd
jbMgYKVoChd8AqY5GqRzMSTxqq7IzrVWzMt/Fhl5yO9KlFjwOIuKIf9mJJKof46U4e2WGWIQI1jY
NldYuUd7yLpQUYgXNBviprLqdtM67+EVHXbw+P8O2cgb2fR3oT7C//Sg3Yres3LlKGdmY9pvg5gA
nrVddYRhOMFXRX9lQapXYMnripXvyUlWQLzN1BtRDpxoKYd6mxCl8wOd3EpxkkGXRoEvm/wXYpSz
5DKmd6n9UnZsfvFEOrkol8rrzVtUsC+PNPoxDRpuc6qe2QCnyJTOwHeDZLMw7HHj8Z/wTKq1TdpK
xBG73vgdR5XdsCXkPH18P9n1vMCoWNteWguyuC6s3SvN5YZkIfPOjyTadeRptB3vKRZFNHqoKnJH
M6DYDz41M9V8gV06OUF4FYB0kft5YVbdj2nQf1ur0lwjQnWAcnL/Z/pZ40ZspiLfJqlJSgeDeBAz
792KhfPIfrXQgN61YMyDbgR0N/9FztnTiu4c3FHfp3SFQQ3i10DFSBeGD+s0qab+Q4rMSP8dBHsm
r3pdSwlKNn+P+apemkhjn+Ik9zgbHGM0aUC2oQ+cgIym0kxJSFh2lgGYuQvdoiFm/4BW0stuvKkD
I3wgr0mHQk13EpppQO53Wn5bcfDFBu/a3XM1zyOc4oCLmxzbKiNrXc+a4EbcvBWNM14t2hXk7U8w
YiMb7tWY4HzMUYs+7p1CwAcrq5elocroIULjzOiqmRQnUo7yLW8Hzs07tCDyJz/EuKMj2NiAKad/
nB7yqzk13iteDuqT3kmsb4QFuVckzttkJuFxGFsgq1SumYe6ZzmCTzn2qWbd2KWfSYscFMSzbF3Y
AM27Gz4DKFttn8ql/6ySpBwa8UkjkzCggKERf9HlVjMHLUE7KJGa+5v7Ppo4evM+iflHX9RMYYdy
fXAUn5QTt+9dLf5Fh0BQkswdBzcpL4/1aAI9ygS2ZBjOWumDw2gmLohLvfSUr9aWRHZnCfJFPFjR
o9FzjMn2zWikyETDTDBFQp8rw5kWHqspykVVN8tdrnKw9fEqoFL05rg6bBCep859p6CgT7omyUTi
u3PEK9z1YAUzdEH7Pb6Ac8Ctkk709HtH2T38kHaQQsHfzEsQox6XVfFrrJyAWSuJzQ6uIsRwyrcj
FdJ6mGpYeqH1XAUJ4LXQBzJ11+HUdosfmdyAD64J8ATIAZfAbHfxt/FSxVK0+JHiBPMBSvB3YzsI
8AjScFhugCL28QNQGqvsBTbQO/cGXQFwn5tP3EhS1TuP1J4UlawOEd6qBFPKER1ECHZpUAsPia/+
CcN8UX71/k9fvh7fO4NsPzuFVTs2Oi3HiUvxam+FxunN2mabUI01qFVhieEC5qtuypioU1LjtlgK
cbh9LXdpeAdKuAMhZz+cIlDeDiZ24uH2RnJbh16schtqPXU01rXix92dyKOXWaHTo9qIjD9y9n8K
/V7Ud8xGWyIzBUexo4RWyv2iNOXSusNiMq964dfOBOlWtbWPeK9fpTt4pguEfvA0Oxp1xA2ygUF3
jhmZiTyHlxudc6lEdf+6f6eWD+1ee1aXSIBbzykGFOH/fNgcZQ/dFbHwaTNam3vIYJmmTeoCnFsr
SQSTPxrGGCYmmkeSuTCLxaAFC3M7ccc8B6vr5598pztYdrD0AGAS1yDbzSpBqouZj7Inv+6YnOnP
bYwjAJNuJ26NI0GkH8dRSSx3y+1iGyUheYXaOOu26Msi10WbnJ3JeNCLdu3TIkDiXk5FGySXcs0M
omzDiZzBeOeKnvAwkFfzIFEXk7ZSNAnVHe53KPm+kB7aTLZkuUXlDpIWPQvXy2wn5YC3R2jCbX3T
+kzSGJ4Ph/5OEr7EIwuuNvhpRue/8FuZdRFd/JrsCTGlSULY5/aElseQX77y8gHcwItLnjLfDwaU
ISb8CcbyYRGtO2Qqo0Rs0/M5Mbg6UvEzlGgy18sUpEE4+sbC/ecAjTGEgvOvvbtBNJ5SZHD6cQtl
X5mFnuzAKmcCP/6SrBERzDNXSCsa570fUnIyVFkSgrnLek25+HhdeNDHnWXG84PuzXZEA5fW0GZe
eHeBBGKD01ZWEOKVrYT1tIAENHw61MSFUWD061pvlLcv6+2DEh+C59AHZh3hF0+3MRGUlE546gRQ
oSgRkVLGO7x6G5JKp3y/bSfTaDWesAKhkRweUBUU0aA2gaBAhCv6qCPJV3/f3SalDQ+epA9J8J5J
xCN9t5XuMSFzd9cRtVpuc+IbMWKBm/LE2tFKfhIOp2jOs8iyOMFTUc+k6p9u6HTZHk8Tqo4QFLHr
SR+M2gARa2a50G/EMoyE1tHGHLN1ioUMMcKraFfKvON++C4XHbwbpdmO819eWV+9AXoudn01oWWP
52qmsJHMUKfdrsTEt+No6OZ7UCcUldk+xXtw0jNcPMEZaykgcAYK/4p5c7plEphjudHLYKNfG5sd
cRWHyfFumrWKAsXAgOeNUPkuuCp65PmMwviQsMEy31vr7khdzSm6WR9tfaetAuT0N/JimvNxus5e
3DTnGXVXz5Gv50NEyvdGowqRSjh4d91dEbwseLE1G2QgLD+/2+xctQGiN2/VcfHAqazOeqBOhdah
Up0MRx0e+Yy2/R+WNYDyAODm/WkVeWu/lwSqTzX/MNg70/tKO/7I5t7b7LTJsYSQ+Wd1IpPvYNo9
Y0fdUA2pXDONSwxIIekEjPETvMKXC5K8A7Tb6iAenn2EsLe0JNyxwqecfIqFJz1WkrTPk7C3cd94
k2FXjBq+7QdWzL5iq8rpA2gKXwOFbQDTBpbdQiqo4br8MumbVflZ69u05CSEzPO4qSW5BQymQGrE
/ykHiUaGszu/BwmniwoEP0dd6ZgN9q9Q4MqPOLVMtVcGFM7xuOUMwGPrXJK0MsG8wqsvyic8sRUW
mfJ3PxLQbyNNFkxy11bBKlNzQGPxDYXwbRu6Nw5WzR5AlxY4/haJp88q5XhfRRmCfUEREEyeQpjE
gemIjQmxKoj/9pIE6v//ar88Th8c7QT0V24kNQp+9M/V7hyWnpIvAHtb72LpZ/vCE9xvNAiMGZrL
0/fHFWG3sWc/PkbGeHelXMK871edcIlgaxj/ReUwVym2jeZGUZecq4vGvtuG/jU5a2KGTwBgF6Xp
77nHkqXT04h9XUVxAUzUtgB01fykhi/bKfx/wL4RRQBQxt3Qj/4xqNIp71FEK6DlUquIuF6PbL/U
ttKVyZSd9q0aovpjKeMshyLs1DVDx4/TfbWiEpkvZLqIlkUGLk+cmP8aLCEVO7SwfFLQV358ekWw
bJoBjlszS7MTgRTVzl6Jb5KlOofW88yMKMfSTBeQyylHQh5TgMvnmfB0o2EM7cBaMnlGKq/lkqWI
Cl0G/0xt6RjXTr2qRZXAj4EKcTqUlAp9btTfGMAW9gAcvWVfjm9ZXrHV/PKYWB5SE/Vvt+KG+7ou
tYbTg5y5tz02sc2IytT6PxJ2exxYYc3Q9Qqco7kqRan9+Rt892DVGfX+1V+29Bi7QYbBNUhFkPv9
aElKc1FYEcRcDQstokeJ2FBxurgT+Y67Y8ZgXoHsvi3d8AiXTizurCGX0GHsGihwLReBqdUJBdlJ
VOc3Av2t4CAJ4MpIvlaZ0x7t90QdscREZ8cZyCd6Unr5Zi65G0eGbpf+UZyFiNF1RWEctcj23JTK
8wLLqpypDGajS3zq18Wi5ehmE7IMC27zYUI5w90pRkKWF8bYmTgBxFMPXUW3ixnB/M2BGcNHKQ0p
j5GUTj3Ck3RtukLDZyWKwstWd8PLDUyafwSf5SIukjhLo4juRLdZZ6O8qiKRILcSqpHpL5uAxwSk
NbilbUpwKLpsZ1LrhVY+1wj5lsa+LJ+NGD0SsUj1YCWfTljsEqolJdf6Vy5NY3RRjl2S6xebmLdC
/DjCg4THS+P147FS5YvhKn8+5DaerL2A/iHKaoLZaZXlZXhOmjtBQRA7jCA0e/ReqJucJsdyeu8d
MGZ1gyVRq5Nz2js9Xuy9AZ9uLCHUzL4DD048XCiEx24KDF7VPcIZFWfZJB2Yo9U3x4sZmp4rH2lI
+4dNHqtY6GTqvy/75pYB70YsvNsgSPj8sDT0ZBTLNnFLPa63JKGeQJEskBmr4aakjTfQu5PC5/TU
wdE53HVl/kAZKlXhFfiJgPvo/gjrekJ5d/oJFFugUXJHhRZevbnQi4Nvzw4BGs7NisA7VIBjgUXX
bNmyUdIxCGkJN8rfHtKTR76t/K6wC3r4Ea1GHjI7PB4zvim2Vza0RK/DylagNSRVbwACIWc7jOl9
3qrghn+xw9Gt/h4JFNuKWlQudjb3yXnNPt4oFeTrnjmMxEWu4QiidrBwA0Abc99XnGDFtbj8lKm4
mYCjuuQQPRKP++UW4vpX0PwNlAeJWn6zcUHq4if2VPnJSxOs5lskM2spmGyID0DooVUAIWDHkPDT
KfX7dvdlgjbel/URS7pA6NxfqirYJsmfIOgOQBDLqsElBCtp/m213E/VOWSOgpkDFtKmauOUbOvI
bdQ+O5oYOCaPzM/035Z3pSsvdJl5Oou55mtzOUofvKjlh5XC0qO1vi7reeFqqZzFC+x5oxP61OV9
cst8NgGVLZq5NM6LpKsujcSs6R4PY8ReyuD5AFtccTgByFRsVK2gyVnT25HwXaN3ulr42ahC1x1l
vCEqPX2GVCQfUnc17Sv004k9sPFPGnYXpP0mlmINJbk6hsFAYAc3tEh2y8hkkXzMwJPCC7GMl6Z1
gCCjwbPlceQuzJU3xPS8T54do+mAOyFGvJ6nix6VwX5sNyVGhqU58i7ms9hytyu+PykQv5lnhtS+
nm9X9TsFcLkMOlxz0fDJRTeVM9XoXSJ61j6F9XmX5O1lUeJrgD7rpC6dR4I6gIj1U5FqgEW266fr
b7frIqLvzkNZ4PbzviLc6NYH4hub8Mg7kgY8z8PZqaRr2BiA1+ZgGnv3eoq878a0RpfmYoLUxQo5
SfMn/ITBwNqyFkEHo/Pbi4C1c8Cu9t2c8m0QPzIM7PKvY638zltd7lw2v60oQxhKmWkhUAVG9oCG
SayFr3IJHC4NZxfy3ODA1pHvIFTT2NhVvw9sblojJ63NgYcj15r5mfJYBdHdqsBXq2BF0cFutCU9
OQcnHa5VbkWTbtniFEjpwWbdC8RO4sQZ5BvRmWEFRxax0raWJsY+g+JgjsHwinznfkryfFy5Avv9
Kt24mQ1bQcMpb2slc/VwcZw3Vw6n/sIJiz0WimuK5T9Lcec34hU+yXGihHqpOT2N6OQzhnA6l56n
fkvDEW48662i7M6fESyyNu/2q7WniTuE/+JZk18caVqypf5dQOYa3LnS7/4Ar0q/ddmtgm93Te+D
JjQfYPuPbY0ssGRG72XtZzmI99ErYpxA0ZR1V0RIxTlazNnzEAJNrwVzpZYi8f4K2rH5UwYyCno9
0wDLIKeqp4NI/tfctt4IKGZ4kss0fga1ab5adby+Tp9UiDX0P1fgl5MHJWRbBDHg+Sf+gvFkU3Le
bakrUeqeSioKP1ocswu1fOgjxiNxw3i6cM9TdBbdLZN8lWy/C6Fu1G/ZOXLy1evt0A9py4Nc34HS
MC3qOnGtx3tRmmUrRoDm6UUOXmjpMqvcL6nxcslPHJ2p8AQ+jfger/MFkpl4ppoOYwUS2yJDqX6R
/1JpKJlRzTQkMH+05+ky+ML6s2h3zorxGM69/PvI4i2hbEoFm1Ul5ZOVL/1u0r3WoelidXzhSiFr
Mf6IdIAkwVYkRRlCMiXH8I2adT0Yo4sb0MMwqOKdftVOcJCpWizMVAKvQPiuSuzdSJmTSNXSAmnK
h4jNr1Jmtb4w0b7o5Y2sO8RQH5EieIQaDm7isolqQ7ahjk/Aq+ishtnW5pcgGsV7k2AxV2/+6qgD
oby0b7RjFrIdszm6tm5qOuVnCPJIrWs/Iuyj+CBGoM7EwLei4gkoiJdNSs+eyaA6ldScN8QA0w/9
vwEstMWkndT8X7aBw9/jSp6nbgkNkbEXEK5t615mFFJypfi1zAd81YiDXkeb/HLXBZfqOg3IyPSp
FMuVPbqv383FF2NzrP2P2wNn8mVvbt0jnHoj8RUzyuwL0Yd/3QIWzr43fYy3yQx2Sj+mo2n/DJ0e
w80Dk5p8JNtFZyi6yR/eDrttXi/1yOPg81vY7QgW8SEXqHcHc9FQ1VSj/fEliNZ28SZ13/27262Y
j2xS4RsKbyGm8NvhBbAH6IRpmuOliR490SnOjQV59IrYxAeeEcF6/XskrhpRis+PblSnQnr0NKjQ
titutbnSKCteqDjhSYkeT0lbOS0yvujSUiFTo3bjzYVg73hKzxIcClz8Pus/Gpmpy/obRKkjT50v
A24SnBfY0j3gcEY81Ih1mBXHOB3rrnSU+WH5IBMlqvlPWN8vMeLl9QSAywsaqW4p/ugBa0HciW/j
1IEabYzTeYRfAkJlALM8TqHiVwSkGnZRA4+wbEnGMTrfGXrqosbiVfddNcXeCAAyYlpvDpx4Hdin
etxgfmrMxBRYD4g0QBpUPyRLUKWCvcwseRjRTumtS1gUzjKGG///CMMCPu2Z0XlHLEfMCFymJDqz
GB0nMm0hB6WegVHiKrE9lbXcy8q/iF+Xx5yo/t/SDmyB4HUgsF9aWT4qrtUi0hTllFHjVmnH5j7e
BX80uU6+xpeElHCmBzSVX86irKiwLtBqMkQ9JC0fSoFyD+EwkQ9+KUVJgMMHkSPCfAcW+6qeRaqU
nD4LedSko/RxLPHkq6IeklAC6bd5E5eir4JoP7h3eLTU8dx5BEbVXXRGuqYC9BCL6TzXmnQcnHjb
cdhFh+rZcFZ07sMCAv5sO4bKcJK6IBDd16FHhtw7pyeY8L9DGJRa0Y1iGtw2WM93YewUbRDoB9Na
OvFe04MnRkUGmo6bYA1Na2Xl5yV6fKS26T2tlHvjp/SbDdeEejB3qOZQHEXTtggNz6YAkNpoCU8M
0DKVDmHSmv8GR+8iiA08s5y+VTOEg0uaPCMuzi6hMtuw+biloadqYKMIboXwBb7FVv3Q6Md2dkwE
PgHrGRKhR/L87YpLjiGCN4Av3r3TJ4w5CALDnsAizzm3TqjMdUzTk58lJ8Nw1AY4j9pes2vcFrGW
/lhCCuDR9xAu11KduM2ef/AsluPNRW99HoWmssDXM8s4Wi/LmHSPhRW5yx6jnl+agTeSmGA+euyi
vq0HGbYIkS58md3OLMDZoJHXWVi2Enr7+pBWhc7mVluqflGydoA4qZ9ZJA7PUYUrZkMlG0NlrauS
RM5oW73AownoYr66fQzC3+CvtCblon78UhABpLHepWuoQ+gyHO36fvRUDfW5r7I6sT8W/pyFV2Yp
YKqKFCXrJtNOXR3ghOsDJXvWE19SEaV2uUATFsPG1ZCVZ3VLE3u5FCUT713lE1asPy/WCCGIYtr8
lCbjUmnqQQz4wXQuBJPGUub1l3/pRoU+zCInx6lNahkev6u/ES5upyh65asZr1oKCZCVOmZpapc+
niDHclZpxazzvWjOxPCDnPdJw6zKEN/TXA77uUMtMhTDNCNV7NsTVvF99m2iZpv0u/W8bc0B3mHM
Ka02DhmfjxB5cg7Jz2P71AmhMR8qvEv/Bbi/HWcI5QFyeswBW0qR38k36lQIq7iVK+u/l41a8oZn
kh4AufjTXde71IMT/KxR+D2OYCg7cw6s0ubQ3u3K6d5YVAjQWy7luaayT0/TEvAyI8BKwZcab3lZ
zsXsCzgnlNBEb51CoAdz/ACCCF1JY+E6/OCkmxwcFvo+Lpl8DOc/CVmQkpDcD6OilVfGTQ0KsHZj
odXGFBmAWPxOfkEcQCTNy5/f/KvN8IFvLPs/2wJn/4uaTHbeGukcs2B+8cI2tmUqb991N0zfcitQ
3QSlcDHB5Sv1PA2DV1TNrTY+kxIMzD4xUpkzGLlsY8SROGLf7elW48nxi8v6e/59vWaaup+j2JMS
Kx5TENF9GpqxCWgZmr5VbI/9uv+o/pTitJx5LdfGH+6FShBJDUe30d6PJP4kzqD1W4nX7UESxP/n
FKXB+R/lwS2WiOpu+EKShIB7EQ2zDO1RkJ6ubkatSqsPk8OZQP8xvYU/GyiMl7VruNV1JUxjhYBq
jWPkFWVUc25TJ0NBMkRMKowX6PqVf9FYnII/7XcRSnJyoams1NNmNPU7faPLJqvO6s4EJMM9XF2i
iYYPBeb18R2vMQ+WdP4BsqE/vhArPMRDXh+e3swzBy0aiQ0Nf3r5y7SBrJorH/AvGBgs06By+ScW
lplekRVm4juXSfQwo7S9Zkf0a5Q0QNew/clMrHnQeGL6dft0L2pgoQwDXcH8SubThkObGEegihtk
9FnrSY5xjvWk5vYrmwlpdLAv+vTcvNsJVkgo1YtWZamOM3XNAkTWjVTBJvkScdN/XCr6do4SBA1b
cz4TkLGbe5iypYJJ7Sb8tW8u8+nO4aO2+Loj8hwylWFydPHIhpe6A64p2xRTZUfqE2Z164aMD9CC
29jMtQg4SxO+TVFrd6+TiXAlJDNBVIKAvRkC4SToO3lyP339sxRgg5RldEDR5kTAcflFuWPBqVC0
rvsRwOeiAEyfQNvpURdrevvzqFdFED5u4Ut7lKC0qN2zAN4QRPYZ8+JWPTgEJlQ3+LbICKzVGmRs
XI6BfaBqsgWqYkqOZwoGRjogRY+aZFxX3OVD27NMzAUB1Xq2+TA0Yq8thV5U/MRlZ2/dqs687NkK
aPCOxMWFBs7vU7XQDwL8Ppl+tNzQf010BzhOEqUj7Uu2bXo5A76nKJQzN5Sr2RhM3GfHbgxQxkDW
spmEVOv3dMUXYcEtbcmIBgYwr05a+k7ZaDIkAJqnW+nAv6iApCaKM21E1ZWUOX/QQIMwkFl1Ai/g
i501PzazsXWiYtKfPWff3VZo9kvan/V63O/8r1YLg/H4SNX449NAdMNEUBWQC47pejsRDi7oecry
ZhfXrOYYRaenqgZ7DMDeph+WoPbnH0BvqG+HBtOYXrpoBXyVvuQOAngY4W57YXYITlHqbdXsSEQ5
L0GMZ/61+JVAoXNOsVjl33nEbPYbesuOg+xgbgOUiHvXQulGkltXpqIDVlEc8zn9712bwPLIakBU
A2NCUkZ4shljUF4HVC6VReH3QMATLevbXPCStxsDZqwbTlKU5no2yQQiTUoLoqV7oI4z6zDAIeA9
dUK2F88q2T0C5GR8SbLP8a5Fs760x+FtJZNfWCJHtGwFrJ8nKQ3u/plxRDqrmsSzvVgNg79FP0tF
dLA74zvhmoFbGFIDJUjLEzXe97C+aSsuLwA9FNZKW8FvVr/BFrq3rwAL2vf4aMyFtGuzgY4rWe88
nrwOo/INRpYVnoODXyUB9cMzW1x6ROGE1oZcTRNa7sIAr3SnAdCdD6dsKzF0DBa1zt3NUh/lp3YD
z+K0Ux9E35YMo+Ac8X6dSt+9qQwohe1dn9ienybfIhtwGkOhLuvucT/mXlvADRSLoAOxcgQshVdX
MA5lHBEKxjp+8MCNOG4/PxJ2oIPuBfT1CSL/TYsfaGL0RW2Mh9/b7oygg95XvYMoWP797dCauve0
kmOtKhDfDRZRXvYWJeC6g+0MjPjoweJc9a/n/CzBfke8UBgxTGuo1GoElTZX9LKLvAHXXQYzQsIE
6ILaqfQL80gfz3ACuWutHGzEypSnHPX1DQ9q5XYMFWtun2pWRD0KvZ9cCksxM7a2jBBHzeXT5a0K
NYCPkn77Oqv4gulJNHMnhR1CyUf8d0g29e3K4NDpQYjyob+7D6KKRfz+4tnbEpjHj1EgSO8SsQrp
UC0z9qUdHk4NNzXQBTvBBJXNTxsP6cXRZfHDcH2dCBw3ZAyowxyEhBv7h13crLhvWdnHyc8gEmGS
sjbqxN2ZhzvLQl/TgGWv0OeFP1A0gfCQH7LTFa4dcKRwBwbbZXzcJ7nnFLM6FegrqfLCp79MtklI
jgjbFlyuMt5MKBnmSxVkPRjHSzXq0OcZzyGp6ZBuqectoQP68EEEXizOUBcG0oHw/Z2nRF0Creno
Cg5DKIEKB1XMEPGMbPLEimDj2t2Eb7NDhPi3QI6UoeMVbyrPbKCWZmJpcohsBlS9fBB7ZWcHhYQW
nCLcu9SpA11Qlfm9y8Jr8SMRNs1e8Qi6HDbHYbtxlZ1VNZgd+mJ0pkr/ztmBs5J0EE57rsYWBtFv
f8iNMowkcFOdiDTTBRplxsj0Uyi3tdUdoUelKMVMQyjLkxLptpPFHIIoUaVhtjxDc7l/J/W+Jj2D
EAikjgn+CZrdw5wXMlsynYVf34h52YkZsIiqbKfZm74aHsBKsd0Aio/+JlMvTbYhhQ4VaI9xP8cM
kIPGIyCB3/UbJePkRfMW0vmcmtiBFJ7q5t+PQEptFjDKaOtuO9m762J/NzjA8IzVLfprMcj0f6xZ
07Zrp70dQ8x0gZRCHlZTJrZg2+uNcf4zhzYJTue4rZGisLvx4O2fqHD46X5yr48lhXZ8DmtbYB5O
WGvg/fHnmqXB33Qfa8GJSMDsC4QpDoBb8zOndQEcMfVAaaxMl1e9o/4TuPrrPqH+EeS1u4T5eb6K
gsuSrEU3uA0e1lDSWM3LDxcEc87uoNxHt3Iu3IGtqJzsTZkhJk5zOu96BfQWCjTD0fwRbhyO8pbg
vmMxGBFlQ68fsMZgNpWpB6ms6iFrV+7xI/Ljw3fjKDE77kE9lCwhmoONsr5VqpSorVDn+XbjF/ya
ELYq/IbM919NkWzCKDlZEZqKIbczExhqzoxufb5v66vtLew5as3YFaWSt2fcfjg0SLDFWFWu6uL1
a2xKYncDKhI18O4SJyhn15pKzmsd9VotwCZf1PuyO8UmE3BiocFoVTuda12T41T/esu5EslWxjOq
6OmtH7jLyZUy5C3h3YZ2cgR71DtS7SzBxrvYFFKUFJynYKxHEE4pVVrDphedBI8ipgcjXIr0sDYM
z8fcJnLASI/czwM9y3azV2rM2PHuMj28Lv8ELV03oRHprqFjWP+q/wtHA8lo0Zw/m7NkX+8MgUwA
Ge3Fyou8Kfad+So5cA31O+ixZcvRnHDz5wiQrbwQQ059fuln62VkmXE9ew9/YfT0RD1YtHSiWr3k
VSrMQNSLCKG1czWMpr0Kvvsfqcpz02qt15PtKS9HxzzDzPoPJtb0UlS5RUFZ6n9G3xJLLCOdKbf4
tKx0DHl505ZdP20heCfjHLhPPqYuiiqnJfKUBJufCxmFf0Sc40EGMF7TvUIChXG4mFSOP8BbWh8S
goVdov4+nyGXE72WCSqH7wQ2wynJPC0Hrha2wXWmCmlAvt9Q2zwCy2phq7HFeLf2l9PBbycpPV9Y
poc9F4zCmlnnVLLmrcbXRWVZkf5AS9H9tNIiq12THLOj2nF0O7VtCBjlKjZWUKFgUEWnpwPAa85p
B1XMogVXBX4UnXsqBLFCuysVcdxwlJka10u8Hn1jy6pIy7hqm6jaL0YXRgwBg0idZuoLVI2KnKhW
Qr7vbfpSw/dJCCL+5RbS58mTtus5HQmArbOTyBmON0/oFsiNPxX306fXZTMWsgyjEZwnrQl7y+mB
UFHx3QbwBqQVfyT69MzbMb4VuiCqnVD0FvDFo+H3xQ7VAq88VhYsoXAyUJ7YJiUvPy2sIBrEjDQ2
aO/WqyrSLfwrio3wH545gAo55icxwqzC4dscHZ5gWLJYNc5A4GrZLLRVYYqX3yd46sfcvYQ3vvym
BNYm6AYm4bIyOkPNxzugFXHM2VDuSRD/Y1iFEXLdLl8NupEup34q3TgnEgt8pnFwYQwvMFsETa1L
Uxwod+7sUpY5NIUCkgkLLtqz6yu7mGgCOPN6yCu6Pme+C69fxB4sm9qRpo23gTk6qAFnzN6FOpkD
ocd6wSUmZ8Gmu2lvZJbFniIDtiThOIlBoJumTp1rFjSWSKftUbnAwxZAvjP2ikaRoAOPh0hkkZ68
LTffIHuKVh+QfzA/IXz3oq2m6dY+5KVnIMdZ0nmnsOWOsIsEBhZTnBvV4Bj+JbmPUO4Ja87Xma4Q
APATiVf0fUOIR0hQTe005oz2soYzcwlnan0bKBaGq35tFXnFExVciGup8Fb55SDsa8Trhb/tCTWX
/5pRP0WlCvDSHIx/5LcJzee3+QrDqNthZrIsB8PRDAoWrlmFZ01VYY5+m5uCFBvD6IMlu7PQJLR/
qk/G/hQwzbdDgbyqo+UbpnKSg6ITMwuyiiImGuQSdIsPbdOtzzn4w1vS78WTalLa+u+recNpbmcS
aUBnaG+4d2TGylG1dTFnqd7BzhEm6s1Ri8gjxpY3ViBhmGPG3MmqJPNs8JO8rxgeMZnHvx7TY/x5
BdkyguVONtiOHpxCQbesBHf5c82P/WmbA3hnExgS3+4RrvVgI6C3O5SVBA6PA2plm0y+fNF6zslK
dffStbUApb52NqADa3jNtllGDON+Iub1STTOna19u7mAoABPh84ru43+AdYEnGxYJqHGuLTEoX/+
SP3NgUsTvZoUcWVLiRkZYLD8LNTGUwfc0H8ihkh1yEsKo1iz9HcDMNrf5g877Ue3ng0S4+l34BXp
0hbNfW+SBTU1264oK3SwOOH0KwNyuCJXhPOZ3mA3LDdZFL5bvDgKQr3ackYF8Q1/6ll1fFvRY2FM
wN9sP0TeUIrBCMrdGqYsvUIPS48/3pByealqJXtil4B3z0Jwwd2pl/5StMKGFyfHq94fPDGCGfdp
kRRRTYbZaACyH0v8McO7yO4/ZbqSAiLTuUmr7Qg1MJUHnN050++uLPIWNduWpJvSzJ4LU/SqUXcP
LBLKigByV0o5cJOjrsgrCbK4F0K0Tx2uCSIfYunTsaKSem2e+ZQQltZN/dMbyKywYGighIybqdVo
ntsohcJqLAUw58AvcRZID3suP4nhoaEosiyatBLMk7lE6aEaFGSa/V5jeQRuPlw2fbfjkou8ZdET
NVCPhtK72PhazxUUSDIfpiBaJNp8SCZAtfpfYmVfws1v0qm33r1BudBjBQAjrQLrmFrW7h37+MX+
8p9k/B+TgRZcOnHlFx1wNgH4va41kATDy0rIlUJw7M7NpsL1Gg85fs9R4N2zNmuP5lPES8WBGKGN
jPa/UX5RB3eAjVrFzffCFTl3fsW3RK5CUG2yAIyDJPrt8erd7UYNTpXLadz29mURPVAI9yxqXPpD
2J6ltT/p9Ci1hEi1DR1ZWXdbo+cek702Gjx580IaQNa8S9q9a1mNuqVfGq6WU9gmfn54ZPEdWCdp
dSduEQ2qJTzQVPw07/N0/NFYXkE+mc+29byEA0XlbtXJe41O2eZK7BkUgIFWeQebv2PZFUNObM5y
U1ySQUlKtfs4VTX4+NFAcjku21K2NCBOntxfLsKjSnkcKD9tDvnajcCKU4dvSPHvYUNU7rpBZe5v
ji3yZakbJVPbW42VPIMmjmQBY9KNcSbhc4uuH+s2zK2C93aNVECj38q7QLRda4SxK6U6bNAMO11L
4eX39LszjdvXEVpDC38CwGxefAke2oiRj++2+lCOb++RvuRVAUsqoVvMpqHuUTi0umDpv0fDbjtf
GuLTv+NxDr3i56gAKkka3HTxzJllOiCynRcgH2il3I2Lej+qC2i2+QONpH91uOhnCBq5c8zFIRmp
pSutzW3rUyJ7QxfbIx5E7OY9sIAr8Kw837Ucy7yaInzhNLoHN1QrHBuWpqK+6ecxuXUffRZ6ZWmu
njcAcTi4GDsLrdxNzs/9aMBlE4MJGvi4oOdsVvj7pwQxlP8F59jb1/OwVjeej5LKuMLpG90ZzyiP
rtKrTJFczKvJrdm3sXcf1x1djKpAZEbaUOxlvaj4ZHUDXGEL78L5BCDkQS6zD00iq70BSLYz6QWc
2fhys/kBB6L7kdLeA6OByDc2tfr6YfPIJcy94fJa2sQVJ99dR/CmzoGibY11VBZ6mpezpZ/q7cpm
r8TwCrMWwGKxviMWpPYiDFIjC7/ueUa1r6ZMlpbqQ/uQ7lBdaOd3F/cSoy9GQhglh6wcCNUDfLup
V10D6vT9L/RQmKyqSqi28HOSoPVEC4d+BMoBXS0mJrk8td1Axs9V+3lCh+WiVOuxNMxl7ByMcnzY
JTm1WE4Huxa8H7OxLbyJWwTbUbG/XlO6U6DohArkXRRqW2xHh0jwLN9ovW+9q5nPaxdL0wjvpuE0
e/AqYCRx4QJTO8OgowOdphLQSTDyv81lf2TltfxDCrqMaBXNKvHlofDJVw0lS9thfI3rUZHyiNZe
uKUD5EHZ95D5HuEehfmcwXbpjnBtIQH8E4O5i4OEO8mi17EPLhzoHJVEQINzoZfEmgDhic36V+T8
cHWC19UUVBEzBYn5218+j0lgoZ0o/d3bUTXOS1pldtD+cE0sHUZz9MoMaJBTWiuvJ+5zog2uqqmH
GfprlY+PDxQESGIp79UYUBX5UBSEbcOULGyopqUEgT2ppSkQTIHWrhhs0KQe3NL0GVvOB70f+2hx
p3mnstJbi43zSb6iDLeb/b/E/i6b/WaRXNKdyIT/PVlZs+/sAaWpXHtu+NyVLwh2RklSrEwWphkW
k8OYR0EFyGZtqH0NZ0KWWlMKKtS77mxjEaiucQWSOxc2U0MjeUAZW9V5Tu5LS6Mm0khRG+WXcHGj
t+sU3uIIC/O8gaFWrbdOGNaBohTNLvxCVkC2CB/G/hAd2IqqyVKR4rBK6+SYf6EGjmLLWNHkU0Lo
yfejTSjBOmCVcQ4rb7Nc9FYYHJkVXDN7u+vC/ZJuLexgSETMad7yYAYfNU5asHDTR5RgYqyma1Sh
GVkzpLIoZwqYcLITwMa2SMwycbXl+jDy69ue6TNpUl4zSh9bkXpMfBrHWi1OleoN6PZ46kex6W+o
ikoigu2IO66zRjOnSZxL+InG2LfV7E5EP6M22HnpVTPD28U/dOxCiG2Y2kn66itC4Bn6NLK0tPy3
DbQGNpapNHfJhgu9CGopmfeOle+AcVKulFeA2vM9G/ziQjbwMZ2QS/LQHAPLffaajwolw/BMKHR5
KrOoovxgyAuzD9VgwsGeeN9GlYinrmM84vmgmbzfOVrumPhte+Q5B5AGfkWC5HjRKmRntCN+RzNz
1sc1YqsOUTqSZSKirHaHInbbrwqXQAxZFkJOPNZtpIPMhtsg8Wl6ptvwLfEFY2wbewPxBv9pPDpE
llNg6D0ERrFJnYvV5XtMyw8FC04NBcZhoAZGiQcYuH+xrJ8Ki9GJ/1A1+Bn1zzDNU8GsPBEfzsEE
kc1TBoGBG+ZJ32RluANaE4VDl9bnkUFj2etYA0WkXSJR0VzWTZnZUChNM+Ip+htlWO0n3GS3QvGv
S6OKiJsUBuCVpjw+cHuhW985bmvxdbJHBGB99qfYAPSdICTzoJQGHy7SfJIsIOePI4JTEVYrcmcG
B8F5rg4GQuTp6tBOEDgcgGnerkiEuAbMSiALlj0h3tDF+hd9aTZo22PnT7N9oY1v/g1Oh6ClJMAF
awIHlR831g+NlyTDABV6b4VsdmVcwAdvVmVmPzO/RqEFonqcsszaSqV6TxLHxVKbA96ToajjaDhB
5k40xvKwfILy0pF9zwYZf6T0TGS1CtTsO4D8fXfqxZZA+CsDte/z3mseCY+FgT96liHgYgleLr/r
kzZzea4ro2JnPAY2XUFS1mp27QQ87/Frd2ZpkLGnQf8cEvdS+vk8JLWEtRAqzh2AOyu8Sop36cso
9W2kEdSUcv20TVBSDZj/HTKoJAn+P6dayTzmpujFD6i2iERElgAwSKPJAsa78ZqdSCZshYP6JlBE
uaqMb3i3O8KC6kNyJBUNfuS3moysOvhWADnoRXZ4tnFu9uQP4aeOEPOLVNPrS/4W/OucYDNC9AEO
e2A6SlrUNGHBFmPc4tVPOWx+TDwsovTPow/gzsI3ii1kNgSsGxPGaJlH7vQubUvLFe5OPVWni9A+
eulPm2o99DSENJjoXBka776gf+vjUnH6vj9r4YKWdiRwoxsfWdWKGcdgSe6TMJ2KGk/DOz5oO7H2
Slp/hCnuQ5hg8oYXxTzTnPRTiIGqQlvRWSCHXj4r92RPMJwM9nNVjoMgxfMs7NzS027/9uuoBxAc
b4RtLFxQtSYp1hTiQA7H9ZPdmJkViKibFiX9jVKtcUjrDvp7xOMLuawKlZOBKqUXIV/hLUCPeIJM
1DXurXUOW/aJjfSthNy4tvX0XMdrHjyJTH32th34kq8GY6i4KujEHiRdteEQ4x3AJJWrXStd6Ng7
dBlSYwD8Y3mJSsGOSsEZ/YYdbvd1VauHh8kWj2lfCRf908d5WY4BO0iuNbbClkVxzsLn6dCyPlWe
joCEuzoGq1qb6NcpAUd5btL43DLULCojPXHGeyTddEHOPVK1VfKUoK/SsjpzUNqtx9IHmVS9Y9ti
XqvP/KgA0cs4UNrY9TR9uGcDz3oZRI0fWFolD8Dl08gvcRmNUbxVQztVrCr2ul+ucBQ/2basobQj
AVBlug2PkJvhgvlra4BSVBJ7H5sy1SfJ21OjRH+3V7ILkpRFeYTyM/y/lARi/Mpy1YPgvjkw6wvP
TvvpUKTGsNXsTddHDjA5y0Q/1zvZMNbbt+tXFtnwF0qzT+kUglml/oVR+SV5OiqPOLLrV4clXL1x
XGxiO2j8stoEnaJyEk+RLZTA6//HuPupAxf9hAuoyuv2mEcEdwa9igny+pJZKRcbeOJZT9y+ZGag
SaXsOE0rqGU3DF/ItJWt+1aGt+x1pfLMZtVdeR5+Djqe4xvTKrOhldslbtoSWPZhQ+m23FiCoJ/z
F4LT0ZC6N3NPinl0lo1tDVXrxkNRge06cpD2LsQr7M1hBgTtvkBqrZccX3HTXptxLtCpLcSxn+lE
NleohQXkx6mOAMdjh19K46iQG4/Ly8bTO9jzF35I9CfmBi9JocZbJX/E9DsYODvL3dOeo5LlxaD3
80FOkDwCxfqHftYJt5oHHgxAs8cDhuaBpdHkR4Ot9DlgiIPubIbjG1B3H+knw9XAUFTXGPstT9zc
4cV6Xl4Ma2UizBJpO9Zt/3g0By+cbjPklg6ZEfJMhn9wW6D5PH1w259Suoly+O+eYWW0tGvhEkH+
yuzOpIq6BDAUdb3kr4jTerxsY+FVe3r9fv/Y9tX5EfNdjpHBVrh/PsC/vm4RjIpuVovEA6P9TJCj
WR1zOGfn2Ba2dedEfeSdXsraW8mHw12ZRbTRdV5U1aDH7xiDZ/XIghgvom/UIR4hTEq7vLi2AjR1
Iw9s9cN2CJNAOjoO/4ADjnBk127klodfWoWW2+Mk4CJY+H8hZtPkiJYE4xP6gk/JziY1ZAF0FxUM
S7tqGuKdDAj2dNeehCdm8r0SFSPIaYYomP/QTVMMVJ2YPLUzuE2TFfwAtw+WovusurRnrWscGUlF
DhMJajFAGw8DXH8KT9QfWZc/HdXGlX5DsFiDDJesDqvksYQtrLtpJtlPA5F6tvYYHioFaMwlpEAN
WmIMa8Jo27Ft7W3vDemDHnB9yJCnFWfnvgV1N/s2FCXTZAz7Eo9AnLG4kJpUqlBF0kkh0xDbWTny
W4AfOAhxrVsCpE/JuFWGpRh9NJCv/+vW2cWt9IeQ+JFNjNZmGKJhzGdsUJeUBN3Soh3xYd35AU6x
L3pPISQL/rEWx9VHUQSFzb7S6zAIU/4T5Vr5KWqbjvhjXqbhG/2MMkdxNscpUgsMhwhxr7g9xdDq
+Xh43ibE6R8SI96aj24Mfl0Y6YS+HO5gjh0jGxkq+XR+W8HckCkG+Oy4+bvVchrlxXnl2mZA7S+L
f+QJuVCjUK32en2N4fXtpH1ZOD3DwsKkKw0iVxvgjOI0Z2F38OSFGoT3xpzuWC+HCbJ8J34zfaLs
0y6Ce6d2Wk/O/43J1qA87GVBjAJYpCxkUu1jHwdvXpv7wbz0X6hDByQxVyHU9tkl9QesdTs4TmX5
PjlSlm5Mb91/fV99D/h0Xb+y+6gBA2IPURXnlH/9ncsvV8uSmltgRSlf7aFiNY2Ob7/WeWl50KAe
T2cEOFOyCfAIWl0XrcWNZp/mJeeVOiF9lEOtk/E3toTfAfnAgh9C//uuA67BV12jnySyeNZj9Izq
cI9D8cpzFoWw1nnv+AOWLalVVO0+TAOA681q1QgZVGP93w1o2UznWczNam/70WMASW+pOyIH+YNa
BQ8kUwHlGJ8PPBiq5PPlhN3ExL77sfqOO194+FcfPiEYHbsjYO9Qha1DKLoOlBSVCMsQk1zL4R5u
ASxTRkFIKReqoI4+ORakMpzu99F2feeRkug7f5+Va5UI0uT72f94bGf/1kAwS5ur4JyqIcjLNXY3
dNGQxcWeYPENZ9CFb+aZg+aG6uhyUgtM1vmfzkyTPcOv4qUPjrdDxDjYhbleKSJKm1cmAuhyu2cR
qohE1T3EFDQIxItrzffpHnrP191yyaCrPub0s0ayDqXaraddEJ+Dj9T2yR48Ac5bUjIPCJAjQrSV
rZ8K+w7HeuEP6sc7a0cDF4j/TUwhlhSfRzL7ycebfgSuJU7tbgKB4OeiWoCWoKT6Vp0OL2LEvX5H
1LXn76F4EoMU+QJvo2p6nP93QZNlL8K8RjvCP2MpR7iTEXjMnDTIFWdj3TWJbUN9gkJ3qRFXWGb+
eYqa3f7wEaJ2e7+553/yQGY8NuY7fBkbTPxVkMYB6XypkAZYrisDUQcGvMZNNtoCwiHqRzJO6gfY
S3zXOu9S39WE8REI9Es5ZSF3l3QNgUZtLfsvX2KzicevsfAksD3v+Q1IIgEY7DrR9VnzJpyoJ6Qk
SLKjyVRChAGdKD9jwKzp9YcLRw3ghBtG2gF0MYS7qqN0ukDSkoy7QStpfwEM04kPXv26hlOCD8T1
8DolqPrYDdNGCz8GXtsyjC8NyKEhYd8gcpMUGbyu/LgyfbW304+r8LugKJIsN5iey4FE5IGJQLze
fOL5K4lV1MsjvbFKdG1PUhDn2438KOWENTkzhF6kViPi324UlviP827pW6zbl/hnQKb+wEbi+zL1
KA/WD1kqOmQlOWmBRCLXPY2Pe5xpaR1PDr6J3+EEnQpyBPaDpxCGJqdEz5c/CWc4oCN7WwZGo3Vb
lerb3BckhH9/VhkcipmqbJIpl03Zxt9fiPxTKhZaKhZDvU9Bi1+/d/r//mWsublVhnfX7eJaeGEk
G6TW2crtGjGOYJZZpNWWrTX7COQeIWvlj4dz0ATpKYIhrjvPUg5TBadCLc3j8FIupdV8z9SscfFO
LvhAHBCaBxP0Xvr8R9B5zON7rKOFNrlzsovknJcX7Jlg6mWyI1birRaqsTqWt77SsavAf8yLkYMJ
sK2lpScvnRu77A4bNn7FAIl1UgaU6P/peB3fAWmcD1cYEzROYs2/v6uE5Pp/P/T8eOO8vgaylrFl
bociuPMnqZrnfFeH8aXg6iNqhCeDdz1G0HoPmU1d5zmtm/deyKJPhaFIx6f7hfC67Q5sEW1ihZBO
Stimz5vt41CMxxBo2RzFT4kpJCzgrGrykeuTUs9cBJhnKX9Xp30g/hSA9WSPwyAJLD3gzudZuawW
TYvbsOpTk2pO5oxwKpyMWDm8Ss0r+ico7DBkmt6NzL3CQ73oMybPoR/snsXRHU0JGsVN4ljKjK8W
FOzNJcLpgWGVHzq/W6mqYl/9YDGXquWwkk9o+RxccjRB8YJgISlzuqjXH4wJwoZeKeUPJr9uXZC/
6latYnIiptL7+0zhrGhnkTS1b2WjrRuiCrg+X1xkntdJ/WGAz1/kiqh6OyGyUdkZUZZrZL/e88u2
SZN/lp/FsCeNpLgPc8WNFUI1a45Ir+iOHa6nCXoLjw2CB+Iy7R4/gCkeyJUayePFxaB4pKYkKoXe
T7ECA0BIId9Y6aORyTSs+wLQCsrWVV/u38EDXr0FfNgbsFf1Zu/egBDM5zFtczPEmFAPsZSLtvQo
ypYUwVVIRbBeq9dwXhRS1RS8odO2HgeqonXrP1aP8R4lR6kXVYBBknNXep7u0fQW//qsZyE7I0s2
KpWmHJTDTwXPJv8sGLauBG8wc4+bb6L55JVNUOGRFAr/zWCwX9+3v3Jg6rvLOnZP6yVKLDyeM/ci
eWCst3n0Y3pl1PeHVSlc+IhLNVYrSs8T+kaPs5P42IQqWco3Lrw92QWnigf9FiTKZjz2BoCPWtVt
j4aJ7gbNaIulUtQyMSMBL3RGwaoDcnGLMSjldxPpyVa5AwMkK8jqK5bNvrzYH4pZ6QeCjJYch2ly
qTMiRe7ZDLUnjCEuNAPsrZ15+jxlJrS40pqctaKroCBvbh5zIBpBNXgXNdnqO3cPjNxXaD32rlDx
XmH0CZS0raa2M9iRT8TYGKb1nVFrECqkwnSdSSoV8mTY+VQHPs0HaYRbE6H+oHozBqyiD827n6kg
DPxiXPa9zYG9y2a2Mk4k0Sa3Sj9Du3Bt9hSYTE220G29muSDI4KFk920CJA4y6wpNit/MpaJ0Xzi
qy6FGzTRnPzeLkoONPkL+4L5eETsbWGtoBBe1f7FSzdzFsHm+h0JT5PwCH066Tnkkf35n/WleH08
0NmSYXYXq1v133y51xaAsaocP4sl0nwOEOP41vJeQMwJjIxq38qdks8qNfPVmb1Bz4wB0LusVezG
7auIgg9yKLfEVPWcJWCQVbtUJ/oVFQdJpOpIznqbt0yPTrnEcbMCE4vwVEvXjh+Yi6sGe9475rMi
aXH1JCx9etldDbZtoYdUJeK/GtJhKqd1ZD65gOPxEgT0KZDjtLFIdGDyIxIDgq+ygSgRIW1Z5A2f
FYGd5dlpT/nGjUnoFSxt6b679u1SVpsmh1HdxL4j5QKDJ2l1CBAzzwx1p2j3O9vHG+h/MZCDmp9q
Sl1RTEFIge7y5/idfXco94U54aQb+urXOIrtzdtJRusPi2TKewv2ogKqWA1ud8dYtrEjgnOyffcV
43lbaUyCWvv5ijokVM91rQCFi6Ool/LV50E6PX3Yg9SFO3FbCpsTF5ohZPx4i+Th/Cqpjwt+WtsB
KnGVCd/TyHkwHsCcCvZRG1bdwG/46v0Q6H4ItC09ipsfEJ5SCWtgiDMdP1taBCv6PIwfXYrXMEJT
mkUXpnIPP7y1c6QlOz65zw3YmbeXc5wgzc3Js6adFm7WNrc0nSKzkcHyXodNkXmOms5oxYXT/ytd
eIKUh5dYAaGdqA+eSdpAobQbanOEDxoR51WNjR2uxZ4B0KVPvQGH63uicsklgBliNzCPb4auWoKI
/HeO9t7jVe2Yzlzngmrsrvm5CmPShxOmSJT8UUUhI2UvNGF5NaE4eW+dWXyoduNOaUnLbSw+Kbn3
66fEbeJZdy/u0VVgoIgvjwBQdGyogHpnIpFFeSoEI7qOzY966F5dRcc5LF4QaOkKSYYot0JIWM9/
5vx6liHnLlCkqXu7cmMaNhq+QzlUs3txHIOo5pmxavIwTeGAVQHhz6e4r22tOx2bqbWhGI2fZ7nx
mU0rI1VitP+NS+JsmU6ZOPmczY8dgmtXt7yVAI+62vuw+dmCrPoo4JGpDR4iRn6G91MILU3Orerh
LWvVw0VuqUofRsvhHA5hV0bBjjrg2zZNTVM5Avo7y5tadKrwWJhf5kdB483+2kYu5eBLARu7Ii6p
kJ77FJLXQY6zmihlpVFyb6aluK3seaBvwd7t+daT4I5ohnrKUPg9Mc6j1xcY+NTf0GajlZxwdIKc
Gy9t3wTe7k4hS09HXuRv/ybKMScumF8viablvJT0P6V3pyZtjPx42fKecIkUF1sMvMIvTCOBoU0c
1sAqa//+plLJFj0yPS9lsaJ3dhUilyQ1yqWrd+QcuJxrn6Lni+2GE3iJpkpy2aWji7yG0PO1BWiq
/DgPZ+jDjRro7ylj5KylzomGnd/LwC8QC7Yw7SMtpJpCJE1OSNSgFb5gnM5vBMDGhBnQFIMGRbD3
pR4fozebi2Wv5k0odZHTq8ueO2gNQDmOtdUoBUFLfVSS0MOaYTnwR0HyO9IQHBXTXUtZ4oNemshl
yd/SpgY5o1cOC5/CV9E7nS42kek7Y/WXdm5WeaCqZOW2n/wZZihHY7cfcj1sZcPodtrljV5x21Wr
wnyJ8ZGK4JneRl6OwwsUv6rhSK0Zn0LdhgHx6rj12aTGWmj7LvA50ZybIJdMyKcxl+UNjvTiQem1
wIOL4Gm9bo23MarIJtC72oMauBLlzfuJZ9pOVR6U7T0wJ182K/11Kv++KnglSSXZ67UdJ7OND5lB
v/YNJa5sWpgZOThW2yCDyvMmTZtwwzyHPNuuBil45ELUGzKN/vVs+Qpt2KY2pQH0cM3CG+CgrFvA
H1wU3746gEdYamwzsOFXOeVAtAkb8VLntmokaLd8waX2KZUvYeaMsUsbIOWiG+czWaLU/3gV0Kvh
WQnbfczNncZunvOX6njzQaj1Qw1pReDL6GHYUdRsq0RS6QxlPWlcDTMDUTbLSHwfX+L8QEyF1T2s
5+biWkkiBUCEfhMYpxXCCj/xiLmTFJwUWXXPVUE4u9ywYzAJxAshPzKWCMS/iN8g75Tp4/zgndNC
IHSsNBIUya8Vc4HZUWEdw9juJhjvfBflWytohWUx0vpv0rX0UmFDDpJf3xPN0LFaNtMwG15V75fz
wMVAXgGvATOp/7fgQOk+3sYH1AgqDLdT2zyvZRwA7zUXBgyJAFeKqN8DhVUX1ZMxMH4PugQ/MR8Q
cyoKNi86GxnhAnjL2Md30DoeYDbsjrfznP5I/FauP/gEfpW3CVB78IknCCBuI78ToVYpuTpam1f6
IHckbhWuzwWbZXhXmdSY5+SKXqOvfwD/ad5yU7KA3ZrKRSlWRD8QDBgzDngcKJ+C6z+WW0YIDsF9
o1FBvkaaIHkXHWqxE2H7nEmrCPN+rsP0yKVGvW/BgblERklbkw911l+Wnkc4uERfxdsSyDSUAPXB
0ZNoda2ycx5QCe1LrlT4ChjpEVCJAOmJTwlJLQZZk7a3Xzcc9WyGm+Jbr3qAVJyfVgOHwFFweQWq
vyEm2mLBuhbt3P6hi8itWKpZamxWnysNB4+7fZvwB4R09CxOoK8Pi9MeCS0YiIeitmcVGBfRcj3s
WAQmwUWWSZBtgkoUwQc879VV2WanE6e1J+WN7x2GeOlNaBYxi/PpXXC63ZYXGih4HJDTYbFR4GBs
4oAi/sn35+CUlHitU74RcJOl9J/Ip9qQgELV5Lfv6twCxLnrO9twyzosRHCHv3NwEHcgi03AuPLu
6TAU3UgjMfEdP+OFjYe9RxXp8qysGB9eUbbiHJgatkThCUnZrV+sgsIq6kOuVskWSHEwgR0TzQHL
W/M50RudyTFa59payRea+5lx2Vran1xIS5akwWHufBi3QjLcktTltF5Kq/do7m+Eo7H8Piy4gFWh
aDQus0yIvlgCDhT692UQ4pteWImOaIStjMIeTNl8e2dHvs9QwvMASxzGZgJwKeT5OVm5bCy5EO2p
ruvjwRYZ3z1tYeFPfkwxe861Cwgy5Na4N1bGYT/l6VJtMKfo5C2LNwEC0CpNcjuXh5hlzK/ZS1KT
rxnwnoj9ArJPE4pmelHhNCRhyM/q8hB1ht6VbiazcmEuSXrXRNxkiFhAlemowKK2dDsdN8QGGmbS
ulUbDNH6C/MjZagVSsiqrhL7vycMIIJdA3+WcTtxQ9mySpsjj6pO0SKNsw7Y7jN+yFH1r0xRGo4J
rLNRdjNVIYJsTD3VCgCY58JyMT/6/YlyI89TRY5Pis+uc7XLYSupd4bFw7POp8t9TvIzOgcGuWdc
IX8yuDhpq5rOkem31iBbkjs4kn/J45j5DZlaygldW7nP6TW/seClYk9PZcIS9KIw9Nyg2370zxYD
mhBTdqHXp95JfusVUftLeRsJklMkJPkTWyDYp5NuX4lHAGt6AS0O/XbLoX0c7UrYztlXoSQOnv3m
y16K9WmWiDDALXHtEo79soz2pZzxCyjkAPlurmc/pk2/g0TCgyEUKkbQj3MhjhwMzwGPp0vLvw3p
5PZgnXphHdtF+w/m3jbmdfOo58Gg4XAtvehegP2RCN0ojYcxEYqgCBKcyBq3DsvtAf2Dn5RBHoRd
i5/lpWuC80r8C7Cgiv3A5V4TyX/OOBC+XKo0GE0tv7w+ASaHdtnkUYRX7ATuGd3OQk5NRmnpaBSo
Eqa8DLjrlEnYCVPqqYZa53C/7nNR3LNikH1aD1JFo661Ddoqdp90JYDZryxRNvHj06it3iEqWyqO
q4EV37vhPA4LckoTqOx4K0fXETmMHfps24FqBYi14LAEkF4Jetm8ymMZ0/3+0e4ZUZUZ8zO6O+lJ
/E0zGJPPwFO+KiKi4op5cz1tGyhf2V/pZXAKnVr9sf4jDoP8H/jIdO89BrvjA0JDtalVSHG9ygo2
1Iy43m/yibGfvLGyD8qnNPSJPcYnPghZnmWkXsjxYMkOR18JC+SWuwHlhcZA1XBFVskZtGMZHeJw
3VAjXN2bf8CjD1PZQhwG2ohlx9vGZas1Fa/U78iqpv8x6ObuJ4jj1G1ZGitt9fR3rRtuhQ/caBdj
aqsJWJ2VqsyFU/zdQZnhtgPp0WRRsnNHCqd3l4i/WfBGIPpxbcO489ki+SYVsQzS/qcaYbyUJBgz
+XazkD5UaAO+CfJ6N5D+bbm0CFjJ9TuCDHtDrH39rZ8i6vBMmUGGmiv5jyFYyklzf1hjKHbBaIeD
g/5Oj99CIjcv/C+OcjzvEQXcocSWklDA8oHC3ur+J0IM2DJHX70h+aSwB+MzexqOHmFzq3guzXTD
gLpf1bEk8nSnZdbalTQAYxzLZ+Z3CkYBoDtMz35r0x02gbmay8AHWcjNKh4EbDDTwjUSFi7ozpTJ
S6IvMHATsErgT1zwnZuNTICv+9NP6g4YlqCfA/2hknF9Mxh3naaRkpbx+xUHAOQekCpZlx8uI2fG
P5A3EaCTDjRKcmSYssAcKxgLmrbvsQAgVTG/yGGpk69hAz7ybV24AmmMhC070oickEWcoJHNTzTI
rAtvCcf9/5gQfyyI2PQwdBQrjnVjaFgwwavo99yBPze46+SbLOj2a8uZaGIDOALWh4ztc0QxLsz2
mb79UCbkeTCy7owHkL7lT6OvyLmXqPDeOmmOe4tX8b+VMj2D1tDls4g70B2/UX6/JcfRMbsPHWBo
4Q4bvC7+kd6oUjd5g+o9t2v+Dlus3n/RwONpkeP4DkNYqdv/lmrqCo3P1EUmyW74QASonq6FeZ3L
t9205IwaGPX90KG0AJpnOt6/97nBgRFCkmKHIGtc3bypANUjEKfZ/Ma1Fu5pk/VSQGDyoPeUA5cv
b0mLGZjOYvrrMBXsWzk2MUXRqpL5sTlRoIZ6WdzV/vF17CtJ/AQJpxTTGsv+Y52YxDjMdrcR3JN+
1NxA7EIMZU9xMdtc+d31WBL8LjRNBayGJxtQ74eBWiuxizs7+CJKgOPmEsJPXTGK/5Fv61wwLXIS
FSKu6xiInnXtUnuf8t/FKhJ6nrQzlJzE9xQHZp7m6opyzpu1uK5JACxfSd7X8NtaJS93ygGyiXEB
YQ5sK/gqiy2xAfBPeYj5bk2AakGCFKaUwfmWihQRt8PpD+sVU0Cg5IeLc0bXg3mB/LIXeFyHaG3d
+s5yzg/fHROcC4bL+GfqjdUaeA5uxPbBytwnvywwKG00UcHYRPh5O52vBP0OvcknsiEtH7/1GnQW
6QjkGJErbwQm3NPRWV6ALKsgOy5mSBRK/ZyV+dNo1ClSpQUoTiocntweSeiG9ZltPTAkBA1uICaK
uRocx0d+UE6xzROmIovObZRPyWypWem2aHKWpqCnYp11DeKEj044qkxd28YRVRYu6MdxneV9fpcr
G1F2VHRH+QQNpLiNu0HacV53hrR4hF4groRwibNLwp5XQ2JJnBRDOLYBvvsZG5xwHCIdD9QszncD
FiirCn37mShlrXyGtJbPDAQKT/OVmh1czBvIYfGd2SyDwaP6Gry84ZEFi53Fw33n+0HZ7++WEwgJ
kRBRZHQ0sd3hUsTrnGC7XuexEMWcukacuTMf1zaVy5K7RdtWuI+Pw6G4Ecdi5nY227ceKPBNxlEv
HV02JjHNRCTKN1YWo78VW94VSR/R89DmLholFYhHoTBp6AoUdnzvZi3ovLpGRn0k7rHn+/8Lvg/V
wBkQ1GjX26l+FxUnRvEfE5BJIo33qUcXbIOeQoFhnuiLv4Fwd/LoSDdJ7d4vGwcLjT99HDfaLxKJ
uOMeQfJ+qFlF17CEvRFIErdb0DkoMuqPIdQKpxEteI35MJ6kVzQ4kp50eHl9ouuc6D6yOrZPiWxB
gUThERUvvijAkDG0JEhSC85XWWx0rysVZlzqqzWtIkKZ5sqbWJueV/lrUt8evFKYmUTxWW8/1wZW
mxpOhF/NbY6QxQvUXxN46OYzx8E/kpl2PNNJnUuGt4YIOeanefTEONW63ntSpgBNu88EkdkRhbpX
n/AO2hG7mtee9z5goWveGWE4pFJkgY8ft9bJGL6ztwU3Ycd6T77P87fFuoqtORIkRId1Keu9LJde
yfeTZkSlYCRU4eSUcW4lRXWnhfsz/cVOIgXTeG1bKMTnGjA30bhYXnbxIDvqASZajQ1YsC1Hpk/2
bo+FYQJO7Bu7VX89erwiMZS3REDZsZ+Tmly4PLTFQtGiJD4W/PZWP/hIqf7Ozz+dv/UJqG9sI0I8
C5U3lLENfuQZgl6MkMWt852Gri152SyITvN9sotG+KyDb/YwUATShd20eMIjZO0Jwsp7HuQzJMmP
sqKXsFaOZ2+eQjb7Nlr7hiYd6dXVPEXUchQRE7mBrTXO7I5S/TJZGHDjpgoQwrj/oU85xrANuJmW
ZDIrGiA8+I/5J+saH3HW7ClVuOm53o7hRZyghbT+YSsl6r217/EmbARP1rJB7wS/g5rmLr0Rjc5g
rftYlZtMj/HH8T2pAe/4OIzdRWQkySkOaWbOnmqfzhEc9JhWcf6T+H/YbtQOsfkhiOys+ydenvzS
riKddEFUZ3wqCnHQJr4ofIJT601LGiAgSBPyzZiVpfbaTI/yw4LUobqxFoQ+kBN0q/5M1ZkQSKLV
lbJc5jRDIDmN/+SasiHr5aWJ5pDI/3kBpIIKQ/PZCt9L9lru8He0Xsglp8Vhg8jaDYu1MM2h0MXq
mkha7ik9VRVmQjjE6nbgputp8HwtwVap4UeoBOE1JhauLBNmh0HdmLBokCGxydft+1he9q5LDL8q
bIseQa+tbBYqxjMkOKWa8DirJQSd17rmOB5+KekeH8Fj0xQFyrkOqn/qAnWuN7S02rJDFFOa68mE
fVVyvc3E4SoGS9AKWXV7fAJzpvFHVOuqx1WQVTCW0G79HSscCKfRmrMP0gLjF2PHoPuk7Hng/c5c
FglHWqZs/h3Q84sVukYwJ8g7QquDEEiv0f8kkuEpInm4nNsIh52OAPJ3HLHPR5lyyfv+guim9yjo
axI5HP4fbeyVs7aIwGP49ZUjcE53BPzRmllpdmrv+r0T1f9BxAFplz5HPO2OWHSy27lTniwKznRG
tCcDUWgM6FsYL/6JWaRQ+izMm8Y3ZlJgSZQHQT5WS7YT6l3k4c2pyZIF1X6ddwN4OvIczTiY6H1g
W9axr3XSMfbxELLOvi319PtRFCJZGnwmWnCUubc9Ap0ZME3QQ6AcHHGSfNm08teMGEtUtsDJUSl4
sO5qKvrtsFMp+JRBI4myvRzIjIBntdTtfQq7sdnsi/c+Jp/ZEN4h8U/VgijOkAc9iFTcQXzwelvU
ayOLTklnJRl9tSOA5R1qkDUSygh+w42Yx9ixnbmWZv+7ofUWER/eK1aiElbe4vWBIHN5Cd/YnHtg
oQnFDaXa9A8DGr1Je2a7i/jnZ8SzGb3kGKFoasjfoKQTdTMnLEPlhU1sc33+mzKXxn9yVVuc8qPO
dl87MHVyJK3JEqNpvPdAFPrAe3caoiIueR4JlIR9O7PmDeWl58d5nqKKrijB03VW0tVcHf26GLqR
2B78G6C3G6FLZLQhDnrjBDQSkbSKkc3IqJzPBJJo2pmMlqY59oCKcKqFWGZno/ECj0Ch9WJ8GLhI
NUk4cFHAKOzE0RzzARhejE4M7PA7H6QKKpd9IHwnNe33dVucAGFNaGDK1t52KjyNRMWuETSKs0v4
oxPU3KuDfEzxJqoLQumv3fbLXk1khTt2P7zEz/v94ap5wWAExhTBU0vp/0wY5l5VR7IgrbiUiUSQ
ZyHRve0ErZyP/R2AnIG9sKTX6gV91PV6KazSLlrAgo/Lh/EF5xnS+UcccydlZfRxgdfQh2tbFtiN
uRk36f+rxBZpt2M1vDQV7fvmBvd1Pd+O+777LFC1oWMb01D1loYQof2c8Hurbawx9/Vg8BwfI2DJ
mnuD4CBh/nj6N6BNtKN6vE7iiIL5d5seaRwPj/qjqy2B+QEypoXYW3n7OustodMLNqvVjCiT8fJ2
WHustEYZyHEtgCK5x+Lj9UkyH7887wAIC0YlSeBSy6C3GJ8rl76vxRAxVFwVLYoXlnWk/gfWwWtV
xk+luhkKULSvGynXAGKszQJjh+Q1vKBCfRFh7X06/IrOiGcotFqNtQh+iw3HtcHeERYVo0dAtDr1
giKgXHfKGYfUCfMnxJ4sJZLyWTNMIH/bi6DkL+C+bTxCdOXt68vLP3XzplFrSqLeKoAKTAeCgWnQ
hl3eW/4CA9hcUrwt58atcxek7llt4bKETguE9w5GNu6WlRYHQEPE4gzcwOOVDLS1RaT+aZU3z0Iz
m4rcwcEjrpFeR2O1bDmQKg+Wc2hGosKxblXPHaRAdjFe+cqbC5iCWSX0nki4bI6OeJcsHaBIlg6L
oOPImD+4VEgWWhsZ6AhxKIrkD7bnRF+/c1DYVBLxdfxvKpjR51PtumLYWkU+mY8L2mWFrAXm9dc1
MSdlxpKLNZCOCptzse3PoATKUvwfhgiVdrptcna57TU6mt36XLMOF4zN4skLkxf1Y53sVUROf8FO
p21sJC4gsOqaRRAZbwmhMoKDmNTyf8YYWnfXfn/ysIltHr5/U6SFTBjvkvUokaHmPmY44KGvBnbS
X4GMfINY0OtDdTDmNjatHW+4VlVjd3ZOe5GpCtdIHLWvy1u8pNZKAN0znCFFfct+9e4Y/0F8EPUL
wdrtNvfO9/FR+dFUxbh5ejbzTDPTZLlf5J5N5GZKMI2xAkQ8qOiJznlObzD6dHrQsQsc5VfQLCN+
WpM0uCx1lO9GwbfX9B7Fcdq2Zk1GZIVBv0ADxVkv24RLOfd6Gkt5uI5wUaR9KnQPVerZhdsa1E4w
wnmaR6uGgiy5HKb/rH37nfIkCj4BoEBU3ZH/qO6cBGpVgOm9g7FVyYkk6xTh3kYWyGwC0htAWI8O
gk2Ssu/C9C273C6CwcuNZ7PNzsuqlVUnejGMLM+iihKbxZQvelZOZ78vEnNnLmtX2nxv3Mk+EnfW
sqDmfijLsO+9xJ6Db+jb8garRoQfE05u/Vs2NghuTAg6HwazhImsIzr4gcgzUjtycHVbRwuwX1U4
9QWWtjcL4Jxf8Y3jzVl6ix4cMOy60IcZEf8kshaX8R1l7gg/Cg68nfGDElyl8Vk0sjrlEBYj4MFR
Cgx3gC/p5dzJaHY6ubKfYWOWjSK5BSJWcGLRZ8wf31Y9D8C06Hb3LkIe5uldeYJ/c6tFBteyddGx
IhNwExyh9z9MuFEYf8dnpkMsnh/cLMRTuTcgWmp2jYHjHxforUrNxZWENVqIlzgRBgA+5JRogc1w
KdVNJ40HfYQdeIHoM8wS+QdFvxlUOR2K5D6HPNpZ4zHEw8OyuwXRzdBsOvupD8z96d7Avl89tFh8
YGYeyN+wzj9WmreDkpYHOIJYFJpVEMuwZQB41xW1F1ZePM9iUewGFo/MjZ09h99cXuzoM6hZ6B3d
7w6GlayHu63ABPYa34R8PNnZtq+pNSg8mro17kNCDQSf+xuNrgb5mRgTjyXSauiG6lQWj2azO9px
f0549CMhQWie85v1AtmiQEbnPHDZi1N9mDNC8INrMkw9MPVhpP++SDrf9V15UvfUpiK4yHv8Vfoa
1DwUqHogbFG3tqawgk2w/3NfxiSAm6An6+rRL6GywAqzV2ZXpWO8OMe2K/vOqPAcUxhxLD9w0gkj
D/rPcc1oqdPKGjIQyldrZTDl7tZrs2rDkM/N9GfGBkpWfVCILSGmpa7Y+yt2hF1/cxwgJNND7/rV
pUxSiwUp/AwbqAyI6JYTKdkMcJy86je2jzHw52yarxYh8xVQH7UYLjtrb+aV/h42t54897k3Xm/S
Ag7RPR7DuGh+Gj80pz0a2K8gt60uO6U7LZFFxsliww8asJ01RNnMEfmjAMe2X02k11ZAAa5NNt02
OxPxw/+8VsadtlEo3SUGWmaeX0PkaYpUqBRqHwY/X20fbbmle0N5JOgDvloFaTPNIGfGAOJ/veyw
Hzi4bdJSowr6kIQRzyOhQT4HmfE8JbNfmf/9hIPIQHSdxNGleV1G8eiqA8uwMT+CAerpWgto/fQ6
1Z/l1qxcNMXIrS2mO/Us6soSdFxeWKosTKNyFmTjlcQqgK92/IBncgqDeq0CNuAv5j8MBBdvQGEn
NHWia0rE4wS22I7Ke81l+JcdD5GSbVAK1LldWvS3h6W0RI7duJRF9TXTtRU1yspKXvIjNMxaGuBv
pg6kWLk6yYJ0B60WmVbsvcHeaFiGgRwfNIHJG0QSaNg+3w0fwNOCnqYkTcqCBvMdTIYH/xqV/Wm/
SOoq4Qh0yeBqevyNm/kPksF1GqP2OS6teMkipCIZp09tF6D7rylBTxeOfkCzA1uFDzbIqL1ZZ2oO
+DBP9ASCG8WIXL/nIB+GB9n2u5PugJQ6UctKrL6tA8byZmGN58oFtUyijLMVs1YM6/RktXlLexUa
N1y23RL29n9SnlH+0hO13TmtZEuOY/oPC4M2Y1/pcSYxin5uAdZj0yJomO2B/nTUNc8+pAiRNKgw
ltJcSlRA0ZrIOtmQYQveGH7IBGCZJTRmspAVNhI6FHoKP5n2b2OTjMFJUPTYxGyuD0RFY5uyhuOg
bOoTR5k+HkscwZwLh4uwCXVw8CzXvP4I9gSSKsoBoaviUDWhJP56eiqY+1ColGRMrrCj+SLfgCbL
l1MGL4lOd8SFWKq3Pn6kAJxCtP4ugjjCBKIbR/Uoke9AsoCSctiZ7/sqTnPefG6YgCmFBNE6AAG/
lM0BMT7zRsWz2QAI/4ctjeqFrgZrn9kPdeb00hfxtsm++wUsRWCbZEyef/lG7Yc2W04LgcZk9tBJ
VJSWkFLI1lx65oCfb51+RKt6dgg2cBHdi244lXg6hM5lLyHpFJyf2+Ttxqoq4slbsrtD4f3vZ/6H
mznQasucnSzhonqt4VQ+9CRkGL6pXAAv0Bbr0OIoUcACL5xFAq7+XEujY5+rMjq5xRqbBmH9WpYA
q1W+iiY4JjgL8izLsuKBP9A2hgnA28Mr5mxfX4I7fnPIgPDoCdtU/U7bKo/J40pfZINHpR4zCwyA
pKQnXhsEGCyylNspFiU22/JtQUXwupZ4vl8zBpLK3KUmeZMJnLvIdiLB29VMirLoRJG8urCR3yRl
xx5MgPWzgpfTMzKzR3zgVqszKpNOoLTjsAFXOqr3aS2vzwyHXSIm7SmBldZHJiKLmfWEPb8RUz9A
f51zBNWboSYCtmfcJPaM1YycXSemvuU/5r2m38KYCEjwosxqqChE/n/M5l+0lr8M4Di/eGivc4+e
FBf3MxlEp+ZBIgoJC9SkaT78wiIujVSfNujn5gKYLkR28soS8gKtgD0VbC3oD5heSho+qH8kZ9HO
8Kp8FABXeB76DGU1CtH/wwMQ0Zknf4feT+JP4f2fXDsajCnlFF8j1l93I8SuRPHkFapHhSAgMLDY
HnXR5OKwFs7YhN7A4t8mPJOlcz0oVK14pxuiR9tvvDr+ncTGEXSq1hZL+O+xySXw2fB86ZxLxz3R
Ka4hPvNNr8Iu7wl1CYqIK1mqI08bgVDVT5jKR5cmpcM8OnP8Z1Pnl0fRMpIBnlnnGp7rM+eXifm5
SzfF/mM5jngUGUBKCAyXjioGLb6/RqTVm3S+SXWcew7zY6bIPo63MHSUBKppZ9UFNMuk1rXkdhrm
psYc/Y4SLfZVFxF2utK8Iwz4pHPy97wARMMleLlg9hwn1HnXMTH/EYS6lFHYxTt//0Y+HJmcpagj
GYLo8evWw+a11VGARbGwdVr7oIQp6Z8tCa9YIOR71bVNCKowgsgJjzvVICGdF37KEEEBOOnZa4ka
Qh7scuIZZtbv1aSdtPACgiuje9IDRG/OiKtgb1u6qqTSbmR+c2uouMUzpOvEM/S0Xi7sd51Ve7uj
UvM/PInfT6qspDs9O7dsGYi94AA4Mdi9ShHGTvQReIxbKve4JV3I+vRrVwloxLixnv/P6ZSbCm6K
6WlUbicxRk1Ep0CDPYFgVVtEX1TIQZSV8wUQ+e1K3kkkcZ4+XN0go8YEv/onEOzcwN+9A5I4fxJu
rps1M+FM+paq5njhrzSK9rLioKmicz20LjDsroMY3K4hUXaxHoxebMfV746K3fRP9RDQsuLLKTpG
6jxZDPMCelhI9qkmnGtgy2FwwvjJTXFLlFleg4FkOXjElu4Lm+nWYmjXgYgE2b3d10S9AgYLyw3m
KpV2ys4T461xWYbEWBMPucDKq8DK4xlWLlSJEUCM1xwPyEPJqnHElu/vxrYZXQAcBYsQBdV6nQQS
QRydx/4+73JMLzdaMhlWLcnq1U5jjw5m42UFGH8He/mv3FnI1cFOftbgGQDV/HILSqNy9148lfbk
0K5n0O23s/ddC4F/3UEmaqF7KfWgde8fIQhKlwYcQgseIVH/ko4MbFiVcxS+x4QoUknZTqvgxW0M
VLsYGoVEVH/EjRIRSAxqVr609v4TI8qDO0RpZxZ1Kc3fO/POKRRst3dwIh+g3FXFuYpQeRo8pqig
CJOY9oSuwykP0xb+JjbdRJHbLE0H8vC/uL4o1YwoQYhg8oma0AzEXinP0smO8GBlGW5uqI5ihJIv
XsVTl7HMS03DuKcCWf0g1vTn90YbQMqwF6L3+Jwon9FZfCHO2f+TKC9o/Ra0JYHCUT3N7lhkhi7u
EOVSNUppT+mKIPJFYp4QSjDDIURgVeAWBAQG7wF2VeRC8Y97zWcVaZsKRu1FY91LpG8bbh1Z3dvS
hRLfvcKerCfW1HFJ3yDaVHiaega+V849Q/yU3OrW/e7SmfLZs+1z0G3bSLndMNnxqV40xixgceBv
nmnGVCHN7jhpUtAqEtLpGLQVVvL5qtSNn0dIQSa+1v/q/wU38M4qfBIA7XpWxrK0boMddnd0p7k0
2BmkGMzy7IyNWIFdV0sBILzz/lEZGvfpjY8SrJ+VeZKmIiFJMIBp3MOpcjl26EQBMJlYpCuS88YL
ENAmb3pwet7Oiiq8MunUjOnyO2ugPvNWgtHteFfkHiF2+wbfFxLIiEWh9GM+MzysGCyx7nkKeQuv
O241SxctkT3JHf36w80CXuLELa0RcRemi31Rnxkg6XUzFvlRMKOMVijj+qOvrHTY5Ku0t+dZboyQ
aw36yBkwGiWZ7KZQHgfcJCtsHKUGttcgeUagD5l8u+2Ues+1WJ3lIhSLCGvOa9HwEAxdBeb4vXe4
1AK9RxabuNrxDH2FyI6wuJvaqoXERtpxRgJziqMHiqu+OL3pGhCB4P68X5cdfof8pbc5ucrINjiE
5/W6uDxqOJ/dbF7mQYmNJ+fehB656folYW3XPmB3CHH219XDfDz0vIn//9s8TKo3E49L1L9Nm3K1
9S6pJF6QA10BMCi+80nCXLokAgBsd+DQKSwCMslxr0s8HaD4pQQIft5Sdhf7BaRMjJtk7PVEl8OX
qxPOTwfRT9zYz7K6DsICzBxzG/7qAqjnQxLBBsxgtgxKEZx+qS6hVQM5fFLEqv31NIIu5/WeMfOr
zAWBxlpVcB/WonjW5gCQkbHUPACY+Cw/8JTo30FRgL9Sx4bIPbYSntBWRBYzrsV22ZrvtvpVVe4U
yuUsZnAHS2d7i7gjxfRRzZkbiLAQMBiu6ju9SjOZXpPrfmfeKBu3iv5HqWY1TQNVqxie3Nmz5osr
Lr7DtAXnC7+je9ng3W9XCVkET1jFO0PWVkdJsCU4T7XKHxsqE4OGIwksaIdf8O/8QBSJqFSt6cSM
oY30QOLVtMenKBDmoxy3Ap8OVCyYETRzCQXD/wKEWGMYoDiXa3gsGpQgdLpkuFNqwk+kaKfjUOOF
vu8e8duNgIEet4++ErrC2ERn348fNx2a6QYCunnTNVgj2hbkxN/3Sx/2K6o9cXOELblBkyRxo9Lg
1qY6oOmOFkpKbWMuSpdgA/8/UBN2lqzsMPJhupSj1wZS2MxkyGlec+EgOOz6BB3X1pWVnJ1U6j1O
RGf8sECbCHNY4EUuoK8p7USTpiCfTFrMk63E4o+HEXmf/9I6bhvMGXkdAPkuODgoaGN7FXgypP1Y
X6fwB5RLo3r0X+en4cFtvDFvNADcmdonETTD6m3gZNJjEuPzg5hdvC1WuDoGPOz1+U8/TTR5sOlc
hTkjGXqn9A/CJc3Hb10sFqA3JlQl0ARRtOrv+hH9Tl+YrUztUVgigQsghyqEkFcNpdQ+iQwNhpse
AqHnWUHbxr47NQb2Kmc/YK+xljAhstIXYr72DoONzMHv4Ddco4ysNUW7QnH+xpJLhPIXBKxOPGMI
jyJMBA8JCO0vPnKb9u3USOJ9CvA0x3awADlTUOaVVTZ0cXLGv+2s8awn3fDK/cJQhUkmL/uE55xt
xMu38p4uM89C5+jmmLcdAeQS8V+Jgio+Qx/Dw1mJiZ/bsPalqV1YrWlw+HJJZcqy+PGP61eBycns
pI+k5r7n0t+fgmem5eo4IHvGGHGO1aR6lF8yo3R3gl4kCzT4XH94q5Rb1UQskNABMqLuhv5VIDxo
qBZ5RP2gSCzL9wE0N3DMx8DTA5Wzd8nw/HaIG8doeQ4f8AALygOj6ueSFzHcPaTS3cUS1EC2MS2r
/qtCpGFr+mNswkjaFDRzajvQdjcTKOaN7cLnZtL7dX7yAtx9OC2cywVxNOK8TAdO0OCvoqw5O1Xd
lcMelnxIV3uFk55jQ/vRyi87JlqGLkUPKAHB6OKJOI6aE6IGoZaWrPZB1mXBsuudL/KJOJU7LpIN
+Zf4iFFTyj8svqN2lNanugtkC5CAphwD/SVUI3OYSBXF+VQ8CZ+5wt4bnGKhWE517mOXdQDh+bKk
iqlDtYweDrGY/Mlt7M/jp62zQTjERvZz6Yt2+jLmet/+F8lldOxBwdBEFUm4fjOLyk0naHX8GW2N
StdudskvL8UZtXjsWt80Xj85d9VzqGucGU1ISIHJX42pPvec5BW5jW++TpZf4i/cDbqvhqsdC8K1
1GYzJuecsoazklFCxgauKJ8Q/CLxnbqggap9+8RVmeCcdQl1II24fg+7dhL2hToB70p2AbHLYXaO
MkTHbHUzpLg8Uf2r4+2gGR2ArjB0cgfKxQiYEZljcumhkVYXnUE9UvALyh2+4iQP7ubWGw1pDPsn
hVkzNIGg+3NfiCOfcx5nj7frEKtpFi9a4GEcox4kFFprXYr9MLSTCleVYVtTNH7BswJYAzIrf6CG
cztGzYLHukdSzuxSzx0LklesV9NdcK/8cHSw2664HTZEd9i6+YG84gdiji/gWcUGz9uQb1d6bAgu
J7exI1TYXdyOypP7PEUaYqA/SEJS6B3xZGb9l1LEKZJsjudUW6xxTJTGihHe7CLP7LRxsieRMRml
8ZWAzcIpVTiPADuTDzUJi7mcTq2EE6HA0kOCYlG6CLDDM1Knv1+GZA5bTYdMur/RxwmeRBzrxp4U
kSc9pgD9POYhlq2Cqs/R/OK5FpWiuLqKE3o5KUaAw+CADCFEZCAoSLDYkunbq5bJHIyXrHdgZQyt
+udvrUdeXMX9gME5uWxcsO8MPGUj4JMODFlgHf7t/XYd+DH+g3qN5FL/z+GBrCjLKA6QJEo7GR6d
TIsOLLOz5qwUK4oRsh7gIC5ZdkQTNHKozaoA88XzXW/j6pWmhHmncuRXjI640VEzHLZCa7f8yGi9
MVEuZ63jdJ5Q9+1458Tw0uJF4kqwlBptkLE2i5e6pzvXkE6g5jyVFzM7wRXrms55js1l6UFOqMCd
9r7XoSvOjxby2Pi/NYBf4JK1qEts08xtgFX6U5Syqh2pjcHSFOgvdgKTJzb4HVm3VkJW0dQj6n67
KprJa2t7AGqTcylJybfgEFp43HRP31Hj2UgrrZxucaenbfWeOrfhsdncHF2AtUC6mDYEac75iCFD
D0YnTC5c6V0TZaUH6H4/qeF3AQAk4mB+nvxkOEzKbFDD2gW63a3pXrglcMFLxrbkFBA3gOY72GlJ
VXIti6bs1xr3zHO7niX6gV1rTkd3+J51L131HWO632275ZbZ2AXIPt18MKglbkmHo6PQGRAjMlfz
74foXcMTHG/FpEPevAwdKSFrMggEJlcDliYu5AG+TQ0AaodYhcNomfsl8AyMGm8J5eniBvH/igKx
voJLQQG9h0LlJ24OlLRN2HH89E7q8dGyxN3ivpZahIu7EnlgNPiSuPS5hs1x4OHjbLRur3Mi/uUe
+qQwdagYR29Nni/udSJZO0a4sRHOxTgkuqFAnEUzor8rr0jYLN+/NfGkmDm02xWvwgGDiHtm8PkE
xQBGCUeG+IJUhgHumqadKGieH7MXJZlWyBZgZV5KJvpjMANQ8IBGSugwam2mf5yr029DtLWNR/g4
0NRnJqmeIWNe5C8P9f39lcd4++g1cjrXHNRZcmQUe/9k+9TY8McTQgmbblrjSuQfkfP+WHZAaRnR
BWRgVd3pZGHezS3GsfeyLumIy488ht8zarKFjshF/v4A1kcFNezlRDmppd518VafMTQ5TeNoJZIQ
Lg/uANWbLfsyIks4aujrs2/1pitlVJIo5h93yrSJ62/4D6YzZ+mIpUVaRJ2T5YzmqHiLG7mJC+g4
d0dcE8I7PFwWXTNatfT+1UiXoKC4gEdWg+IykfKlmzzg31KxOmvO1b5dqsrG1MLQC99kA+99QxCR
I5cj9s2Let7Oa1Omte6EQZ437iyup5qFhpG4F1I3BGQKQzPAevyAOAhISTi0HxiCFwtvzgbwGY3w
bk6Pumz83plcGn5biEaeDiNledH/+eE+5CFNX/c3ghSB0biCnvsVAtLxU3lTDeEPqPQY0RMomgdc
fYPvHBnJzpxuUaS5fomEiThxS2Z9b6p06nrMQlDNntQ3goBkwxLsTlcESW2uX2FBIPVVdVm26xvO
xxEEO+KHtlOMBPuHy/9G1riQIT6tw2VptY6QgjN2Is9q5T1IRBr270MkMh8q+XxCO33zkJ5TMAF/
oLlcueINABph1BbpzssQ/nzhEtThniwwVg9GEotYgyQ/Vf82ZgvcEoMgVqcadxWiUopZEeOtYtuR
kgiYeGrAegOPIadFGAZs6MZsvKFdls0mwtQvS0citthTU5rQJ7JDIV/JyZ180UOJd6NhR+HV23bh
JsD+4XmwcTJss4LToYIvnrTby+A4N6vUmZKGZC+FpJ8WKYWKntyurWaXhMjULq+jc/uvZ2++f2tk
QyIwyX4vvAh63hQO6bwuZ10NIVSNRNzOsXTEsNXnR23LV8HYy6Vi95mgY16fnwUGzRKm9SY+xcru
vkAaDIIi6sCQHONsYpoxPkaTEIGmfDAz5T1Mw6U0RU1LHXcudmt87x2zuOZ+Yig5Fr1lfuxamWwH
9hlNMQSlGwMt2gJhA8VigdYUsE4RFJ41ubQ/xO0tbUie7oAXZ4P+UP/G1THXZCsjv9uWnd/vZJp7
RL+cG5mytXY/SXiheToXq54st5SWIDtGk5Ihk++oZ8L/ETpjvkJ5HL3473t95TOypZWbQotiGaLW
HU26+WrkCLJ0nlRJgJFWRvq14+4OBVYBIOt4cXU/t3aDMTN2dGb9yTThuYQMQbZ8kL7QJLXj1bnO
mz1mdnOQaMCy7ius4809wB516As5OWgvikGH4RcD9y673hl/veUCAulXIkdQn+wtgD/70F4uDvDE
ntGqf0lGRruzBGjwqZmV+h9qpFj3JaGlqd94yV0ccm1vtOBHFnY+C14jjkXUQL/QbMoLRg0e6LeX
VHQxHykjQusmMHa+pHOg2Y4r/7pLW6q9FE1eHx3+alpW0n6lkwY7LdLrSFH+WWkCu3qvHI8xakXE
0QS2pXvYDKkqJOaYlzNZ0Ld10OkI1DcHV79GyRLoivMbT07e+WzVnmkfIBKYmf0DYbHZRApGtvAJ
OnZrBJJy5puOIqmCw83aAh2nzIUr+HFOXws2A8ULhBPDueIect7fLsF9Ylmm9kv+0nd8H3qjSLiF
HY0i0qZ8Q83fzSzi7bTBoG6xBRdXkbFPKWzWX1HuzIZWX8AUw+tda4ZeNxsTjefpUlVshqGWmMpa
8Zc0I21GX4ZSmE/yGPiJoQE6q30txxk8s7sU8hluVfNFepQd+FsPMhuBZE5fwQV+8OQ6f7+ZKB0Z
r25rru8kRbWyXgkzk3P/8Vz0iXdoeYj0jNhxnggDfyKqxioC8UWPCfcK35yHVeTk0hqkGCNoizSw
CBBb/jFZntF1ueT8iovR9endmJboBeWaDtDeG/6FWnnBZlQsguzlb1h88ut8am97rG6V+o5V6Rlw
se4PxeGAKEFgHMAanP6opImcbuDyzVpVBK7BNN728URcVfIM7SfBT0fgbDZ4SxmYUu2oVsN93tZu
j92yJS9dmx4RIlUcXhrSscbsQ9K34fS0YVJKOVbHT7krGRiE/wqMPKvMNQuKxnIYoFWbX320iwpY
q/GI7ZXaz24g4b2ocqy7jSKZwNs5Y87lRVmFWOoNpMrlDFu5OVdCceu7Y+90+vmSfP4CSHSVfmxJ
4SLb/pTD0VDjTVY2x1oZERV9WwCK7b/UtYbG3+dxN4vmGI00HYJU4Lf/iAOH+jzWk1BGOZnRifZb
ODuvSlNUIi0KYoUZaxm0u3c5mA1WbTIdhkqntQ+GKIwnbB7ZZgee/uO2fiv5MyX4VkVqRA7lG2Ae
/GuunhLm20EYAk4D2AW86wihrMsEJWJfgzKAqqDxb1J6BxDFZ86FK8PIE/JFXo8+42aJkbhuyIta
h5RDzafH1rkvD1GDxJeDAOcAhKbx9Vq9lrhFfO5tUvvG0437I1ENdpFrx4moqe0cS4e6aCIuRbjW
RE7OYXN8+/A4iXeG7nhc4o0jqB8eb8oaSgEsJtFBKy3mlgcWEZwsBj4SUU12SUJC8+87dZI/nkDY
EroG/+Fqml9GrOqbJNPNn8f8O60u1sQ7g+EBowLLzoAW8oRwBJzAEj1NtDzu6oHvFJAM11S7PFnN
0MrHEGAEImKAkILy+aG5Sc0ilXcKgbWCmOxOukhkNQ/ltdTWktJDoxLB69R7ObUKfJ8/mAIYMmze
Jd6Lb/A4njl2DTp9i/tI5ODc3FvNodimRPA7y0p9+FS6UnPuzVV2El1rYqq1Ynt1sUCSk4EKPhRU
024J4z0d5z1kPyFKThnUn1iFYQO0FFIzqAjDsfzeafZCTxS/Di2kFTCQSuJ3cl7UnZfciLPcdub2
dIhxT/Q0/4S1MibFhCKMMKPqnLML1LRpT4R8jAmOwD4Kd5xLVC3kC9qRoXYKdL4c/POnJjO5DxDQ
ZxoEIdUzXRsdoK7zYgkfSwak8n1V0yhcbNgo/pQ34yHX4B+VuYsiy500LJrnf064M/gQhi+LVZ92
hRSgx1x8pRWGqhoWlDaG62bltievziMq9j5crnmGmMWy6zgh5NNB9PPYVLqEsPibyziGdhVF1Pva
+9dQZVQA07UAxPyBKL00+abSxydH5AIM6sfM5xwhC/y5kaXlSgaCd/e+wKqJK+oL/mjFI4Ps6AXX
seMzFkgLMr+IlS1o1cB/lGTwBiVKbwRNh9XNlcGjcIl8Jlp9nY2qBuFU2y6M1pWOlwqVKDh4k0aQ
XbxKWhmM7AvYzAQiG0Iu7YwWscSM8NqsE3dC6+Kv3w8cOM73I2jvG1MAcZCNqQMVMPdQ2EX1QiUG
1tnIXiMk6qla2vhxbqXOTyUeNXkHNheGTWbZlZGtsWsdbyqtVxpCosZ/XumAgvEwPhipkgZawLCk
kcZuI0SeVo7XIheiXhaurhML+WwzimG5h667LnpGrEVTZlm1Na0JwXgMkN+8/v0V2x1Bei5vk75P
MT50ssEIGWF3f+DIKp1M11TQLcZKum8uuMvXE5Kea2YO7LIFIAth7+IS1jxGihNC8JcrfALnmd+H
q7/74SwequO9OyzknuQwKMe04VFqXLy6+Vmf/4jurLZ3LmbIwFzT4lwUZyA6RxXMUAaXgECm0iTL
UvE+N3bwVy1/+C7ROkwdPsLOLhTaKiTnE3Aczk24Y09KwkevpKPmgSaUojBIgoNo+WFzQkgBzw5G
m8jIE5zkCHAN/ok3bsXwGUK6tRwclTcu/jDbms8+4bW+0V/A6o+5y9k+6J0ZxIHpZEBL4NgySL5v
iQ+3f/Mj0fxjZKlIjIpbqiyWtBmul4HhsntAhu7mQXGcmdejQK6v/oSg0WBloZ97jlBuNm01V2hq
8OkPjtOH0NfDJpRqKmBSk3Pl7nUMwghGCVZ85AOr6EaOnkMKbIHNamzSUUgs5JNeE3BF4rHQZuF3
aDLiAY35TMm/hjyL4JAmPQMQSn5lF88qO6EnsCou+2IzVgPhISfK3dklVYfZ8ymOCKTcCLIobbX+
OxOLqyN3bCi24MMYiz6sxO1qO0B6oEEUhDVcQueqoXNwuMZ02CM2F/PPQYP/guBOy7z3sbbpwCWq
77u5ahuGfThdtZfQ00mbcoh4Rja4Krnhz9lp/4/3IBE2m+cgyBW4OP6pL5snrOWUAYXSQg9ZZwf7
yZ6Zvvn7sISAW1mdEnWOkDuqPGcUPjI26wjCz+G4yD5bcFIoMYJKMzbhP/Tn1BlEXgxHItyLikHH
+c4tdg/URITFDrLpmasIeHHG4JGh5panKH0AygK8QS1getJqiy3YuOny8uuR+kMrEj3GZ5Hk7PKt
euSVW+xpl7Dih6GOVKggb53ufkcyJr5eAyEt3zKMpbXuZFROQX42HKmqjT8+olyvjKtF3Yqq2xdz
w06rBA/WmcijqwJ9xW6eCYvdbrf9zsJMMBy1PwS+SidlTtmL6XKEoIZgMiUjHbclxkw/qq/A0wUs
uuQzYCEK3whLAYaNZyQ0wvK2l+CfUwnBax2dCjIwsHSUKJrmPSja5PyCOnj0lBNFlT6C4niJTPlG
m8ZpKalS/8hrhyBUEq32WsZb7zeju1zqssXLwMR+fZXzFOGCWPhVq4CJuj157YqaVbtfhrb65rc/
yCeCGfOy43ERNggL3T7U+9yupzSm0sDSin2l6bDSzj9uPSMXdDHn6yYIpoc0V/JX7Hg8ml8gsr8N
pl68K6qG15HDDiBSjef5hdjpa9HiOBW9OCeydB1iSrECOrpXQ7RckAgHpQyFqh2PUAA1gwbM/8Th
M6yZBrjAqtp7HZj/k0ko2L4c0h05/mRv7S245zNaUqcf+AZAf4wQtAsNeLQyu8yBPcbOprKZS//2
rjXl5Z6pX2XL9Fle7uTf1T49rkB0iQ7KPsaXb7yDmF77Jh8rit6i3OslyYI7prhaf/3gMh3F7d0n
VN1bQrcqP/4GPKejr3a+pIk3lujjXXxyQfbaf3dIKliRs/ENV2fmImxIEwd57hWVTNYNOkEhotAP
0pjdBj2x3t+rZ0OiruULYM/m/yFQiFmOexXPrg0W5FZkb55IXIc3N63q6U7gS95LX3YzOGtlvJI2
ullUukCLvOTZR3n8wrUygFuc5anjAD/zx9pm7vy3+lZMbVqkg4lRZ46ISW6kAllbuZotnQV9dPaW
wXdricuANmSLy0OVBlyKB6gqNjrtN9IlslA8nCfPxK3Vl/2aq8k7D9dDCAGuT+3XwwZrqyJNY+qm
YCfSiqPigZiDrCSir6fVtwklnsnPeAU/5cwSuEj/TE9S30dBV7+usOtHl8XRISf5RqRAguDhhMts
D/R6K7YgsokVqJNxcoWh706poM7dJnORekk+PxFEMPznginldhjuKRb2XZWOnhvkeqVTejrjxCUr
ftANHLQ5lv+NoYhkfjE3J+btcQ8A7H5wxzQJ1OGMA6mmDNp8ataAIZU3a14Tvu7ISP34qeWbNrr9
qxv5F25CtCB5vcB1wZ/yAPkpVrypq2QurKhfABWcOeM0YwlesPWVm+ehJBFYOoRhQ+Z7r8JUHK+B
2x+Ayrwt5RcXn+kTp78wIfJLKCX5JTKx/HXx5t7YuwlsOJaBXLJ/VTidGMg79KsZ01kqOVZWTBK/
c1XqrwD3OI0wwjHCpl3NB4wlJZEHkQSCKNMPshNCRBTa3Y3eCC0xXisMgozCo00iVcFvY0q0wc6S
0oSMp4u/w2vzlSSMC35ONgMrZc26ZdHXllnvJoHvrnTdRE38shUJ/6OmX1NNrZ9FvPo/mIAMivTZ
O8olGCRWp3xLSRIddynFpcawsnXQ/YIF+eYUX8qleL6UZ/DAsWyoOzu40t3USbwF/h+UxKe0Brsx
Ac639tK+CaGZU+S/buwYeF8hjiciwU31PLJaQPd/UMDJND3FX8FkD+TiptJTTHhLwO7AGRtKQVRj
anT1PIz/yarIbYcMBE241M6W9YKtZoU7RTNCccOSa8ETTYPMRyOEbzEm3WY06QE/OTzT0kRtR7rR
YPGeaYA28NPCjf9aF7SSPganX+flv4SIIHlSclop5HuPb7Q70qYXrUhfzKokBxYlmJbH07VSzT4K
/Y9wWdlBFHaCsm/f++2MUtHV060DsHQ0wU4084S2GQiYwlyS8WsP+pVouXNU4o/+AQCFSEFrKQnr
sI1Q24jhrHBDwm45gWipJYeSrL+t7J9rqLVIKl/Vg3cVp2atLj1zi+IPQjacAw4HOUknIByGplHI
e115XhxbTPienodztLeOKXd1Ic7BLDuN+iAMk3aBPoJ3k4lgOnSLs7BUmpvURv4BCVdN7KaGJTD8
arCkJRFu2i2svoxXIiipIIAv26dicn3xQP09CBiXAxTUxh3+a+JT0gpHOVBvTEtHsfyKF5Zsm7mK
TmBn1fnCv8cvo3pLk+Nzbr085nnY0WB7tS2mvMPX77p4aaVJp1bYCJ2yi3RHN8XzPBYg9y/Ucbha
aM3nA2g3YuolgX4jP5IA82B9gpqirL260F7t8K62Ek/oeszcE/29v+mDG9tgVRrhPPS8FJCk+wvk
z6ItgSSYH5HgBn6p2ka87ymgxnM11irr/YNulFZSsOsnEzU/WL1Q/DU+2lqXxTaTTlgR/muhxas3
hhZevA4E5UQT8VdT9UvnmblmiqSTaz5ub+cI72Ty2BG7sxJfvMb1lmanjmEyHoaS5aOwaIJqUuLZ
3P6c5EERrhu8p0FbUKIxtP734kutGh7sohnXEqRLFF/tpnxiaUov2rcrrRm/r2fMrov8myeLUl0z
nnjrEZLSaoPx4h9UWim3nJDwY1qKdtFTmEk2O3WtUclnRei9tL2ikslbyZQlzpukD/4+3dzUhpkc
FIqvOSB5f3YFkOn/r74jj8c1AIuSU2GB42l1IgxBrW3DrC7c6FG1fIdSiHnXmlRHaZPsllZJp2EE
J/EkUAb7wyQIbT0bPq29bD0tV3OcoacgmkjiS3m4OoeAyhBDxXCM87IrjrTRoHk8Aa//BfsaStvF
h034V1kog8VxrEzLG9FI0MSWqE4BMpl7Ort038Z6fUZO+leDDvlGKBBuJc9iptGF7WV2VftIH4sq
6mb5fE6w4uFCm3i6UWGI/mE5QjpL90WXckDT7XxXz3VuCO60qXpTePEfEumyo1ChsbxlZiGjNjSx
JYYIIAWs6YOs8UDcdt/skfZ8KE6imU23aW3L3ZvU99d1YGOR+u5VfNcq1KbK2bzDmQWKW/THQYF2
cpTLBEwIUsHcVp6HVZ5o8AErgf64XEnsccfSFRIzjdRDE4QgcYR29VBXYco74yropsEr/jmv8RW6
LhY4ORbbYGPEJ/OUUDCJRoKtKNlvNbdWGigmTOJbHwvR0PR1qammyviXULtzXxZqIlssWwQd7CBk
tqYBD0GqwV/w3AJ84oeF+UbJZLHikOBt55GLjAeKv9R4fPpQ3W74u+vIz3owao7iL3+vcZnINHaj
UE+Zlrb4G19sRcBGDyiV2fiKuFdxJiHw8MIYxRbDIF2QfbISkOf73F6985kgOFahDBl+9VSSmGix
GutEqROAhKVIMmtCuS1kPJ4WKll5c5HfxFYpqoMyoVDluHxJkQ/7TP5gmW8knfrbXAPd0voExkIa
F+Il6aLnHUrdNVGYR9t9+sCERTWmSn99DPdS+V6rUm96f+IJW1JwWpqum5sHkQ8pE5xJZ0IbS/XK
4NjEx17kAB99hK1J6qOcBUJj1hm0NSlamInWVIpaPfRhbr3HL02YjsbLrXNNAduryJbou9T6fr4/
1FFjZ3LmpcdVlIyhUoVSnxJAeEGzX4I7IxNcjEYD34ODv3VGS4hNiR4PgcORF98xMwgzS1OHdwwA
OZ2kRWlkijls1BIieuljQwwxb2+w0zAUnQy+BlF016yeHxDR9zGA67cmZjv1bBxOO0iycVwCZKpY
HPEIlTDQHROHm+h0ILP7Jm5eAq0Hdlmy5XrTvZ5sZ/i/A6maiGOmV+Bk7ZwdDx8wjNbtMlUtGRvT
rgum77jM/mlHMKryjwVs6ffFV7lHCY17Yf8/FM5kSw1CDvsx/FTSq0M9PQkOS6DrI4NVs7lVuQKn
i206bVzJcrGOzdZJioRsnZ9l9cfuMAThsqiPLd7PUEL2yVYwvNWMk68laHp5dT8MwiyqMvVYuT2t
bOFn3+JBms5QeiujCZR0Yk7xCSSJpPHtbOuxdCuoP/FXRsMAH7peS9hVy3yFrAs9LOnaoSngtK/7
/DoqfK5MIg+XA6C0hJUy+tXLpYVswcvGBUlNUCd6GpmOI4A24iTJq044oT2xP+6/NlLsal4NXUei
ZJdg/mc8Ox6SDnNQyquojrAhuPCPs1lxmilKzFb7DqLwBdN2ZL9vuLQBl9nTL+EHuBiGRyGG9uFr
hXci9Il96dqkPiM60HehuLZe4QwCJUzyPUlExdofw/fLxMgU6jdS+u2hL7qftR06Qf0bvMSIkH/X
KyQb4i2K0x4A8zwKuB2b0JbIFIfAOx75pPPmCl+iQpM3j9ZefefYBORn3/CI/PBTbEznqQBuwhN2
PZqwizZm09X76ah5i9w/0I+BNeHYZ6yLVLcvD4KyiAi79w46KtN7FKlidzIeFWkh248PYeSzCs2M
YVwgxFUECbiKUIP4mOairVZ6Vr1W0LZE2SBRoK4gOV/+6SKGwsHqbcqyvHjHEGfyHKj8W/qWq7Jn
tPxYHRalOFU0W2HzNa5UxpgeOqlAs05JnRPpit9aaii1MMM0gMt1Jf8HajfDKkEEs1+C/oGI9jio
6H430QU06Z8p3g+tsQ64iLpoCLoJnP7HHuoXO0OeOXaHGU3yHT1a3hrWlBhQ89Aq5rivopcPif7C
3fCqVskzNWSH0AGUxLTMbp10lrM2xWdZ+75jWaeglSsx0wh3D+/PiFFMBnthStTz1wBjJu/AhhSf
NsJ4/CbOHfBn/PMMSyfHpuTM4y4x+6lbjGzMSIS6N0BIqp2ZAdhbP32/fsgx+PxUAgu1neqLvohb
dyYj8CCtaa5ubssBnlcKrq6P0y+0vKi060OSlEBSDhex66CWwXoT7hTgnQKJzLgjE/5Z2Ttfy1q3
qYKYNwaAiDj1rIYQzKYXlWcMbW1fG90a8+GArwUyfZw5wT7KeTTmF4I6xWsW8C1XaS2e2ZVYfQ5K
f7/zGsPABxmlSSkkS0GONMdcHFudghuFwJi3/5LxCeAHVmBNLJ9763Tlmds9SJFlUa/UCr909NCc
gnN6K8JQtu9EBiTu4qfQjVKdXO/8pYrHoVdxYStGzSf86RA19S4IndzNj++osOgqiPnMN4Fj3WJQ
Uty+lsK8hgrXhV3V1LiQEqWl/6y2QZN0n5n6XhebgcBAbHvSkVNUGnIWWo82pHjAj69mk8iG48iK
u1O0Z/s1qLAG/4qri8osCkogm/Wj8KZ4GagxnXOLKgBNTECV3/lJP5j7VTjR/LV1nhB6ESqfFnxm
neIMaBZfXEbvTBaz7cRqzflA1gcVMe1ZQYB8kq/aYBbIv0p7HYAWDZ3O5xwqD2geFoMCtypCLPw3
W+d2xArddeh6qt0HkhwickXnE1OwY/ahMMtVO0cK+/APHOWYCDlSpGlWaLIyjPhjdTcfAgjFMoAx
OODCWRNspLK8NNKXUx36UzPBtDW0KRDyrnaS4AXV2/SzxVe9S6vAihtQuVFoOoQhl8EHOmV1USk4
wyKTy9Q7EfF7+C6W15GUNUS3V0W3U9KfpYMLhOTcEOYjq/PrlI5cJk38auRFOntr8fm9iv/Iyc2x
LrSlvqrvIBxiAfoWtU40MiXMCDSDVa0fbfXQlCjJ+w9L0sUeqUgw/SWIiwO0STwwiDld82ZVf/oA
bkewQyyZ0tk5RdaAavF95Qq8ajVgK5zok3hY1hL43AZbMlhU15z52ZLG/Q5gpW98n2BEhGAEkEON
rHXz2M4gw34UoF2s6nFcsFLs2/UiwIz2ExbRmXveUrV01h/tOKXEUL/9qBGs0JxwW/QifEOR85/T
othjhUNp6QAbtEaoWhA2j90L2dbR6ORnqPsWBQX9zDiK3U2DV9ww1eCTQCDwAgCFPi9RkzuH6HTS
CQqx/FpM2XsuVuZgcYMV/9AO6GH1n+e6Uv6G3/2sS6IFArO4MPz/jDXmxkYt5eKcILdWI8ZcdLzx
KhID3u54m68AXh8O3mjJJkVCg13vUXQ+vWP6XVaXNonLu2GwM9Q443MUH9RO6oMcA+BhEtJU0Sib
XWX+p0x5MFp8Myy0ipS6bkmJn9OCpabTXbocC5HI2u304kOBtJkBJ/imTuvn/ZiK1zMNA/psvPue
oWkK5o5XRs90ejk8VzD+DuaMlmKeNOhrGeE6qbX5FMI6vnzz8F0NSeDG41GytFfLZ65NusI4mxAz
aZm1BSTRRT65UQ1UD8Zd3FLHKyjjmZEPBg2EYgHuFWwl+MtVxn2tJuXIdjsOul+h9/1ru4AqxV9v
zbiQLxmqoQt8moNeq9tQc/Z3zn2JH9r43Kw/Sd/Tn6YV03y+aFTcWSSdc9FcOsWSbxDca6a30iYQ
K72r5FVuVVui7Bh5CSNLLshA8d2/KANzzDbGMs2eYMvowHdbAVQlFFTHHJ7BzpEhA1Z0RHf+F9TZ
ItonzNcyF5xNGJvC8WyQ7GfIIsolNiBe2rxGOhzzyqkMpHYxM4qQK64h9MYLbU+2zTFrwe+DuAQG
VSj/zbFCcyGKizLZgl7opCab8Ej1pYYqbKxgacyrQacAW/Ewd63APqseWH46oLmOQ+3b/DxH5Z0J
BXlVAObZwYsg5247dF9QmZOlGtt7YBkYQYqezw5iWtR3+RlHg9Izdj+O82ACpe6Ew4w4vWvjr5Vh
VheA9Cha5sAt9fPJwH3eiC2js/vUn8NaV3iSHh4n7RydXlLW0n7YazYkwplrD4g6Mfuy+3De8AA/
Ckdrnyi27Bwn6C2oikL4AT4fTWiELlzSyBU4FpA4uwH08TK3PoYKFcBfmAKQW2XZhbzlt5uZc8vM
3Sd27l49p7ROLarcS6eHhAJY3RUTMl4yZrKh9ILDCOBe3hZ38+YCtg9RvqcDjvGTIIbxJ872iNbz
FziEyP6FQqixXuQtpP6y1zmiOXLNp7dGpfVq1pUi7Huf6EKT9yhlqS1buz7jYABT/1qpoY34FREz
/FIBBwE0WZko/1cpPQiXiGLVHquEzmr4a4Yo/eGQwH9tdMcLxxuH2WXvwQXFecJLN2kd0br8f32k
+F3RYaGDL9xySeXVcHGAyf3f3pMhR9W+z1FxhE2oa/ViyG6bj4tQAp4cT8qtOXx1H5Xu8MHW0q/N
Ku0GMweFk/dzXFlSJ1Jpvr/nRnxRgBaztN1oQnDElATVKhi7JzIlbLwXyDp+LEQecFGrJQnXWIqj
ZKudF2aah998QwTtJ2HgA14q2qnKdJEG/ZBo6QAcIcgx9/y1P8N+EDlCVp+2CrUFo18G1ip0rKC8
g4MOexV909mtzce7SU8gdtb9fvwBC6UGJUFTTQxe5ecDfYqTbKh76pL2w6/z3wYcBRNyDHzvKAnn
kRQSnGkQFn1xxN2oAi83hNwBf5NDpFHBYiTbylyyG+ofG05JqpYS211c6mXTyQVRgJQ2gO+eS/E9
0fhbq9cdMLIGG5+UfzHznjEEJDbHhT8iuk18oCDNg6yB/rW2qevFYqzbNRbitv0/MaNeUISjJU1F
dwTopBxs3BKxmTGcJoAiExUyRynXApyEPvmorOkg2I529HEMdjSBZJPLrrqAK12Qv5vIs1/giH6I
sU/y/ixxHNnozJOD8QDMAsSi9tMbhS67MO8GZVPMqTQC2qthneNrdYTC25z8Zsm8fTb1Gx8LNhQQ
V0RitKKA80zYe36wiQqNJVPiHlP5SoOPDRfv/O4/E9/afAKAOSGBYTt7wIrId1RtSTH6wcWiuNIp
kuwF/oh/Jpi5X5mJSllXVseDdOgcNPTGrpkCMOnrkIVg9da8370wLhKUq2STfGfWyOQTkrDgt+0b
s2vsv3Zt6r/mckmgnQyl5PZt3iJD3OeAapjmJ9yp+SQfqyvDsSVJONeCMvtViwuwWkV/tyly9ysJ
/3eS/SisyAHQVXxm1yTHPeTx0/Xx5jvca7fvlhPOYA4pGKwBGvqz/DdyLV9w9pXmSZt3rj9q55Zx
hA06tE/sH/2v8C7hYN4TbUGu4FYC9p3KylNnuYNL4giwQbUVURXffzwhX+tfX4BZ9tfin+lyZHH6
GTcE4pkIAG8By1v2LKNXRAWU44HoPKBK5sfvT7SeYRuT3/Hq+hUBwfw5xV95MuWugjk7sZjIOUS/
+46yT4/FxvfMV+FptKJ6sOVfzu8P7+hNeG5+VFTT2aAhrB5v+L5uRy3LbRPGddBzc7iNu7Hw1kYq
AjXp53XeCc8ZZv5xe8uHGv+UuB3u2YAXkV3u4sZfLtFwZSTYPp+FdTxpBLDh67jRzT+sQQtcdP0e
PcUNscVopyLhMyvbqbMtc/glcXv2EejFyZ6+2YR9R644pV67AufurSH19cA+2ZrAq5w7vx34q6u+
Hr1P3U55l1ySsb5W6jg4qZhVfru+Szxf1JHJaoUnHUOvncJyUz3Ir6CDgAXyLlxHL0zXR4KbulPL
CZYuNwuteWXVkDUeOdTBdpDMacRN7NK5qjyQcpCZCiGOFu3Tpi39ReJUEm5bsOq18cvoWs34VuX9
dsWtE1OF9MmzOkIONaFzmaUjG5CRR44uzvRgp0EOsk+IY2IcHL9Jp5NFEOLMeNbqtwo7eUQGt7oM
w4f9gustH8XzigijFwURY7/Ik5C0knmaEpM3OFBXzbdinAylCrirLBJmvS1vUw8PMna3y0Go7BZF
fSNVs+UegatUTliiHqWXipdDRgxHUrbeHCIQNk1mqlAMAFYBJTxuojAzIsIZxZ/pXGkK2w3UuaFI
FPOnYWixVvEdXB9DTnhza6XszOF806+hnT+1eCq+hxgRD0ODR6T3WIoF4ME3sF9ViYvyw3WgXFg4
V2S2c0e+4UOG1n6zAGwuWxRWcd4nNxLRezQTTaVUmxRVvacCrsRr6+6mdc2epxfKiyg5WBFfH60z
FzOWo/gmRjYXHxP3Chy4OPceM1lZphq2lYLfy2eo0jJ0DL00f7YGpKwlaigDvjHde3V99gNX8/Qz
HP3ghy86lL5umNPusBZzDKKwTHvVCWOU0Jt1y0cDeyEc+8plopih7AME4ebTyyr2bczoXVvfZwIX
iYsE045XcFtCXaRVzPwkAITJeKOO/AuHizdTiaNunkDfC3pxIR1V/3pvGQ5kf/pLqFRMylpupuGP
fxnIBTnfUkuKSZYu9MSjaj1Hs80R+O09ReybDF1V3XZC/2QfYI/rK3yhO4Q3tMtGXmude/enMssR
6AQcPLERa5ykLKtPI22OXkCzA9hVrW/lxgbWQhRCWzhdIcQgcVmmq5WWfaQvmhJNBPII0g/rs983
KeScEc1vS0hNoxZdPGMDM7eotNRp39N/DFgfAPNi9vzkwy+5/0mjQd4DCG/FFtCwfKV8yL7WX1uC
9yl6j6/yZzZTvZUTn1AQvohZTqvtdr5VPFgrfugSW91V7FP4wmfB1XU275NEs+pPIiie2GaN/fWv
I5EgouKp7Uxv4d7lDeAGyd1drjuvqdbJOSyr6CjJOq47WcfhLJ42tZIyEOMiMwG5lrySHsxH7EiS
YonUWnRp4aX017XyQ2TLE1IEr804AraX3mEg/w0SV+l3YAE8OpRiAbMDH2UeKf1IxDolK2zYrYIL
r6R4q0pDxkZWRPRDx/usLBQRH+XDGHPQOFzCQtGrxerA3d0F3gVg02P2JoOY6lYrm1/X41OAv6Sm
M3ZoYDZOZntmv6UxMlliw/1xgzsCR5NLWA6PKzau/ojGu86qSjlw0VAi42xEmMZXEFdWoXAuQ9LZ
54QKoObufb3dZDoKbGrH+x9+Uw2SwLH6mO5PUTF2ZF+tVlo6Oq34rFF/STZ6SPWYVKWntTF5eQWU
mdNwA5h1cmv1iHL/VVOSzcs+/lO0YSQlnPIYTTyN9ngaImzw7LYQN2CBWFgE2QCOUzXpi7ICiw0v
T4XiQsxzRc2X7RSU9Qqt5k4q3/W+eUG+oYzmduKYvEdp0mF0YrUgVUze7vj4+35Tp1piLSl9yfbs
Ob9QrIYiHAN3Xq920f0oQg9ayoAjp36MuvnHg2kxR48np7YPOJXsmfn/6fRG67mKVs71V7ni1hon
KHmfHqxtHxeM2s3unlIKzmZAM5nUMdGNkMGIXfQ983lg41OT5J30HBZWOn2xxtX3wMuUVK7MEIZP
13rwVk8mortboEA4mhg8UwfUbQSJA3ZPFso/PisXCQiBGDZ6ZsCWTiSyZwTq4oPKe7PFC45BF9iz
GwaTBiSlO4rujXgENsta+9Doky6eUoS99DhchpenpTW8rGCZY2FT4ptxXxJ52XckV/KEJjNvTr4c
7OHZD/zxMGY4glI6xl9w2WVWmZJXGlqKzAFGX4Qi1bnIJUQP7yehwPtWENyJHJaVYvEFRjEvBs8y
0yubEO5x9+fBz/p11wWKqt3Sy2JSMU3v5EhRwgBiWkLPN82/PH/PBdG5fx3kyvUoK6Z3jUtEjQaF
ibEGsOwWq8bSyMcfs+JNolwTGbE+Ur5z36mXUHxo0eHzwBrFpuE2gcbsmlALM4gy4iXHgpoqE0Mj
n8ydC/bYqrb+LZxL3nwktYwyCW6N7edCeN8gLDEP2OPQg3r/UEo4eaK7qE5zWtLvGeyh425dfRPT
RZI475anbuDI+brujecV9+8uuqgt9YbTHF5Mc3vjUgKgKXbAs+fnrDtGhIE6lw1cAxAXZJY8KCuC
gJXBfzxSeCGPkwhSs7rAWIEwxXmU4usVPR3zF4hJl6yASyhVhzlwBDedX7KKUCMsMId4dZraOO92
uvz6tzv9NWlDAbpXeMEiEt7zaK6pNPpj1xyoVFLCSeVJ0jybErE01+EJTf5IN6/0Ft8NJo76VOEa
QRqXmRfqHLS38JkPvqq/P44yOE5rYNdY7/y7HFHxw75WjzJGYC4iZTNGwtJFuQFP4HYdctXclkZG
RZ7O2oDlqmCUFEA45L87WAsBYVfdEwlIH43K+y8WZ8wAniE35LxZtcHwjGdlFW5M1eIkzWCgNTfF
Vs8ZDVoUjuadoTDprnS90DT1xxFU74V6y5Qz0JlXTeLt2UpznxfOF3bAqrwGTNn//bXYNd/D7XT3
XnvsSZf950NO3bJBgofqdfBNqvPXIY7jJZrmEI0sYqTOvWJh3ZppYR6zLK61myUTgOJbyMzrL+8R
amjWh1382lshktV9Z+TKVewofqsJYrC1WgsYWpSwVa0AGVJioA2MV+HfQSvFHngwImMKQIevGgh4
hG2sH2eUSwTnxsqGI9fAuAhiFWb/2Iz7W0fRUpHCYKM8PIiwU253+wZB9G6LktkNHDxsBSWBf5AA
+UFDvP9ibk695sR1fGzpnt7OffEv9OFfdprQfXUwzzr4PWt/ywH1bDHuWGw2Zlrdg5YgNCOXeHWd
U/spcZfPp8krOeGYqqUi7SYGaOugda8fxBv6UBnB++7g4cm7M3RPvMOHNtYrHhqdK+ALoYad1ldm
cG2TFnlLeehQKczNg9jM5AA1y9MiwDkxtK2ThWzjzygicQd+C/ymIPJsnRqHPqH1aeootGad9JLU
h6Mwh2osyvHstjWotuTuYGN3yM3cnrUEpMxbJUGyNVMt0VwV17ZBs6/HnEEfvEx/ZupO0550Kskb
OY+8OzHR405ZT7A3Tp75Am+CND/nwNbAjbByW254Cm2pYBQ8biVdJ/YTfJBnGePR8xrZ9u6XRUO8
CUXB9aQsV0SPVnGDxKCnUPgv/eCyFQmN2RR7PPlRzbnqssT/1F7n1uhZImhWp5wRk3eDls69mrM1
SKP93CDTywk9yGf0XXLKkSrvwvi/P8lNIfnzB7mAYsl7QHl5f0FbbWiVcR+Lg7vTbcBmm3JKl94V
mTTcLwXugy5EjoFBGGGijjBrWuyeu5zQP0oIACR7sYy3d9NoJAwS0JJctvzyCQ4LFG+1NRQta04Z
Ga1fXkc3oJzCayuDo/D4WHq246J4/lA+XzTnO9tUj1FshX79dNNiE7czeeNACWSG96LJ1ExJRrcE
AtLxhgncz5BZqk6CGSGPcup/jzhuBCvE4mwBxFZO8Ggb0xVb4xwj7UiTXrPy2Khx5ZjcvFUsuFH8
4V1k14Bsi3R4tAfS6KTJ9qPL3ZcCZMwhGJ5qv4iIb75W9pS3Ii4FNKTLPgPd6ZWG1RYC21nvD+1v
kOwu61HHSblXGALl2WUcjFHLetOO1dfyHShh6Zj3LySe2+yz0q2yLimhH3H5pIKwIx3tx/Ov/uzs
PxFhjM4yKhWBPh+/w8Yv/PLQp58ej2WLVWzeU1aXGOErJFNwwzyWj6f+egAexSCWxSjHb6hYxtOB
NSBh03iLPv0mf0dDDpN1Cp9I79eHjvqS2AzXUjFgqlW8joVErMmDzYvmscr0EXCE65uk7rKulENV
f0vBoTD3Awl+RwlDijYQwms/KDadhcQIfIVluutWJLMV+oi1bkLaXURQ4FR/7bPJTjbvAQrI5A0F
ScJvqeYoJroWLiDxbJYuAgdeaqFZSbmO+38yG/c3xjGZU9s7L5nGjhPaQ73yyhC+qUXaMiyUbE72
4y2cUWXoVACK/tEUXA70iQGWNrAzc0CZ+cR5h2ASMglCXHrwWOS6y6Pipw2hol4gFYW0IVLsOG/m
j3s88wvZWNzQ/e8NJ1ULfMjaw4SxZR00bEue4iz2VYT1tekIfbOiEwBzXB6K1LpMIxsE+AYzZXNu
Kj/vCM+OZVjYK4lAwqxh5z1lwKHSv3E+sRaSOmMfzoVgLbo8SByEbgF4QRjwgOF6VLZf/+hN80nb
ASWKkpwIcXT9Uc4iGJbXguBbNBFK6q7GotFUVVGIMTK8vGrJ4udety7eUHC+smZB1XgtjAeTgW3l
nT5fNvsRAczHlD/zuucp0xReqcYr/nUCcHJBLt4pwfuDwi2M10/gp+6r3NbD0/8Zm67QNJWiXiHs
YSIlYibb6UG7V0AZagfMBvF84IQSPgM05+WSWrV7k6HvfI17Ee3DyHLr5jaEo82EDHCDBv4lKBT3
s4b5POnUj8tlOHxWOs03F5k/gRq3FC2tPEAlrnPK811vN6r8OtI0tnEa3KhD36qRlEsQZNv1T7RH
ePi6sjteU5csALe3JoGj4DWSh2fgokz9zyuuhxyaaVsFxIOS1b//O91D/JNvTfoVUdMc4AteXCGI
XFBXZumG4hhfHq2XMKaXPWsmM0YxNgQkERAM+geBRgHrYBU/V03NgzmyJvzcP5MbJkwPck2qgnpl
u6d9s+SkpUI0fXRJPY5f2hvmZ/dLVLd6atKHJplnFvdtIiiuq4JTeHJfV3PeSB97pXeUZUc7uNWz
HVS3hn7MySspeQTen7IH2uLdQWsyM5IuZuelLSnvduMTUE766/7x9zxg4jU0NCc97Dwlcv4S3Gci
QeRnwIN6R3cMiEL2mrbPxpTOL4Dxs0q63Y+ILqgeHf/oB7CxHaqm5pD4h4Cz6jnEGY+TtzP2cOpV
cuEhbL+WL/cDsn9UsW+tw9kiIQxl1roHuF89cB84jdDH7rqAxEhPtr8l13HwFCL9+LbDqVzGbYwt
0l05ZdkU6Yb4+zy0GsppyEKwF/APNV/nQYF7CScXyDUgnnh3i+5sdqm7AiWCeBN8e/7IqRheo5oq
JYkZx6n7JNgw/2hLNjPje2vb7iCcO73aw+WaLhwkxctGUFC1iF3v4hU3ckVZclXTa2q0af7U9/Eo
Ejlrwqk/BGw/FX26IMvMS7PZiyPsYWFer/Z3+egVRoJUxbRBJybS+Z/Evaovljoj8y/NFk+R8WGz
DM2B7R0lVfpv8O/14upkmjoTOWYotW9Mj+RvRDMVAkipONyl+76XHil59PYJ11IauI15kX4KokAt
wtFbSaL9o21GZwu8knYElgL9bOWQXyBzu4p5EcbGSlWcenOlv9Nvang62HMbR/6y2ymrcULB5m4l
SKjcDxhHmaSh/uY9AZqj+YQg+wlfJKfCfhx8SIjeFpzoPJw/qaQHVEqYfwdhNeU7gVGIAXCs8k7n
EhvXqG6xAzPLZPSD4elT9HEEeAJzMEiQTxC+1hROQBN2WC7fhJLl9vUFZDQ9wjtYB5F2S27qUBhZ
7SFvDdrtf9Ism7ejZnL3RcuuR6TPRa7AeUCGfFatG8OQ0B6OW/0vvRX33o3aOGXr5eH5OXnL0iZa
y1zrovLPDDcVhMQU3bup6BNe+ihG6Jrd6pFjgDqB49qatJxYL7d8+II0uunRrOI7tUvEypm+i2UE
qka0xBHUPwqcfs5jACPl7ddn9RP2CUwiOZ4Dwjal9EsOWjx7xDLEVlIvSvAotvSQgGny8S82NYzC
CueJcxgMWZjFZV38XjBPzyO47tgIww/nf0ph8cLKFbh8ELEfCEudPW/M+nI1zJ44t/RMoE+ec5fE
kSukjNDSp1H2lrvllfwrQjkdCypkqkGL1qMJHxkcb8gBt9AbJ8SFyyYtfSliM8b43BPEUfdw5lMf
kVhoDoF/ojT8p3wmX3oGutRQPt57TNgY92HVkc1ZE8twj/rTJLSwtc4LSdQgng3P2SjW19guRyYf
uUXEkOFtcQO6jzcitPH/LWAupwzMs7z+pO5G1t8NIfP+da1PIvyTpFQo4y6px6hWxvT2K7BCClmI
5xUMiObL0JwNbbiWtoJzZxk5blt6zk6Oq974AjWU5udZQLGskFlZstQKCy5Z4VOmw8vjQxV/ePde
tsR7kZ9tUrehZyIhEGK0jXWt+oCNjxDNLpHA3BTc82qWQPPv+rafZ4oVo6YAQc//nYpP4ssnf0pM
IjtaPsEYLmjKjNY+oyolTGKCTkS0mNDlnFIAu5kcm97LEzh7uahCj+6fpd407+LoR1eTm2MGx8Qp
HFWsf1B85U83lj++UAe8nZM0o5xdq1QeOJNrnpu4wHeE8RtoRBng68KmELcvOBNupimV+3VvvFhV
bcABtngC4Q5Ihf9J1ZIZzbcxrduw7t01MWzRLpZAouQQJpGVVQQQgcwhi16TjL3OFC+s83lbNkNJ
hZWI+ZGBd3a0GDw/pMu+6wXeEAZe0hBgva1pNS8JtDZzTHYCBct7ShGQyq4Mdz78tOUzPrtF/eMp
uX2eVeGjydpAFD+HA+96HddgwMMG+AqNzs8A4L9H/8yEVvp/yGem9oVfuK2Tv+/b1m2iv21cY8wV
2887U+kca/IHHCPvOMe+Km5VCnGnD42YlXd3PsIcMF1kIBIKpAMc3AInir+5jh/mAxBpxkxC4ANz
YRYQFY7a2z+bxOGCcohI9rmLLnUwDfRJ/TbwktIn1Up/T6Drh3/eEr/rCDoYlvPBXqrFQ9nUlfWe
slu0saZun/lePjK5oTh5KCOB8j29LeI/EYWqCC5NtPL4JVN1QvlYIZEbSTAGOG50Grm1nyGN6271
QsAf9I7lE/8mYH3U+Lg39wLW5YzNl/BpQRGOR7BFWFTrsYMwuHIBALqigTsNmzXfy3TXvi10BnJX
xIUcuO9BO23lbefmA5hKr5l3B3B6BucjYBzc5HgEXlp6hU/7y7Di/gMhr2GTasTkdnHpxVkh82p+
APrVV4gaRfLOowp1jORpcx2uoieSTq6CurcBvBM8MauSisQoQ6FGfQz1damyLAQf4zVZ4x/Uh4LP
xtq1H3oFeVQGQ6s5Hh0EvNk5T+ftp/i1ZFjpFMi1b0TeZj37XVprjFT96FEanxufM8Ele5AgZocU
32JsTCBKWDTAcI2f43jyI1ZIwc9QWt+ieBA5o0ZBk6hbUp1d29dkKPwy2PpDWmzXdVyzJNl+Fh34
Ea92WRDBrn0Swlohq3prd3xltgmajVv9QZWMuGuEnBU8snC/h3yhRh46tWYxe8vGFe+BsNjbQM6l
pFGRx9t49/AtqEeR7/hwTTeBDT+KMe5+PSDoBo7c3LJT5vq2ryMILlZsCFZYQF9439D3YS9SuZMG
BzAhXER0ZDUrVD62KN1I5NdGp1wRRP79zkUoaE1PHCrMJ2Sjr5trh7ms/K9LACiz1hDUsuWyKCli
TpotVCqbXosaj/k7OczxFMsMp9SrNBAej5695wvFOhLBkVqfueOCwfCOiK/9INVR0B3nX8YOWAGU
3gF49arg4fRAwPxYEBGVOnvajOsEeSB7by+tGsFRsTYzeAnjf4Est/5V9Rqb4RSSF7wpOm9+XFO7
DkWG06MQcd6K8O8bfCsQ4lwtcG1yWQxRYa9thALuDXlcJKdQEk3D61Ci9rtL+81HKCPtmNcMDS2h
CjWDaQN7yLL/WCMaDelY/eWjDBaYWJtr5geKWI6V/0jdGmQZ4hS8VelxzHokk8HlnOvNX8VFVHbv
1PCmgl5pdpaAbfEffGsizqi8+HcenvM143lENVyIscf0jhyvwQ8SfRHxs8bfJy3AJvwjwpfWhzLq
NVJWai9GGYCmhMJ40v0GhjmDT8hd3TFa76XD52njFoV9jd6qkMHL2Bn5Xi4RUxebhEwk6ZdfVcMP
n5cxlYvOYro9MMni9/Cze3Q+jWcaviWO8L91ZASgSV1FNEKsyM06zfqlpyWWdeQUPy/PTC2eWTw8
9Mr0QesVJHokCFD7QzpitUY91lhAL9sbz0XD2TFntnk5OE7rdXUBmAG5Oq0h94Q891aDTEDqivRK
5tb2nNORqPJS4sR8mfjDb16EimmlasZMCbBFeHvM5uAX/+Cv0HwO0Ftx/06qiDt/vzImVn2dGC2R
oUnNp012a7N5q+c3D0pVZn5JuVj/W1gt+CcF65FeAPA2d4HD5DdjT5Bne8SAp7lFHVKCqs3Qe/22
Lqg7dSFHHpmLrBuRASg+aRAGblczZb3PBbRyMIoX7jaCeaigXPj3YD0PoErW+S2vgvImL1LGRPgO
Byttq5sR3j4FIYtsUnrVJrEngf233SIb0BxrwWwYKTsMh5dun6jCgQKKo6cGEKcRVNzvofF8Gvxo
trC1CX9xvH21DzbzHB/HZ/13d7XZZZjX5TWNbi7xx1XL/A1P353GMQAgj+7u2eTHslkBbdn7Aycv
Vfg9rVI0Hn5nGorj2TMa3uPs151ZoR2ZnsqNPei6DKIWBwArucX0tBs/ohsN6FL+j54wHd30wVb7
h/D6zhJPLOcxz/ehD/EHCtvtv0j4UAuRS1L24V/DA4H6gy+jo7diS2pvuBKvUM3zwvv3WAe35v8W
9JZf1bn8nAljNznBXekasKiE7AAJ4mVvj/SmEW2eQpOex35gnazTUW8KaTGNMJRbMrW9XBtzhwSp
bIKd6FxlWLhp0pDHshdCvGK0cSjnvcSf0z8x4VDLQZCIbloGhbF3erK/tcB+8FJeTus/h5k46jeO
o6rX/K/tfxIZW2gFt1BKpPK5Mgvt315XfrtsaIxlqQs9G2oppt+cTarTaxpUbusQL0noCuugLfqj
uneLamSwhNpKNYZagF3dCUs+GG1U783yAjgp4BnjqobywBhMNxKVb5XbH/eKGapinWj74IN4M8tz
kbggrWD8/f3ZtaR5uVxyb6S+lj11mEEokmrZq8v33ASm1OQT1ZJxjEfAsES6ouVJkYCvM34nAzp8
jovfYkgxFeUfGr5fPvjOvLGh23OE+wImr2XLANWqPAgujqtqovitbtsGbb+gChgTH3o8iAC3buqu
QZt0jhGiiHferFU/5dVfmSNwfP0fG+fLnhoX1Kaot30KbGCsuBhltxHkK377H1cyl0B+nkP8Aw3g
EoosJe9T+aSwWLLmH8Aq866kKFBnm1x+Si1bbo6Ebw5ds66H0ME3HPqjHhJL351jUGXbrxRxTtqw
QIUg/hrguTyDeaSn1lyakdB1JR23+njDYhEcNlUlGt00TN8ARzVIK3MicYuH+9iUUxcQ01BhJ2Zk
l1cieq4kqI/u4HgYQnwdsFn9ytXn5yFsvW/ojcfVh4NTzWYeXleMuTB8NLGqLtykRVh261JELu7j
aVDKZXh7caEXsedGm+pU46walaBmJYdhS/YMsfoSjXAQt+BtBYzCGSX8agxmRYK9dBrGKHgZ9nRW
VSDxitYfMFsBlPw5HA84XhsnTDnIPSNHJu+ZkcEBdK7gTl6LVEhk5DBr9+s47Xb8fPMGLS+2H41U
kU52XYX63EAqJeUyUVgIqZUWX0yRz5c3AZFVTPu6qb0vi5/M+kHSlpc5m6FtObuhMBLpi7zaiQ1x
e+rASdnwMjBYaSqLOpFz+Zyspw2GowLOpQYwxnfJVFPUGe6ViK725xA9mytZQ0EBCkdl6RT0A4iv
MZJiItT5dbBPzUZWvsJ93F301BH3lTv1/JoXmQM9CfXA8+0/byCy5mScL7ZKx+bmw3U9K4AwUfbe
FmFepret9J+Buqs8mdANPxdFTS83+yf0Sg29A66f7iEq3MD6f/ySx8ZTfFzbRddxeFJettyDE5wI
+IKwA9lDq5HgZ4BN6YTLsKOBPBvvzU0sYHBXy8epRtn7zNZtQ6OoF++ag8TUMKFaFE4huG8ngyWu
3EdTaJifH46TpIfJm+dTCB6gLspyOo7Ijh9iPTxlu96hCp7c08xVrWjrRFGZlfYSIUVm79n6p6am
REqwvHMBC1lrW0Jv7zzKsjb2c/j5d5FboTReU8y701B3vn0O4wWpCBNmA1gP/DYF0S7iuFVfSdeo
zkG5jQobMSZwp8YXQCsXLheZXwLDcHiaPYrzxzBdBRUp/FK8WXbICsXpIriPcwvJtF/nUIfTeasi
3KuHILwmZjk+hOrKK3Hkaots19W9S8KW0nySZ/hn7w9Gmp3YM7bJ+077yWQTCBKfdgo+djTPnKO6
oJn6f0LyrO0ye2BpXML8S+qYrwQf/IozP88rBMEy9c0CAQKPPHgsHc6s3zoG2TWaH9ycDF+xZ/0F
m6C65lrII+7oXctGG4CzH22HQ6nnQhHk3vbdnuXH6EPRqlH3FBGp8iaYIuORh/9oM0S6F7Yn9A9r
pk2bLA068OU2tkms2KxoUDz5DQfdQfPROClq3RW9X08+hgCrSfIfThnPJ9T7FA1w05lZmrs76q3J
tGv3LQumO/hbo+d+DBLUmOg2Z/Hj22SAJCxTtJDWxfQPM97tDzJ7thEmPFPh0dPCPcinOf8rm5/5
P84Tzdbl8vEpO9zRiEukVS8C/90M/FGEW/POT3NdWtQXDdxTncN4RWCTGbHVyNXCJ6SlCXTcT5Fl
RdZpPp0n39dc3IJu7Kq9uE4CaEjQZOk/D0fHUQu0j3ATnfwd/kVoZQnGXbk7LbCxdIMcoRrsFdPY
MBurT89yIf1i4oEgY9P/75P0EJfVAa936yhZbZB+8a5oqV7hFq7x6voiigzGq7XqiWG4nL5q1uIu
G1R62xaPOqaRzprewNpIiM+NfJ0MSgCUUtw8OYAl5J7CqLLnvJc+NZhJMygQEwO0hAtC5BmdNuA5
suYCH9WNS1Rhpi5dHXMMdDryX+tP23FMNr1AEHxHlpOF9985bAwwMqKcwe3hlOWssoPxc/ZrKczY
l2ALgDnltN5HD5bPMkaENZzmv/ATKMLO2rlS8ENAczueQXJgFsVcjV+l2Tw0sx6AusKjbw3RtEsW
cBDv/RVKIiNhPcKZSCax9egAXyMEwE02fMzaKpY4CVluRR9fYLKe8HJJVHtfOMnMM3fjJf5K/XkR
sd4Zi/5V6mnyV0e7PyuRqdBQPk6Ffn8XHIJcvEpCFXJFazhwJDPV/1dtqaoSOlgOu8/jSaSYOkCC
CJWIDNM2L8pnE85KEKqr9U1NqmmAHxfv3JUcLkFiXl0FPiGqB11DBHcnqHJB0uNHOHEOxOfttKs8
geeI92NG90A6dd5/7WPlpDFzGVgbALCGMcsvtM27i6ct/9bUFXIAF9GCdEE4eXmcluaR0oBED7T3
mQb9F25CMfyg4+2CjqsW+zOjjncW0olsvWFBMvsamql3cuIuJrGbfzz6r6LnmCN3Y2mDJIBASlhp
yYwMIpTXDy9R1N08YInXqiOCteKq1Cfn1gwGI0Vgreb7jqoPychCo6xbbWqmoka5qhQn4RqaWa36
dcJtc7ZQvpj1HNhNlGmysvpvUFrTeSCHjGZLLV3uouyja3JIG1Sc1FElEtbBX0rqKBMKy0jxeejo
6exE1lVgk+p6EyQMC6CvqfW+ORYw87cMYops5yGCY0dHdvwB1uDZ/gf6p3429OeaU8uMrJj9M4Ue
qShvF1XE6j0hhBen5ySvP8dfERiSYRPpnlSN1C+FgTSP8sU4cttOded2o3flCqyVc5xre801jYCd
VV3mYv/3kZO7vuEwSnNog0JQNGJ0borT9lTLokwdCPegWmobZi7SDmZvM6Cetcm6ZDrmRbfJ5AQR
pFfq2Nitjmzy5J+xS+IHOMtjKYHbpftcQPiHdCJWorsuZeUYZCJsFb83NzbX6U4QX7hC3yUvxi0U
yD+4zxk8J8uAB9d+/EhyQ67e+5JsK8vlJX0MGVCH6IFLDzt63StEKnsTa283eeSr643j/vAG/g/X
XzyoQY0CFmW6rvTddsUCr7AZR9/aB9GuU99wjhPnbBwO5weSeXn4D5bW6QRYAszbUBILRf7/Xrtv
e/YfiK0vepS7gpwXu5EZqHfJ0bcGI7n6b3C/8h7GptD1lepKZv5S/H2otvwPCz8gfGY4pDVOa4WB
XWQId3xLNwrtjMut9FbA4746dbrd4IZ94IcEWD3ixDpQRrgiqC3HVRtKvcyOODcTVFgRXZTo+cvq
HIki3ysn3Xu8jaooUJNDXZAgJzxWyyKgkY7dfHtLIhMt7TYtjdUcvn8fFod2whMvNEbpSQ/n83oJ
arU+fD1O6MIXNzr84t+GtUniAYM8WdZNltC9cfDaxkP5RNjiKLBNSXrLPQ9FLWU+otcrjlkiax+J
Ri7ZCPogL3IUKaZcK79kgy6kU7U0xh5LIFLxlNJeG+d/zEnCBXVtZ8lzigdRp53u3YZl9xwqe6pW
OGdcu+X10gyNU0zAzDARoAf1VJRmXZrqgBca8PepkqN9Wz5eO1hnfhtvjDfFXrd7YERKDuc5weqL
vqKxKNEwhqbAbZSVBxRxlaN6lDCvWFossY3X0dNnBNyScl9r4NdCZ5Fvyba3CEOqmM2yYKgi66L9
nzkSu6US/pa2SHXOi9BQSKhcLUIrFr3KeZG/Pzs+jQReDm7OwhRY4/LJ7lnnquPJ1fpF9j9YFsZ2
4yAM9vxNl61mv8lQ6OIBIlFfhVQvvcrqbAvrPlfPB7NIK0o7uh2Hg+9HK0H42qJAPQnngAchwYjj
rYHlgoOzqnwvg1tNVpwo/U/GE+zM+ij4ChUfe6h3bBttY1Tje/GDZ+RrDL85Ns3kBrKyG1aw+L1M
VXWPwPrZLmc+nW06SR/AvliJjkkJOduEjKHpaepb1HSMoKkCkEODdCVx/5CO1UvA6xBbYMvGo36R
orsx+XwR+Nmta6E9qGjNgUhAPxnSSZS+MY2xKg+B8/PIbzL4nptTdr2K3CmxpPoBZjImLBzxQzp1
ZH3oKzVctxqllHJORnQsN9CG/Dc71RGz8he90EgvF4SAuw+TGidpuhjDNIkqYhYaSlg2MDKoPKT7
HyH2/Y1YxakOc4lAMgEmbtLEp/bMm6zZdTZzklaM3h2EWX0EPK2Ap1h4xGkuPPWidiunEBDnvB4Q
nJU1R1QwOtnfRruYwTXxH/8w5JElOpr+xHbp429HotVryGTJ9bZaf0qyB5GNhOh1LRfcOcVfODrR
ZfddcQ/BGZB3SVf7u9zk+fe/Ffxjqc++ceLVK+uEac2JZbtZ5EYa6EYoqEWlDAsrqu+emHhUrA2l
k93t/BpOH0BFjWFI/ZLfsOdCEjKnT5DxEaFofkLgWMx46vgMfT0gY4V6VfYXM4n9yXWwJxo63Ohy
CW6OaGvFuavhTdvD8kGRYO2PIYk3+I8hNQEeOlXN9jEQYPJa6j4yVgtm06DRrS3M0yCtUauphe3O
ZLE9xTj6cwJWDZjw7p1khLUBha6xngLnSb/gkspkpMJw3qeKVhakOYjFwOiiJcLXZIV4B4OrA8+q
Zs/9LMOtEjiNRJy5msyzbMOF/U6LhKo56+UNb9qBc3M993nns3XsPSYVycLhXjgQk04am4OD7hEu
RxYy5QBS4PLjv17a9THVhv22zRivqi1NUBE4PSbgq2M7TTnS5xwJYBXrdTQO6CmvA4R20ZQG2IdN
ZaoyVQ6yBSLs94Hh4E55fvWFIcrRKlQNe63dJWkdZJu6l2tPnuSm4x/yu96sgzR65BRt2tbV9CDB
nS+F1/09JoC5a17vTsCrHiTF3ujlUHneWGxVmdrXQ+VZMtZzIasZDmxEppVDWXhezjuuEpSoPavD
QfiEYea6WUbr6Ct3I1mLxR8BxCba8GENFYR4HFfNYEQ/JJAi4CeJuKatxy0/bdBCuCThzDQmtAO6
ECd9cAJtaAlS/mIxOqcYbuUP7dFqYgHyasZRCeLRlCyqpdnNEf8Md9O/qs6bpBSX0rxEazBWSQNG
3C/Fj1P8TbBiLlMWcnygsijO62IK4g9D7P2Ino2NYQRMALa2gltGroOiTShFgv1P/D1jpfXycRnT
ReqL3GGz3cfzPpNxdE1gZd9oGeu5xk5wvKGy1/HMol43P627/BWPf0prWmQmLcm9JWpI6BLjcRYH
Xiy58qA2uvpEcBpjHyyKWdIaXTP1QN6Bn4+brHS3qJ0IyEV0DN2L+cIM5Gfm2g9pI0/7h7toF7ms
eSwv9WuGJpQDqfRi/qjQoCIrSqgWQX4ubc9mlgEdCoD+rjPM4S3WWI5O1cTZvEEDY6cpTVgjPLAy
3cSLLfsQ7AGKQ1VOYfik7xu4YRzRm8wcputlbi7sryaeQ5R9r+Bl7v7hy1rBRUwbOPZDeCwDc4ah
siwWD5NI733WVsPJ1My0cm6vNx0QuFXRzkFof+MpKsES4XLuiVgG6XCAzYvNK4dwN5lJc+VBSMyJ
JshxKaVVZRrmHY4hbSbl8JyjSPFjy7gRKaE8iS0ZDDFdS/kdX4ElV3zEMn88a633Ddujn3bXCkfM
tfxWI79OmMRn0BiySB3IkwJhs5GbJnqNJjBc0CiMbLkZBuAk5ObL1OguJHpZdzRr6l52lbZPIyX+
dba1OXMTkjNDvHKyIQQCA1oYvlqOOCqnJmknpAHdPKuaudNtBkNhp05G8wgIjJTBAsOxEAglt2uG
78wleOMoufKmJBFFGaJq08JfuVALMd32I7LPhlV9dZx/pOpR3XgLD7ILTDx7cuZ3+/ZWrR+4ccK0
pquPyCBBfX2QZrNppBbCtoBL7Nk28DSvBcd6onUbNmf5GBYDdiukEjCIype6MS1jhiJq7vMjjdCi
2mRx6vB50ap5i78MtWarsIKtla9hw+p2M6qz1Tr9rgIup0IgoOsYrzHYh+tFZJ7S+B83tfob6hT+
3dU1+fYrFajTvSM7HlU9/N3lvqCkA+NBRGLhTYoVp3zAO6erkBUZb+ylFyMQ4OzIKO1NOF5QetiC
QPBFYkQDBp3KUNczq5f3bT4NLUkmN4+g1Zb1L6EpsXjg7QMUQaoHQDryL+WNhmmMbZhzl46zkkdK
sOBBt5OdS2CmHfTJbvB71VXwxPB1PuDzo0HmWceY4esYiD1H+jdWEVwtqtAZ37kGxSocxsUj2miP
nYp7xxWKG2RzugvnaCF2rLAeNLfG/klHpQdohSiRaRExSxH55FnQMqsfSNrpoWUixpTj1hJ/rsR8
25UUM06ZjM7j3SfpXmExz8CfKDtIgua6/iFE1ORiaar6zgnrnLaX5PhiLduHZOn9JtKGFtQpLTaX
zDVU5bOjwnvZ5fJJhxCwKIsMIdPgiXPjIT1n0k0UxpK7pPOb/6MrfEbk4UC2VTxDU1XRLWxzqh2B
bweBLD33h9ihscrl6ECrPd3nB7pInOfZyKFw17PaCwM1p3S8dZNcKGSR4t6tX1FBOmyuaK/3U2FG
WNDxdhxcPNuSr4J9YYwUCWRonZA2EsGbXlvYLqM144L9ClKbjbd2BrfrkrubY5jC2/SGZXnvWRSv
3Mp38sHjxj9q+vNVji4bMvk6NTq/UjPeDyf5/BOgVmftysH4uxPGiFA6a5HKq4LJfOCDtKv580iA
l4fRqjsJfT3XttL+U1Yg6CcvXd8NlcKHfm8qgMJqeNt/I23QaibuSEehMF5+TfVguWD2wrzkvyeT
HyxcpcDM0GOduASt4QcrpuP+19wOGa8JbXb4GPVf9O6MDdxdwPt3+7ZmBLXwfXMNzVzVhQOgrCNw
ci4W1FA+MEGEiep/xfvlRRLUk2Ts9s/WX4muSs6QQ9dkaI5bt1yv7qIEpCR7PqNj6gBlyEcPvCHV
CZGdksNGpltJpOflpps9KN8ujQ2th6Z1E7BaoH68YjPR6aFqZp+/vnPMiaePkzugS29j6/uRboJN
t35Tj8wkl3uFsxYdIuNFsx0xidVW3x50YWPK274j7LM0gOck5I63cfS1UddUIct6e8O2P3dIrQVz
Fu3tc/i+yZozBlXw2FVngqofGAK5dv4Qy48qSmm8W7N6GNwOH1NPZMGNDRvWsBctQpmBD0DvWdVm
jpI3qE5/SGbxq5hUdf50RxuJb13upBhh7rSVtFehFG2f+x61ufLykmpLKl55xF3QHEM1cS8QAAXA
fifVn7ZQ0Xws+XVZHqIIrLn+nr4n9Zq1SMjJ97kWF9ljaVbt3JE57o6zZ4QsgflSAeaY1naswqUD
mBv8pvVAK4uYWPHCOdMkCbI7CR/ydCFKTDo0AD451ttu4wD/74UbRiGSAz61az8Fm4uXiwDu42Js
GmZ4P82Wjn9qUl8PSaS12VhWAQO3NFSczwzLkj94Numnmf4mPOdhxNSASJCarth3pdSL+fCkkdqf
YovlbqzVy1MhGdVJtxPsQTfHLojisvK4gN+tIYSkgCZBEw9xD1qKnng+AQbN7U88wktvECBzjZz1
cq7ow7Ooe9HJxFI18DwPkoqGqgzjJRHFUU2jAGxvf6Fo3j5IwN6UDeKfQw2jHuKdjw+VCq5aDYvG
7GSb4dJ4icdtZ7IlDrgC34vL6Fc37Nk/bkk7Xj6Vas/xWf/IE7toZMuc5k/GZKysUdATy73S7rQE
tNF+wW0SSlCq4B3vteH7UNssyMm+L3iGbgA9HgfI47o2YPpkP/GpxbEmb3asIVhxBE8HddiC7soQ
Nppum87QLnL676jlDhJu0yEd5xXeDdL0rJcWxMvGBiJrXDOMvtGbikQ8hBEHb3S8kNDJE6CmC+VF
Ob9t2epXsmPnQupEldUAIZtbsIW+Tk696cl0Tgf3ru1R6k2kCZ4K/LxmYGEtc7Hyvqj8qsRqjVz4
vRM6wQhJoXE5+y7h6tWPZ7pmfxbytuHALETFyirJQAbIA7v0/0psK98+gnZCbnxErp6hoERKmcAi
JGLn90YC4iu2Wds3ffrmZD+Zx62IxwPADQPHcD9/WWdp38tR374dzEql29IfiiI3nEw2Wcf4QNSs
PCsq7JS/Xtv4onahtP/sINpfSnDPxKCXRHYmU1LJHGYy0wRVyenSDIo7ydEkaL05BE6miMwBrGfV
ECtaXRsSMJ5UGh/xq5iqz3IJ4+0zSJ1RvQzRtTKGpoNH4CTxi2gLLYWCUfF3SdlCjlVorCRTavgt
Sc30BNgBFQphw3feQ5F3zHk4gcwAZcrEqkMl4+aZRQ2Qcb2oxEI76DMSmCmrg/kCOzC8vy61NZbJ
HutkZ7iO7caLV+9ZuiFppTxlNWNAL7HLsL5iUUzPgJyyd9PC4Crk++IHQyF1f/z702T3WfdVbttJ
cHhGt3b7OHJuekagW17bzN1aMJ1HKsx06ylo/bQuMhBPc5BJGR1JSzE3YfuF5J479+eXgh67wKFB
WMuJt+YlxVbvsnxk+iVsZdVZZkFJVLuJwsX7DAOnFLa8HBrM+lULmY13xPpoAMTk4gNND82QzClS
aJqIBrV7HzoNEpaHer/gt0+X8AtMSPX001LghIKVsWi2Zi2ndoej0kpuH1WuKhPG56zbYs19ROl6
IMyS6pUaWOiJ7pwDsKmJNFfQoSwxfQ8luJy6CANOpZehXVNuJNf+uULqCAF/gP5W/zfmQhw130QQ
s1WgG5M+EU2l4CD2YVQL88gntxqB5LI6Uq0J1M5yqaEuu6D/y03Po7xP0PYc79VsFOFmQpSAErd+
8h7icK/cAFC89r2yPN4X49pTLSRJtLpFQ1k9dhj5unytfG8R/yY+YBkD6QNYoy+Cne9PmwHdELK5
PE88dzfBQj4STZAfw7EjUQ+0o1fH9QZ4xgf0BT2XbH2cFM09bHws6cDg+ifaMHUaplpXd40AuRej
rE7J2Q6FrM5+gI9lwlBLP4oVoJcI25KgwO1hXohzqC47twOfiv5+s0oJ67mc1W8QkstwqJDaG/hL
QuXMTPaDgKCI6PG68FbBXpM9Sv8uVgMJqlmySPac3GoH5FwdqFOvwe2k93Ypu+5pbCT8Bs1Ak2aO
/NM9zN73Q6EWsswaK4bYkqF0W21V5E4XIYIiKSzIgf0edShPXHYLuyzZcg/q1qTswg1T+jwrg0YX
4XnigfyhnPQsrduC4TAnyj+XUBxwl09QJdTgNL5ZOtLAa1cfLT4tfejjoY0qHWLJr57YXZAs2QlN
62nr8N9HQaha5eL8IOdM+wkY1bMuYH1QhTKTiAkwLknyeo5Y+h9PlIYR2t/GNuL3geayu7fNdHeP
iP5yCkcDNxHPUrYRf6YmgYkv2Epy0UAYTknmWN3DvBIzmGK6Redz9PgKNGzHcd19x5c7DWh0xJII
X7pxpKxZLCgsv5QHwKDvmVgAX5ILgiMyslE3+AiCErtiEAQxtEgpZpqXPx3iA3eRgwjYhK9h/kqe
WyzhU7+ALcBsOQkqknhYrh8Mjg8yAGsqzQbKYx+jlYarfST5iCDFVv/p9Y3Zj8NuuWYpRGWwdRTj
vYgm7odqlmcgDwumaV47hEqOArRha3QxlkSwSsJPIFR7Re6qj6/bksd6ukiGCVaX08H9m4X38kb2
XbSGEa8o8IbTEvDDkgCR+9mTW29+zRA1RjJhFObWw/aGui2daGH2aLNwqhCSDsE3MNaZNST3X9rx
TDVfzyg5VUgglMcNl58qST3T1LuhMnRSCoAK6CHSeGBttQU8zbHLvhM6L8gQKD7t7SGzYHTpbzDU
0BRL3S6ch0AoxRu633Ok92fgCRMZ1TxyqGuemOjEM/a2hStVByytiRLGtBLweWPyc9TGnDlADK3K
+Fm3Urh8C9/yleeu+WTk9CSpHLk2jiWQhqW49FS+3yRDRtEwJLOAqrlcTawYY5tf2s6ie6W4BQPa
jfiNaeh/4Z85K9U2jaJaAVN2C/N+fE5sHNCxRLHIAmdNFVl6byjBAvLo+6vSqxBapjFg7K6D2U6b
NDddWPWeqT/tp80KYK7dh4qyyxByornyLLzR9m+ZkfC607/r8PZI7qKSOkcUqvsxpqZGqnGj/iQ/
bwzpSkuH2b/FzV0x075YjeqmEBHy+sSGAzqg8DSxQIsb434U7p5Jo7ASKjVza7bLALFuTvLTJ8jl
rDmMLgR665hYMGppnmFQVARmVOpkT32kt1yo63lQ5nwwVBTF1mIfUVlrSADw1aY15Lt7Jf1J9TKh
j6YPTSLV2LJOdbMR4AEgFiprXr+GXRxyamOaHvuiWiqTF24lsnWvLFGaPe/J6lo9ORou0w5U3+fu
8XXdjZa2oz5baoM7EsENTOobcM3sNf0TzfYkIBwY9GeIVp63UGnBxz4VE06S7U8FjWpWn/wr5en/
1zv/xOXl976L/v4CnO1eXX/pPGH2r2nWb+4Yzch7L4rpyWjQQEAolfvMbVe9wrIA2E5X4nuB49rB
7+Cogf/gBkx90LEH+bF/O57QxCYXSnT8Nwg/EiKA8k9HVeFJDsVCy06cegX048qiPN8W2Pnns2yh
iJdhHb2sHZogCWI6wLx08L+p9dMsnrGpG1fWyzWrxC6IvwyYrx/F1lMK6bwuGCg95n+F6WLLn1Fx
7IEZSG6V23Eau0jpUHurqFOG9BO6xfug5ixRza4du96M1+LQKh24+i3OWEDGMTsbXuHgZgXaStGy
1NlpRJdXVoJb9gBD1Y+dOycHWzAY8hjm3jwVPY+oC7A++xgFptmCWeaN9d25AoVqqUjuUCI/x6xo
pC5AvSsqU6nwC+1ljcXMtg+gmgs0r1xUCbKltmTwMMKE1fh6x9LFnKeD3zlTz1GEe/atC3Jnh1xJ
aU57ogpMOjn8jnzl89ZSrLMIVNzSIPYuhE07GzCrLXggP5ptPj7FhTjcaFjnF9EqAUqHz17hDknd
24TAO8dA3PCJlV/jWkAKI55asJ/rqcdf9K0OuqwaGjiAXLTbg7nrpcAzKeG0NaikPxGkgfa3635i
UeQb6QkiCTpjwXWP4NsXzu9norCQXVkbb/OuNaVym1nXMpDqTnMO7Anj2FJW3gpylTb6dYuo91nh
j6L7sgdF2wcn1neHG3qW6bxO1zX5n99AJy7HefaWxYC0D3DHW1NPk244KBnO8JFbnGfCJ14shRIu
e0RpL0oXH1nWbORDH3NZ29OUJoUXQUzzpMC5e0vT3cYisiwmJ4LUfSsLs3217flRfxMahuXbUc4x
nC7nHtWBa6tTG9eoIw+swZ0A6oy3q9OUi4/rolDj02mhlLAJekB7rGhh/PXjaPKlc88RNl+vfmLJ
sSpMDzLQvr5w50U3m2PgI1f0ty6lbOgLhltvTTdTXGGTJ7vm304NhXhZ+GqJpaa4XtUzVBncqJq/
stBTSLYdfPR1ByDnrnp+NErhesZQRM5l6NcK7tqeTMSnd1e33JjQ/L9rJvcOPKyG9jdwA2sO6g9E
bxvj5jVpMZCWQoSHg2agvPLZZ1HWXH6T4ygbK6VGxtsDBtECAXdVQ8zl1zE5kARvVY/vJytOnNkK
f3x5Z42J/UV77gMOR+h9eWdxoUvvWC0anHTa7k0UeuggxFbMsJEs0WGyvShSDJ020+fPnLnk3qku
KlrCIb4kfBTSigcNJv1pUbIkv5vMGdmgmtBbkO/QoPV0V7qlSC56K3IG6Aq6DGYfpm52ebsxGUIG
xUXD0CO+7wCJT2DLWNsih3RBSJ8fve/v+0K/2kFQqcQpK3zuXPuTSRzfT+3HW+AaOudZS24w2f4y
fJMlSmQnnJqQZrOiOSTJMsqcAIOzGZxIl3oHkOQEOwhSpniurra5UKfcDJwuq3H7XX+UMoKV/yOY
VNuuPDlRgDlsH88oJKkY5tJrup52g7CQi0ggtuS9r3cGiUUJe/MoZY/bKDRBcXux1QqrJOGlB3Qb
FZcpu06+3hmH762yMIaMlZB1+eGRUz7sngCN3X3XRV1l2540zhVRvz3JCuD/fVDCyXVrU7mcJGRR
o6E7JBxQ26IlDWLWjg2PpO5qdanJmbh5oTuqkJsG0wV2hCjqB9jf5L+BZcEB8pcwiR0U9aW4TUq6
Jp2F1SJ4xO+8mKpEIhhZwrELyuwXl31Tz2iTtLYAybV7ULZkOD9iGOZbdeIAsn+xNqsVZE7mwafN
HzvaIREJ6FukHQD3M8Rp0vWC3ZVu0/9pfTbL9VDtcEL/1+XwmGbW5RIPBt0FC8RXw9vmbTjHXWX0
Pq+f+lbHAkxXXYGEx0dmdBb2afFBwvGOMzG549nuaKQWnI8A3T/Z2ebB1P0RBOjF194Huq2sIbV/
rGfk7CqPXAkpVqklHzoNrrWTehXr8XjTEtDIu9FLCemR+wcDvZmTF0/zpdpBCn0yZkTXYH0Si3aE
nMp2IZpuhkvjaalKhsc5HucD64xBadAgT/vB0uP9dAz4yIAsgsPgLYidIhHreLmkeGniucb9ihEe
aWjOv1Ny3Q0mU2YunXKk6XWSgW28dtx6Zk6XeQ55Quxdq4Y5Pf9D+BEDxzJ0j1DdfeKkQjx1qtB0
PasDbPIauIauZ877jH3JhGvcVbmffnHBd5kGozruMUFH0U6wvE6gjdH5ZnhSJDsj4TW30lAMIqbi
BonAqFJ4SQv0egOI3TBrRDTLJ2U0kVB534WNdci21s38+cSEp1gIp4VLXquaLcSeVbnXmDTck+os
wxUMr4t7Ybwq5CXqqDla12WH1PQEfmAsQO2PE+Rhr8nxYazfvb/2yOUC3/rwVIgo5F7ia2a3+Yzm
XHLMMWlTzWuO3UKqLSpJukC1cVoC0bODLXBogNcwlx1/PdYUB0x/phrvXUlv3A+/nwOqQvdNOQvj
MIL+pXyjGBQnnRcvp9+H0wrEEQ2S6JHmxeKjiZdcCHssrdJEN7nDw2auSazwGmOSIfN01YJoHuxv
9463juM8vXWym6wLsctOAm612XvWEHeyRCRnlSIL4gfr9xWyOv2q9lh7enKK+xxJBjVADHH968Z5
5C7FQmuSVhbIa2qWi5piISz0cHRCRwsT5kyOdYLzFav3zWTBDBT2AGjb7MuBrCrRn6pfmEmw4D/Y
xycP6K47RhIuTpIGyef6Fkdd5rxLLSwvTQmxFSkc/iatXppnByvaDdDeEdSWHqQcUtFf5JkI40TE
3pGCCvPJX4KoAHI36u5ppMKxqXiBNrwoygQU9VY0o0JONEexsP1wjhs4T9ptLk2q2ngdXGcmezXI
mTf4tX2NRv4DI5WYLLNgaD4ts+v3zpreULjcCutYTPs9ahaFJXNWtVVAER6CR7S2lrXnbL20/dJA
jjPHZNbet17Mr7GR0xTsd7+VQFRyWN8GxUKN/8lOaQEuzfWB6JF33ozMu+oSNdKxMxcooZMbdu1Q
HB9JMmYyWuqpqmXS1s4Q4zK2p9Qd/I/pBn9RzREOcS1cST4IdqZcsDHL9+nBl6by/hT69WYpRtMO
pv1V6YKkVd0jz359vyXEVd8Z73R8EnAHokjz3smyzluTANGdMTon/mATAmrwbLYyILdwq7ttVisG
02oXjd5A5bKAxmDw/GkbKZOetxqghRjr2PZz1hzBikpi2ywZ/uAHxEbJpKXx35+UuR+q3xWvI3MS
Pi0ulCjmxINklrk8tGouFSpE8hww1KXYp62W+KdH61hpVC45ENiHOY+SyTSoAwGO9mbpSX7PqYyd
cXyBz0JStqoKwIMWNbnVSRysouyTwuFEw364mSg1UQ2vek0oQnXF3BN/KUw2VVPG5LHwHTY9bA3L
a+p17PY1nT7huuLMKEoZFfuGnMY3ri5Em7dnMGyuevg6JY5leXXnq3bBqxaCFeEi8jdb0lQV/1K9
1PCyluRWe3kI5ss1+UrDJz377sY4enqESi+qwosbeYj0GDV7CjNc3yQAkG1VDejV5/Ujzm6jQY2S
+0pGvc9XDTyqKhnu3UuCndB4JoyiD44AH8Qg1hztE9AURIGdajeeH6KPAxFGSn2wcVEda0cxPVz5
Wocp53xur+S0XKgyCZ1+lqpLNnu2Gq2MXTRWTr5jICnFIhv+RewtfU5U27K89WGv0W2m6bpvJkBF
K19ZON1KAL09yu6eJPpos57VlVnLP4MZV8zRHiLxiwwkY5rCZLeKBKKaoOV/4rqzvQ84U/vZjQR+
7sga3AM4ugoGid79HxQvxDZncsgM2IXO/C27ckYekn1VkJhqlcwrlL1tGSnIRD+7svfx3e0QShYG
ndD/VHoQDUOjru2/3BkblhMW9J4VxOEbkEi/eCVV0JmcJutp67YPCIrKZoTKgUXlmN/I6cVFt5+5
aUIW1PqjOX36mNF59g26QmhuCZyMhWsowPYfiHMiF+Y3Pdk1eNeZ1wEX6NPHOIOOPxKGV4cv68Rh
+lsNi/ii6cbQbAajB+jkyYEOa5MKl0Pz1galPeM8usYzd8u3LyhFHnKgMcpDx2xYiYlDkBJasUss
ARXJTdatgUV7YHPRO85MvCExOwl+vpv7ruDaLYL92skPL+flEBYuFeZldqdhFjWwoJNYO8FehnzE
1KP6gJnwZpAx+AhHJSHp5omGWk9jXz9se9SBFE4jFiVT87ccH3NCvW/9SYq4zsw6rRuKb58IFkgZ
sfOBekupi7kwwSGtBkv9YH8wmq65ZYUDo4oglE+OQKY6Iv2GmbO22WXnYXfbTPU3u5HA+HZUrd/C
dr/K7u7zOQkIGmj+u/t4QynVVNO8If2wiP4SkelvyXjtqy57L0mYclAogO2EhQOIYs2cANcGdRna
y3YBCKKVDJuWBXXPPVsH8jXnIw5Eylmvg6EKWTHmKDRZV4L0rqVnHN2myRsgzKSUfLcB5YWGOg3x
6M/7tSLBGHaq4iaI0/eNI85oSR4yCzbnUlRvjAmsAtCwCLxmrjuQOHff20SdyijQBFnbw8+hN2Y3
qb1Oug06hEj6OeLfxyPZnlrgmvRMhE0kGPl67jnF6ssr5sRwYmyWliXY1GvQTiHCqDxIVg0hYPt/
z88oitHUz3aA4ynMo1TPumpOrqPM2XUEIshOEEp9DriWBerppeh4ERlU5QR/1ZVuT8fmfTXjDa4s
HM+wpEmUaV3lbBmRMkArkuLPRzW/7lpFaBVvX2jJvgwS3m8JmGGahW/miGSwOiiBD4uali4ufgk6
RroYOYzY7thtOU3dOLzZ6JS866eVz2zAlH6g0DMz1xJi7kRGdu+G6w1g0uzos6WoA6K/b0zWkzP8
VuL0aOkrecvHl6le3KqYPhHDzlg3BA0WC3ncx7M6WISSHCoueMdIsiOMt1fJaQZdoBg4hWPbN4yl
mLf2TBsRkpleD4FEVbh730FVArXmzkNr1WOw/vLmssBfJRAYJ8EQEdPy4j4IhX1Ljr8Tj3RjH84y
kjgc3IV7q8lQKcXKg/OB/Txs7e7oWKLLcTCZUEnRCetyRCGleaTblA1HnSH31vFcbhKHtRRVPoUk
gvh9dDM8D7VI+clLWvDIMORiHmL9tGZbwx2uvGvCCrZW1TEwT5mpV5pZmLXZbqhCnAi6xoY76PNz
L+WZ6T7ntnLRuUhxPNI2zqxatUf1ArCRe0U3KWZvWwqMlMGMnFkvNb3YT7Prp1rm74faED1yCEdt
DN1Zvb61k/Wt/H5ZaVE6w0jrAVxF4et1hm1EUq6LQ/y792x0GINqEq7N2f9XHtQqRzGGnTIEvXzV
EubBzR1CHxFPC0dMDkxOGOhteFxJFYLsnBfP3oDQaFV7xk2M89J2hbSfK6nA74mURq4cDvLZbtFk
ceVZxCZ0eKyJZ28om4rPbgzqnocyuQZM0ghU6jJcvgcKWxskgbPJrV8jEuItpYDoi+7aMaxugFxK
5Fm5XxRmbIt2pKFJlrgChp5+R1fcCoJWdAj+OpKbRMb+w+3ph7GkSAswQeODCTY0NlLF2wstlR6V
FDpVA4wu0K2oz5DHKGTrfRLrK8Vt+Xn3S5wjm8ba43fOdYcs6BTtaqUAVmX++8XTT2TKP7u44aUx
nKmVw5p1F2g31mSisHCmJOJi5RmxAPZ4ho/AxyfA6iUs1GKgAi+PPbACGrYx53CC/aIs1eDC9KkS
W7C2/b+WH/v1mZSM4/7HZMYt26TBLI3HvnGb4w3/L7az97V77lDw52fII6TrUPga/UlX5GyrVsH4
ntEKOIj7T5KcMvBmjfZOiumzoJnAIc4GkS+VH6vHUoO0bGyFm6kDZd5MVi5BSylTQ2iq7MlTwyOY
vR0I/66CHp+hBanFQeEGskNFTyRhGvGQebKBk4K3gRDQD7iirMFoAFqZTjlHal0jnt0MNKtFef0A
5ILzmXWbw86X6zOK0vxJV1sWB9+ZZEDJcrx58FyWGrk05xY+1k56jPxsCahH6P+2f0hgVBiffhA3
XnocHkm2xv2BjgNL+sbgQ/bQWJa8LgQiU3gbjxmx/zjgl6YmYx0p9hHXDkWs5pKCgEnZ9FTUGkBh
1vHOewtnSong1XvdjPQ3BQG5fj0JEWUinC3oCvQZOM7vym58raoBZhmU94EBqs9i/D+arbKa8fpo
FTSmVtRfFzWDM5mW5i62sllGxVcxqWYDLnqjyPcE7wNSEU9FdEeWsmOwihSxDYobeU9XjvZ7gQjQ
q5zwcmdC67/ScGnQTi35GJRQBrsrc/ExwcxbUec4G96FzMBLNyO1IejRoKdcXV0uqkAgk9BhKJ15
iWnFC6zTZY9rz+rDy1JK/8tUx9AQDUTtOihabAs2UEasYoWZNCXGxlQrPBvvKAD6I9jGSF3kxYu2
3ec47DMUuCWNyZLjmWJUJOG56jv0EInchqKjxgQ0ZLydBnS1+qcPvuSd/VC2K+4QsxMszx38pwyK
LQsU6Hcy07mnz1fwJPpKEqCAQ1bqI1Jbs3aOjNPrvNB5uvqpUbpjaSLLEfXOkS/do/gCMtKqlaJX
agIJ6fE9AOydcRHfUhyyyL3b7YQ8u76qOqvda4InUlb7NChPknpj5KUOdaCqk/yfnsJBOCqJmIJv
cFEgwvi7yh/LHpHKxV8+1N6OjoOGNAQKCiI2MPlhVlM2J6p1WhVEee/M3xDozAcU/pnQH+stc9Xz
dlUmNVaPyST2xqVv2cRho7oUBZ0DWoXXZXYMOZMg5NR1oub/Xg4+W1WNrfvPJzfIJL3HWI9imm5m
J+n1J0pf0ieTdsI11psqWsKTBWG384Ai4bwoEC6lXOv5xaEGgtFDKcCmqzYkLChsLBJDTc1Cdy4C
HKeMMRghuhMjTtgXMGRv/VhWbgCcIGUzJfNRy4pTf6S0gaycCfay6iEIgtRmuDND4aOyWAmhTHC0
FzQZ99qau+sC9MiKNN35eXGMfZ05slsZqBzEr3/+ncQAFRd1OsBelUdx9PGb5tSuS4uOl2bVzSi6
F1o/4gHgSF+jp574d6GPzemGYV3VtThPnYBv9ua+4/M1LMY/Ul9Z8SvSVpjszBFF76YAb+yx/ErM
89EHc5i7xxMHyDbotgRZM+lG9denGhqWd8pUn3NykKafv+6+Q/A7zGSJH6+G1GmBgYugZJBhQBKf
enNeEohKO9KRA2Q4gIZyhXDrQjYRvxAp43rCcRcOK8XahBGrOZ+5LHMec0SVp5r/nhDWyVHGrAiO
/pkT8llLcH0xB+uIgmRjNWnysJZWm/g+Wg0uTZjOSJeOO87zRf4g2gxjM1zRqgehKd2Kmpt4Kfjy
ngLL22ZHe1zdGCCNe96FsvuugqNLCGHrmDW3XvhHmxGtNzpyFZIi4bKTx21dq6tIF/QqQtkQhJdD
LyieZ2399wLNqUdBXizQrO/JU7ebUA8pn5VwcUEGle3AWdYfBbpkMg5zZ1DSgomZW3zrXfKdHesY
KSLd79klvE0v7iqmYHuHB61QC8TMMS52lbjF7v7BecbhR0eh47eCrtMe4bD2kBOck4Ho+651sBA8
6TM3WW44VzMC5BMEUE0uDrOcCQ12Wd5sgxNZQGJbqguh/TeEvH2z4WlTnQcS7IuWFIzI7oyxzUHm
ySwQytd/iCYv/HO86ehTonnDfkDBkbPDeen7rWp544MXM9w+79H4GnWrxgiR7u4AM3mGS9Hy9krZ
+MFhqPjECw+6ns1Bziq7wHFc7/LqzviZr4ADty7zyih3dILspAFf6w9Yucp7jrMfOo87u42B9nXE
77e5Y+AZEv9085tJDHB8Zu+XYU6hRkG73eFy4U8NKny+tLYSGxisehuaFruMa01aA+Gakfp9OUax
kOWUttyJXsyUZ0ummLsHCNDLaomXyoCU3EexgwQLidkuygNkePArtmdfiw2PmpCsW/lPRTUwmZAc
Am+Io7XRY5KAjBcthnCxCvilNN9ilDr2Dy1QEEsFLz0sbXYABMhyW20SmTorvBf26PmnWmAv+XIK
WFRs9fFbLq965t0wUJrrW42SeEH/n79/OnQXqMWFnb1iRNgWb3Q1K7JFPqkMFncbl9BMlj/E54Wf
iN6X390z48x2a7wi0f+7bQUpZSczDzF+peSGN0AU2D7kUXQROjIMPXVIqxB/RukTQ9JlQSiNslHE
C/nJ/LZEUToreStTpLJ57BVIFks20IPjqKR5WV4S4nZdxQ1JA/qfXhJ13Ty9MBPVjvy7tyobbR9p
kEtbDefhBBc5KbF45y0PgSpQ5L3rIJTDj7iNNkIeVnxsNGAJ1rskR17G0zrwL4FBUvNKYxlvrYj6
8NSX9xO8DWOK8TeguMAblS3ENrWHJzc43SsNBE4BaNGuaCGfauQLwCF0XH9fchrGKrnYpQwgzN3P
Knk55B+2eppd6nuwxizYLE5bKuFVJhNqpihdyyu9GSBJ4SFgb3AM/BStv+CBLTLulNoEiGQBMZBp
QiRwM99bz2qeK1/Y5eJdPP9PSX9ZWX3Ez9JKKG0R5Tle3qFdzR+tCWnOradmQogwQyKp9bf/4Vvr
PJzQabLPmdRuAFKgp0ffoG6CIhAvWFeV37QWmTw2yLQGckVGWoUZIQ05AmPBt3xI4lcWu/Q2ZVO2
71If37rGTgSXWMohI+XEM3gLFbKxu8ls2DXvCR4ZCy5j0Yr8RhOyqeYG4j0qJGx39nA7NYqZzUno
bOFhltW2Qh0C/53hg/XzDmqDKwIdGz8CIkPzg9lRaTdV0YLHb0U0qvBtKtFz/Wx21su9zSCFMueN
yej0JGVRHCyItfDhQ02K1DxNo5Va31z5BNyZb0091FTCgs/qZqtWddEpXyFIlDgmysLvH9qmtLj6
NIRmM6fOSKV1o5IS1nkof6mX25Q+HGq/N7/ABuS5Zs+qS+2srSl+MP+sgfvE0boginCmeJI9K3nn
qOq25Vc+1SPsOOieUKLtq1HKrVdtrwHSl2AOe/lHk3jJs7dp7ce6OKQyMFPmO90KbxqPbjADEmZo
aHOdO7iEuLi18V5Acd9xQbtWzYThpkjMOMOn+gXHRI03Jl3uponZR0pqLpcyvQTXJKgYnSlCQZ08
5Vg6ku1VmblFnRkMwcHcLOrN5jzrfHD99eRkdsVqLfnKsPtcavULJfbU+pxiyEtkH9WWWW8INmFW
+EvTb/SgMTAGp3XpTgkMNfWbRhgGU/f2CzbwtviFZq5Mo4vbAwzwdR5rWRsuS6zZah0/YLCU3+1d
LVdfgp2NcRF15C9o/TEyVrYtuVXU9QCCbDy5Wi5xn/620/jnQLmHtkUR76X4trwXBXCgWUqer4X1
lkCxvsL54UM/DGKEkW6L0rbHftZEiMsqrmw41InuZBSSCigJV/ELTrz2K06V90AC/mbWPy2n0k+z
X1GlVSBdVMrm0wuDYSoyRJaRO+IMKmus4tUAVFPXV5L74CPbaK1nal5mpBvGOnClY5FTQNaF8gaG
sQOxYvf9G5Ecb/jPhtKu6Z0Seg+R2RAVbLiBCGzTl6HYZM98PciGvoGKM6YyxRADK7TZwmi5bv1+
fIs7AmPvWvP8scO0OG2paLbaMHSsI7FhlXroDKaJGUdAvQBJ+Wz1adCKh4qyfRCu45Ei4mezBzcS
r+7n7GPO3uVOcr8YFdqXvlqOok5MglkVjwnb1HG6knYZlufO7mdKzhFwqs/jZoGQWpqSKUparj+R
QNAXf1F7p52qzny0xXcQItgFc3aJzc7FDfsWrWz8LVwoO2+dRQziHFVo3WOuejXWdM0/9enrXHwW
cbVFhcG8K+Xs4GSZiSbura6vp/wPeQfZNViXx2Z1rLTBx0wumfdJaTe1tG0uuhyEwXIdHoXomCch
9W0Zj8cr70f4hj0FhlCWixUDjbe6ahvvCoJQK2MBXoTO5RHBweMXY6Pu2kQbtmVolemOtMuGN3Y9
KHNLhZ8J+mp6wQuULRI1n6qeON7N9hvYVpNjEB0azPV73/ypgryCBQtn2Ev5GCQ0qwS2LczRz+Mx
UXwvT/9sDCpaRJu3Uj6llrM/ki3SS7Pn3jsecgNkO1cFK56ZuQYOKk1ryYvnDYQqmG2odkS0IDyo
puxFVwWxvnimEBKddmhZ9bOjes1SYaxPa22RbiBjQD5f230iGrJ1ICT1qHxx4CNhYaTww8Kbd4eC
8utVGExArCLf5eRaVxNBteXOe++vNAMEMwcawuN0ARia2Cpc58FmwPwyfg2ZoEd38KY5HL5ZVWfN
BXbEO/V112mAEJqYvN1XzsaU7oRg2X8j/TXtUe9y1wg5jHeVqpsGTABMD76z3E2S1jc5Yc3GNDtn
27KL3zWNRHZhM7irmOQNO2vrAs8qr0SZzCfP4OIT//Y1M2MKcP+vuX+VjThbo2DAWZx5SYlWRTqC
8wFEC8eKukxoHXZlV6dmXPSD6K0L16WF2n1cradD2B2/XTblYZe0aMrIAIZ6km+8F+rZIDH3qLyl
Fmr2Z0Nn7k4aTitCbPHbWgsSwCpnHZ390KntMrMsbVnA5F6XJ57A0CXB1xAWKLxip6cb4y/RL1mk
FKl0665q3yERy1Rmck8Qkw2iY74WuQl3kLa6FDMzWnAwAlHQADnLGy8jjRPFHm/n6ddJvwX8stGt
NVamIHbp8+Toh29YlojVhmvydBF/qjvYBS5uOu1OxJ/It31MykHdSEr8738YVoc2s2sxq5/ZttZO
+17GaG8kr7hj4b7O0Lvn7ad1jj/Gvn09LIABef43sL0tvC2H6wqA79NohacFHMLSSjc+kNIGwN4O
ClSboq5+vYXApCg8p5CbQWTBdy9qYzSYVIh5I11hWu1FxeS6xbCtA/SgvbrmQaK2XFJeQX6epLNr
xRVjQX+XGdY3dz1OT5S6RrV5t1zQIJDP38eHiIVo90sPpu36+IGse7tXWZ7FbmZCouqwOPXOHw/W
G3pUJtk5VFAjj2kjF0GOR7qUjGCOiXsNxVacTxvMxW/V4vcTrOFrdHaNMTZmuofyb9uOj6g2feI1
zseGHyzAFKg8bQU1YxkVHm5w3C9PdO11S29irT9VxbfGtRS/inIVEDsXFCfKykp4TU3fymozHaKD
19Q7cT/6XXLL2hXMzoCGsHKgXGC6AXJcVlJzoTIgEv+waM8qdA2F5dphvqHq39To2zPr8J3KjN4A
v/BInVt3Y/3bB9QdrAHs1yBUJBiwqjlomGJON5VaDLNoYy1eFnZgx8f9UTkUMLjEEgZWIkuIct/S
SELMaWaB58hJdDOoMb86+jQ5IP+ckkP8xemZAo4fRDUv9TG1IW5g46HPrTkYkODNGHaw6hzhZDBT
BUOaqkQr2QMsXQE+52lhbpJJxk2dbWcexxij6Jhfit8QViFprMqptM8E5KUWPrGspQHWGSNVN86S
NNqw6B2hRYBnh+xrCXdsphzEBgv5tX82QitLV55eDzI3IVONhXBxEa/ExMim2jXzUJIx0G6N/+zo
vgh/H9zDIfBpysATjMC6nTXZL98BAgtY9IKVb5czk/Qf1yrX97qI5K4i2RzNgmmWfJaVY6DMq147
/0U1SDoWo8EVQNE3QYDKVMUCzNwp8h74l/5EaMPP2v7iMzNdg1uVtQP3k11B7NaNlgfDtzaU+697
4rRDUd4JCYyAtowC+akbxHPZptdFPRAH1xmRMlI0iW9tYkAQyfDlMhjmqzZxsl/2QUUvp8qAIfpQ
GBsLsS8tpBQSoT/d8emXALvJgYb0yAeiXCjyg5QyWUVt+B3w4mMTtEsp3BgskvC5OO2YPj3St7ls
kUB6YWo0z5oKUfMSh5+PBRa82Q6nY05iudBYhtv4JLAOMdxpLHACCLR+nZNMaHLmTXyVe7968mmi
R6dkmwMJMX2uUXg5QMX+6FVbjSeMES8IC3AdYIsltvVrBj8eps7WodQ5SzV3jgdWBTmFZaE7NTUf
MZP9eDitl7JDmnSLcVCLRu5cJ9hmkN+aIrInIDYg7WfNpOfdy2u2s6uyPlP+zTkJuK5aZE5AQyFc
kTxmKSMyX5c8sIbfg2BOGHZRDv3N8EKGi9GCedBdiQQ0V19aPF54HFcElrg7AodxnH3WGwoSLmIf
evi6MozSTCgtE5YYFWgjEliAnDbUw0qLfO77RE3tweKVZU4OSOS79FLia0XTh7wYV9iVsnkvvYPv
VL2ggIiyCs4arfsxMi1b85g76L5v0/afmoBnOqhHPTSttb348cEx+8A2DMClTy7h1CC35h7EN4Ww
NWuaC28cSCcLBdVBc/WerR5Gq1YTJBgM4e4mQc/bPDHWBiaa10EWy6wbn7h23Y77mNNTyh0o+p2Q
NP/Y6dGFqAB9GrtZBwjjuAJvxrRJpj84luzV+m2jvtEssvNqutbGzFewp37QDnV/AyTa5Aj/IFTb
2jG6bDR1/It4oHBTkcjYuwAJx5+7+fdGwXXRoUumAn8voEol6gDy8ls+6tzYV/FzItfq6uXV61/+
dlce+wHWEH7PvLg7JOJ7N7IPbqkAKxodi5hovqSlZG1mTPOg9jlvtbfzbyydLGkcTM4osIP3HZKN
5IFUBqG50E6Pe37962fLRBYrLzcj3xrQQD63AVYWMCbetaTXWxqkQPEcVuA3eSJEWaZXHR2sB/FD
iyJHZj1AkgCOMfbdwnViakMFgBreFM9miDC8JFbOH6kIdrl9Dl/lPwrVTtj2GGG/eHkeDqC7CnYP
O8+56k0DmUpxSWz+SlP4YRaSIBB+0sIsQJ+P0opMWdZor4VET1H7K9FltmPinu4GyfmlrATJOd0j
9YVwvK+EsQDtV2bmG6Fcel5WgYFye6r9cKr7qQzivsNhcC0H7SPLJE4VB8V+vEGp4/cr7z0YYs1n
OC6MhRZjFqUJIbZ6U7d6YPGqIAN6taQKIiBRNlaJDPLNjzyoqUpGiw6aCbPjAaM+EQx6pMy3vBLo
XS8TKeJyVMH0DkypNouhwFuDJjKLoVT0NCKsJGdq2MzlWZGzm9rQcYMPyJXFH6duwq2bVkEsMVsP
Qj2BJyiFdJv66dpnpAICOhgl8JNMGGFYcMfrZfjgmQn8v/c4twSBTDHCHeu8G4xLXXipWIpfQDvi
QF9S1t+wwfVZSGFDt2Ja0ZbvHuoVix1G50sK4tKiPVXfCNoD8Q16OWqjWrtpO9pM599smOCg+3q/
s7Yj3IDHSH9QTQdoBrfUeahFs25MzY0BwQK/dcqYqFJs3lwEz3FQS7Ibi81Tg8asc91hKfn7ELX4
dv/YaIT+Tr81QYNIoJV+fZ/VU8yD1ijA81naf6bZsE5yzIDbgIaU0kWD8pOi8FZjG0nIsl4/EVuQ
Uky0oVCwvw1bYeYfHMFuTIe1PVBlcBB8gN6LTQZ9FpnPGHVKpoxaH5kMMpEUI5Y4XAUWbjJoXbkC
JnKCNM6pPisv+pZfLXj06vxQCPkcLnPmuDKeWQyZr4pfQncXSWegLpejY0SF1137lgh9slRxVGkZ
24M4+FFueBk/TJfBsO0r7LCAdlqQ1ms40W8/UxwJTrxu3ZeYf0iNSlpn4cYqFffB3BzSPYuNjIuj
8dqZbDJi9kUsT3fdYX0+WKVSw+UOyciBnWaNIFExP7sEekCToRVuPt6jYvX1rDPWJRYCOKRvNVUO
3Gc1dQeMMkhKte9DDpVL8K2ZJ0iTSUFQheaFmSMIgoU3o0fyKy1v5+QW+9id0RlSj6XYM3tCsciD
2QCvp/nx+x/D+2aI+2vRRh39PGuRW8QG15kfhw/cC8kuKiZnVdUdKoKTjaJCt0YZgT6THOnnWS7K
okkNHJBmyHj1B/Ej44FEFbN/POAkpiBp05K0UBv0BbyX7e9+JSgOE09dD5uFLjOgAuNgpyNKWIoO
MKHtjGXlVW2s4NgbZHIgSaENNRK7okgSm65V3wyXaLvyUpkdb+L7MO2kZSE2x4fK1zX1LFhbUoLo
ffpexxwOU5oP0c2RWk/PnrSQR8bSMuVui7L9GyyMB0MXdkEMztATFkcbDIA7xYUotV+vxIts6iJO
sF0qg7IKjEwxCYx1kQVcTXQi8NLpUNF8YWdapWFwdue9IdUfKfb5zuVuK67uAcINyIlojpCaaDDk
aFOxIplpO4eT0N1z2wLUChVVBDHOibvkysvIz49EmEuz8bNyxk4LJEK4Z59iEeDa5pCzZwrUBk1s
92a8j0sbPtpvV7gYOxN5x9L4nUg1WeQc47/8QDKLSagsl+hjrR/WIBH5WcjFPn51FLukXHcHeupv
Hedb1SsgxUUZquTI2FdSpq7MOcKRbEA8M0KEz6RSPzvI4gAkEOKAWfwHSJHnEF9vJU34RXFWXcLz
G6s0thT5SzqR5AFx5K1DAngCaG4gQAEsNGXLMcDxZu2AQoSb8QFs5S7twwwCdTdOu+KzRB+kAcmE
/aOLbWLdrXpvdUdTPGzo6LYjqsHQkFmUQk5+cYW/3nR20q779/7uM85m4G2qjddxKrooy3hb5sfu
G/X0iRf977P6rx5llEdxOY28S+Vw8BFKXuIHopOX1GAEhl1WaouGJDNEOTb6NQJTUz+Sk5ey3oCT
h1Vr/V8b41AqwIpzrABgAe5Q18xMHqortEMX8n58/CUkmSVYZGAX9XYUQ6ey9BEmaFxCRvcpPlA8
i6VZOPnwHEzvO1STVHoRSW6CN1rkWw1T0ItE38r/djkz5uESWSZcOXO2NjBN+Uc1yFR81MMkQD9v
nbFe2Sz+blrfbgpKTUswqnMxA9XC/OCGBn4izSmmzm9Z+iEkJmRY9bRNg//TvYwjnN5XKR2MZzxy
EHTHYcSwrWzr5D+AHohJG5YztzmXvGi+8r7izOrNBsbrbPRZc3SOu1CiLJagvRh5Zjk+c3Qr0PCt
ZUguJz8DHkiAh+zYSJ/sNxn0uCQc5FnBdXXH9Lu2oEar74LfapGsvEFfqtEVuQXV30L7sVnJRaVd
5AyPx6pOGUr39gRF9iI9UkVnMfEJgVr6qK1kLO1xMzaZ+XCFGADLK7Vv7lRkLtu3Rhm05cpAaHKw
RXClyi2tbdbYTpWc3Pc4bOqIYz7Vk9EpBOKdc3DIyoEwWW7h395Po5uXwI40cfqWdRFmqmp3FfwP
KnWS/X3DuJ+6frlbekBAWr6hIEScJ3H+NCrJRl83hTzM1gtohIk5OqLBWP9CKa+Bov0h82/EMSvc
JiekSL8jiMth3uK4dQaBCFaraK946REXaiJtXVogVtu1DWFDvYpEWHZaLufiCQce0eJktMGTrVoZ
EGHB20qTFGu/VjPMynjS9B2eYLnE3kCiBJMOXoSShc5SDDqeWTPbzWoqvkQw+EBgjLpz/12EiaE/
cO2i1ks3kcV7GyCc8czDWOWvVtCQS82ZaqTg8XK9Tq9cKcbeOHemeiEDH1apCUplI9V0jBwk7S+i
aVXZxO5X/KGPhNnZm5cEo44exbuutAhJ+BFQuM+APc7hTZm+NmW1J2/AhVxI2tUltWi5KMQwkFMF
/L+eFr1l1xOsZLCE8YX5XPltejv84BDruOaHOEhedtaUUtCyaj0j0by/MjN6NU5I6PoqtBEPFadx
ot/00QRMqg2SM+LTgDPv315CwfwKJPdoSr4cKEs8+xTTovuAxdeJhBzUYX9pGW8ufL7OkRoA2xrt
Hi2DoSqH/Ng/WR2ve6xfd1LBexxCFt6FLOrSO26Ve91QTwCem+f1YlClwUEA92mesDth9jWO20br
6bz19dMEgG2VuOgCcXdtD+LHFF/P5uS7b7Ny8FbF47pjs0CT/+7MZPseCZWR1IjLVlOl/jz3lDQn
yrek6wBlxsJWwTR0pPXn0gNVxkhBpeNhsUvQAfiKDji/gcoFgnly34y2SSZpl5Bu1uRX81wH6v6c
sBqOEeS6rzh3vh0GeWSHTWWMvRrKbqEx0m++on2dpyH0D2PVhTZltJOLDX5ol3HqhvilvQk0SSm+
PtZkGs+AbdxYOPEKxGILbCc5/WKDyeKxGUBDYpVlGTvz+sXAeDAI4CJQT0oJdc9DESsbJ7VLvuBy
1quu2tIeDR0ELaIeScwPkFp/vaGs/29WkowlA5izW0Pmb2hurFqX4eOyA9eTs0aF74mt+nKIaV+P
gdxN9RFb/xlp3u+PSH+6DguelZdXwkmIIwg/78J643glUXNsyFvF5T2WsLRhnAp+IzbLzDXO7H1l
wcQMNEizNopbEhcv/CgthF0dB6sPYifRGSNB9I0jUGExiLxcBYZOMQO0kbY50wACCzJCsNxFv0WA
hV1bzMHQejmgsjfdeVMKUrghi5RekS6m3z96Ia0QL3c0vKzmJ4+HOF1bPFN/t6tO0FmVuz9FDxUr
lhNyv/+Y+Ig9ZgTAYDnP3LIWeA3uEBtND5TOo3Mqeu6UpjzrE61rtlDy7lQ7P/W8sgdUzJ4kIs5r
asLI5PnBIgMfTfeNZ3KRKm/0bHyGgrL/m13K8WzwtM9UTCiiSg8gTYbHg7fjceEmPl0mvGxEtSJ1
8n0KFkjeCdJLaVKJFsuzASrFpt2UcpcqfnP0B88QjUIysV3WCAQRFU+ZM7r/VjKhLWFIu5rJMNTW
JR0h8PP4nUTQnqhv4NAwkIMH3MxHFsUo7sagqYP8MdgPEoNPHLoFTLOAvBIaT7tgDbzRZkSSULog
RXjsGh9b8fRpTC/jTLDlgKSbiyNq4IWnfjrQozyMFLfbsXEWiN6wcMncasyYsMjw87g5kUAjceWP
1FeyZnGeUFIwEWjj3+xjH2VXQQsIq6m4JjlfV3js7FquL6MBciS4+Xe6bvuqPa0kygq/tb2kjQfl
uT65fXq9D/DjoKR+vG/Ij2LSdMIk5UT+hBbtB8D3j2l74nKgxdWuVReNs/mD1XwXfCgPdLec+Wjp
xvDzNhUR3QLDKiK7x6/UIMZa880u74HtnJMza9sneQKc8nGzouXmKWyKR5ZHYVpncgZEre9dLi9B
6fAwpjQpAqHgxRjhKp1Yph3zVnja715yg4bVwzAaxfGEtNFMSbKk6mzrVT0QKmohNvyPr+1kbdGN
TAm4q6Z0XVSXitIetn5Os8PMXSbXezcP6hOc8+t82B8CXz/oTe8zt+iQBn3emHmKL38k+8ph/piG
WQxVoX7viFf9U5CeKw8FxT3h7WsubUa+oW8cG8fJ5tKxdZeR35BpWcTxRNKLZNmBiSGifpE6x4j+
edEYWMOl22SNGZc0+M1lXPzVkZvfUGxT9Z/jPofI7sgd5Vcmd8X6GxBRQCW5ljS/GrBZ3B7/LHfA
8D8FbS39KpWG0jdfbanA2qnf0MQJXnjRhSNUX9W/cHjf3NekpYQ0jkPgQ0QEUlihPJ3ltGt7YYVl
uOmZwWrgI0WPIQ7uFJfGtld4H7H+hT2QH+fl78FU8Gsq6GlGsGOcJzXSOMsyFeHDvY3fSSykZPyv
PpQ9k9+mtU4p4jWMGMcXygcP/DgdBz5TuzrCe71FvZPhKJx2UFv8x8HxQpi+NkBgEVxp+NPMMkEp
og7WPP77qIXtcjMlaqZyfESsLuhPTBd7uL1GUvF3vfgZR4dKV0S0sdq51QbO90Pbwjvo+coYDnHL
PATiB0gd7Kp3hntue1jGIjanVEMotHMJv2te9fn2US5T5YQJI3PHznxQTHJDPUPQaErau7gkrz2M
fxbiVYbLpK+Wc2OHRMgyyOEF+XJoP0whEzOGi3B57bbHLL5dJ/tZIZuMVxCtSB/kLTI2S11NZJKG
dqQ02UcGkQ3GpVqpCIijQnRwkIfMTX79iK9RHyADPf/69/eCoiIPzyXoo4VBw3f5YWiMVWecJbJ+
Un5zQjCBNtdyX8nDqdw/mPsp6CZ6uwY+yyMEozvRbl3QAQcZoJO0ZVEz4nS2ZScDwdpMtTZLB0bQ
pzd09n9IbXlrofkPqYXtVBfbda44ywwBiyJ5NufuasIcEQxuqZVnA5YLyQy5eQCBm3xkQxlQyhSv
tT2BFxCT4MbTp0ZdkewJdO8TZ4v0C4D4/l9IwDEWaa67k5iZnH3uM0zuznXs/1pEJnq3EpWv0oa6
3onoiHrFRNVoEgFi83jTLq7PsUgerGrVQDQdd5M2rJrZkj3E5pXvLa98w4+ErLIO3m3q9CCHOS3L
QmthUdJu6gDnmglmQUaRBfo+i9kQ+y3IpQB3Rc49tN1wp9e1WRfRk0U3D3NQZ7BnEoTGJkwGO+Dy
3UHJkLmZy338Tbk8BG3fKeZhgxFhwiayoLvsGydZky2KLgJrVIPWdSCVzDaRMrXN1mnIY9dxH6Bi
td3HjYn8w89eAHFmSkWrZ6k9syT0JbvMig2Di7zywEIpIsUKlVLLMOjBGeg+2b1QeyIM+oNU0xGn
clWdQyT4WiwH6A9vr1o2PVU3V2xukROI7o8coDXGQtEG9sMfMojsALYUZAT2f4l4VcbXV0T465QH
lsjScliIhJnHPeLNNmOmC2PLOh7j1AcdgqN6wKpbCzpEEJdTIyCRQEzaq9DQg+ANIVV6FxIjoa28
9VxZQog/hAPor8uKncqLE+nPFpbv2mlP8Pnca+j2DD+cC1VIqmyc84rVHiMlh+8naxktqILYN6kI
m+L5nfxTn3A8QQVMs8ZnHKCsews4MBAzUtJ3lV+1ShcxncjfJl6X0hx1z4lIo4XVjI1oxBJ7wzfx
MLJhUF968/hznJqjlbZ/d9rKhLXnDq401QuUOoTW98I1Gol1xyndBcVJyg6SKAr1t1n/2x2JsnD9
uXdBVRyPRnXU1sqOD8l8X4oZgYxu/ic0EGJ3/NnAeL4BS335YoIM53pQVwSY+hjoYvIz8Zu5uAPI
ftbQIC+/WQn7ZPW9PfER+pJEtnsTF+TfKDV6475hpabf3fl+xKdLke/5GX5s+0K9Kc7f5yPt41Dr
qey0Q0mLc6yso2gU/QeNgmOOWWhxPnySvHopQUF8GQ7vCxu50mSGzdt7wIRRoIe8OwXPArfn+k+t
qJG5adLKYFGq/DkmzW/fx+jRUVDeyDGyXmOBSXfjh/G2TDhlsjnCrPjbUMchKHVEZNIREfqEn+OQ
fHnd5s5PmId8MbjlalZwVRO54K2VH7o+NrdaE/9feeGbKspVmd6lKBjtF/gANtNy0daji1ICaLQU
aGzNwRY6+Mf3iTngkeZalYgR9an9x0nDYL4Ms6S1eZy8s7figb1Ban4+7yfg6z5m2O38E2t08bTh
PKUG0oLQLpvNSJCNGHhQMFeToWYESOkKAlVqNpMmM3xst1yWJrB9wNRg5kyeNT+ZMoDVkRO81KH1
9xyoq5ipLot6KIEycw765bY3Kz4R4Qu0/zd4VY3tDDFbGlCqN/1xBqzR+rac/dtj2lCTt16dpaa9
2a20kallTWCrl1QBwLqOp8f97J1ybeTuLoh2IDYsjD67OU62Tko1HR+jNbo1eFk225QbrNmRsYea
Z191Jkbe2e5UU1mpYB8y0/ZV6UdptXrOYop9/U6sfodJR38od5g8VV3pncT5u0QUTyymKZRsbU0K
F4sNLF6jVc2Fwj+jYsAFy8QzYWnzedPeJwp7kEAfcEixLkvpUWkx0/QBeTotCPY3pgEyK7fSkq92
XkXw3pYT/5omtCbdxeY7s/wPdepbq0bTTIM5aadnrZMSlk9sNzgBKawa9bMqQhXpaRStmGSIcHd2
/JVqmdw1YrW0bT+xfd4iJwrvIwAvATsgW+VSzO0YhbN0C7d83FTl0g01zGSuap7oED7ni3himDQh
1z2QnjyVDZMWDoAFRiEPGHCnepZPlPQQds6Fq+IvCOJU+HZGUjryW0dgn6jEUjR1APv17ekkl1QH
n7I+U2wYfvECf3lWrNIGAZvbE9avxNGmyTeVE+DldjRl3gz4yY4K/NLpBINWFzDieLHKx+n7WEXh
nClx3SUzJ+VH6baEJ+ffkk9OY3nbG9pnWFpiPAzU9gG/8h7SNWDlSihwiy4/LOpZGm3gFn7yQMFq
f/9U/Bf10Vb9IqG7RkvBKKJILPh6AP5UeoFauNu7FsZbw7bwGuyrNCV5cgpJ/4d7zZUlFhNNn8iO
0/UCRvS3WOQNFuHB7aQA3A4tDLaqXKoLkz7Uow/Ggint9iXqyc5wlRUaPPHtT4dQDHx46iKkmaV8
415TN6ksg9YRUPmidyKU2pU8Igv8lDY2osSaAzzPari75xcBEngFu7sLYMl19gZpkO4HdWgOci2N
LKzdODF7gyOYnUHAVwVKsGQT8u2W5pMSkKAg4shRjtIZ4hVxg9QGJWQXchTIUQQfKl5oN8Su/SnN
zqD+YXvVuBQKFmEMLiLIFU1n9UG27tRWgvSVIiyrVd0XE1NpIHT2X+7CSeQWXSNYr4ecKPHUzPHW
P+TGL2WwpqLmMvdtPxf1XB6WMvQ/lX9rTR6iR9BivGKhbQREyx03vSLIeaT+0rkO5QLYUccPMHjA
f6IMpDDb8vIz7Oc2QaH02ufEGf6JNPCIbgwU36dVPClKs+P+VdnrIVSlr/zjiEUppnsQwl7HBhJt
YXnHWtG7jCLc4DP36UMMXteeedESdYlh3rHH/GoaE4oSTU5VZLx/YUPzWrY7ZaaUTIEN3+YDq47n
0yc6b94M/ry8PQCGUA/5o98GDzEd4pdfMeL/DLR5boOuw4Nrae9SE+0Z2O0Qy1cP0gj4TdzklKTo
d7xxeajCMC/hz+XYZuZSXpyS7Z1IX3L2FwF40bQuKDXvYitWEYDnDoxGNsOwR8/2rg/DFFa+MbSp
IgJHauF5iABrVpn6ALkBE7TyD17NGJkAAuL3QgjPoYS24Gzt0PewYHP+t4LvMyLOEx4Bw2cLKbnU
utm/vyiC97MOclCFaxvJ1Lok2W3XzZvy/anqRSBhhpWnK+WL57uNDk1++t4Zh3zZ7Q4NIvWACc+o
oI54OIkxJWUQaQyAerleI/1hMylY1kz+JCQXqfjEGqJBa1ojEwo7Ef2NqyLzk3+QZAZcXCi4OR92
HOlowtEItKLZ2Z8VyIn91+Yu5Llhm0ol2ZHYQuNSAY2XjkD+zkWPYjN4NW9ZP50qjKGHBZQqP0ae
Sl1XBYH3RqljiZMn/qrsgfG6EfDR8GR6/UE1+SrPgceHgk+Ms7yIVvsFIEZAtfpNLUCb9R6pPvcy
5z6m9q07TuQcN8cs8yCFLEdTQI5/ZqoMgcAfJW4jdC2fPIWZ4Fq9EOxzFBScePm+Hui9aRigCIWW
Y8QvbqYvJIrZe4qzB/IPeTNglwEznqLgwVHVEgGJmx4JuXedFhjjbOjYQ6g0biE0BDn+sdHcfUbN
DR2Y1hxpMPifkNJCvkSU7zlGWk8qIh7ghPD4f8FgAmXTMmh62+hHe8q1RBBWqAqNXfHsmpzSkLKQ
auHX88eaxoHN53SYAUJcQr6uOsgxabvT2DRdTXVH/fNzkfTYVOPS3BvteZy4+/WO+oopzis8QazT
frsd+KyjQljZxkYV+7/l1hEVH0RRmPdti84iJuXeznKDzOn5e7i4mTfSq7KlRlFqTUoO8EseKD5R
P2RzmEW62ZkqyTKSvQhQzzMas5WnrAUbBcPMXouuNQ+iR3j+ENvGVCDDOzS3qGHtp1M7Ivyqigpc
Y6lEJ3R7dwa724Q0Udy0GpqA0yQ/YegLvMxgovI/O5xVHcg/BF8OQrcr+gmlpV2omJjGQH2l68O/
WT/maa66Bz2BXBAePICFbw7xYQOrZ7xsShwMlvPRyyR1CZDkzGXLTlR0dsY/JhknZU2+clcgiPaS
kguetOU6cu4xU7mlrNE1lPEz9080WYOZpJzdVPa/627q6zWltUmzFLgqiJ2LWhu9L16Yqz8pbIH4
a01n/ydBFNoWIYxQMHk2F/J6OYzoCb0lZ4aVkJFtF7fwdiTUObERp0GP58UtEGbHwo6KdaxUtcix
w8/mOobKJmIKokmUPcO0Xxeuj/DogkKf5baVK/dn37lY/77nWHboIF/feayHm1WKpb3cPnhmEfKC
K8teUVequ5aTjFjSunWLAmr0wd5y+ifomNHoG/20LQShr3icaZcsNZAyUB6r/5DEdxIkaJVhuSZi
xC0YNJQxPqp/eKu9xgcMg37rSVVZh9Nl6yeiKMazhWcdl+8ypxmyNxIL/466st1uPBybVlKj8Hq+
9uoBhH50oDx40WXumeX1xCw92/7QC+OMPlQJLBRft9lYgEmUCBvR6JKc8pFl7TJAki1DwRxfAt4J
Nez1kJ+fGeZWa8Gbh4KkO7PyURQSSdKWiBENxsS9V7Jit+fGMMt4SRim/Ux4qA2kDhDOWx+sWXGX
cvpSmvGfywgtqhnqeRLKh6HPW9VAzSSbk23wIUuViP2DqNgyVGFlKY1quBoqHuLOpN9I0/9tEglC
7NwxCH4EeYkhrzdEOXwPgG+Mr9D6Z55PCZjQdBa0Mu2fHylG012aY17+r320S3gOlSNjMrmanUQm
lBvnQhPdSnJ2qjQBei2ttYJxxmuxFTK+PTE/9Bv9adw3XhsYwtmIUiBaYzKaXk5w5FHFsd/rcKVr
HiN3iIXO38k2n4jkDV4jj6pg+lZZfxtfjQzKJ7GiOxvUZX+YisdqMEclTpF6ZyXrRQ5WwW7/AmPm
gXZfsh12+3Vl3IjwhPCUA0uZQX5cZW3IKG5kNJmaptj0qa8rGdfjs/DaabK98riGUItOqktMrEo9
VKVuif9KaprfV7HEZeoNevS+JHpatHSXsyN1HSD9a6MwQxe1tAkpP5XG3vsOszA9tukv2nky96dP
TbYml89JdsBVLLynU1Ncgt2nxADJxhFAZTibTX5+ZRz5857navwjIMlKR/Y4qaMt9fI3OIWOT169
j+I0h+M7WGkpAHGNjR78vX/U3Iwdb4FKrj6rd9nS5UeOvq95Yfwm3j6r+pdm82j5WODTeCwr1kGV
b9SmoMAlJNKp1FFDzYsF+pIa0LdwY+v4GXiShOFNRJG34lRP4IzKO3lwk2GkYhrrMzbeOjE2tRJP
xt75U2D0llXl0tbm9adqVLvsHZg/ddhZB1t7o7SudxVJaExlEDsmciHowL/fQo4+ELByn0VEaFS7
qQ7evIeqXDVn6tkG7BEt9odbxXotnBAFvPb8cWKj1jB+OhdMlyzrrYKSWmnVBNkf+EG0t+8vnacr
kDN6exdBPaoi0oltF+Xj/gRDHAlrFOWgkiK8QKI8iuDCM//o3AmpHh6wkKOBmjXA6C+tTuLWxuZ9
cmubSQgHSXvw+hJTaCkLZvZzKoZyId7WpHp93fBS+HiCdkJzfdjh8IUyptZm9MwstzK924fUnSY3
SleGW5HFEgXnYY6tH7lUXqFd64SQYXpOzi61+Dg0wHdpxmdCt8qYEXC5ztgFE/qlPY5xfMmMvwHe
XX2rKtDTaqvSGe5nhnCXh319Moiq/kxJ7GxHGPjFdN1RjKtbSM0d8o1bf04u1lYVptGUEowxTAIe
zOIEXRVRQE0H9CSAkJguVZ0MAG0rZcrqTqt5rvj0ewRsVIgScSxVjDKPGAuNDxe8dJXMkIc1p47H
bOXU+r4wKa5lCuAmlJKIw6UxsEmOb8VUN4t7sq8WF0MjnpHOYyH2qvuQM6Sx57i9bx7g26OJbIZH
qPSLn2QTV/u7oGQwSefLpalHHVeB06sLsoztsfawIIQVhPI/jH19XYKNRKctL3FUPS3EZsCNmII0
TzfDaA8X4yv+d2UAi5j72tkC4mvJeWAFnrO7Ozq34j048OMscrmWpqUEEb2BtCEmPEhXFXmNe8t5
9E0UT+3TPZLl8WGCvd+Rgtdf7ze7OWTSKlP3L0wEuuOL1MtEvOeXpjSHoJMw40ccKCguvlyWYu7D
B+ocOs5rRnxf64G/2teoKK7z92yHjGoOzIP3wkSRISnDguDOoAdfnu6bI2q+61KS+uaRRWFqminP
zN2kuSsi3B2fRp6q56pp0A2UlgAUhg7lXFGqYJZP40uisG9iaQzImYE6ExgZH+XDxi+L41V0FLTx
CZFIb/LY68Dont9xVwNop3pMSR0/FWpelLlSC9kyiJVI3LFBgIU+pECZy3BmeoKbrOqcd1BVBNy0
4AlC4S/F+4WUC6Du0kUjOe0x9OJ9aNhz5YFe6QhMvCkvWhfrACHbx/FKbLA50ERZsoaQy3aWZlMj
/IB2LJUvgOJHyJSoMR+KRS0TcLX0yiin9Hk6HKMe6RMPNMn+TxkSxH9tB9g+sFRYU36fuEQP8Q0V
X9Cicr/dTaRBxWOz4x2xU8UqgCHAAgO2S6y5CL1uGfGFar9/7dwreoQWCbZRgIvjvU1+aTrRXP7a
cHtRuWJzlMaK6YztY2NNQYsHNwDyyii8wLh2N7Y1h/kezaQHl5gG7n3jZ7TiiZezMwrDE3WZ8Gqc
hGER/PmdIDZy1Wa57No1Pw+8h7gPQTlAr6xvK/A0DLzabUdcnsUtvPJd09GeLP3UUn1KopGuE5kS
xV3ifNFayUuMhV6fBSzRVHKbJD3IbzXJzRsjMNmFowZq/MKoru30hnCEfzFZZQCSZJ8IQstF+wU/
y6TGNfwgmXKTmW0Ugilpe8deg0tQwC4McxRm09AWFVJzY8dcT0HaTKoNqUFOexh4FnffmgZR1qfM
vY6P7NV+ttpmnBVqE+vAydjd9/WRakFsAZxJOvbEDzZ22ebJMGfxhCq5REvWwZikxAeEV4VBLMFF
/G672kajtcSxZW0RVNQrHGOK7HJ/fZonrdhuw/uFfXOIO+F+7csOMre3dXpSitKL91B5DUlrIiHf
Bg9HFlUpPKw9iIf6vDEdItJSzK0wlqxEAM0JvWWY4WwXHYjSiAiPaTTm5gMO0ZpRevhQMKAWbk09
pJFiCbXfPEmRg5wUTuQpSgIUmT4tJTNtrkwYYCA8ei417iVaMtt1zNwm2Glcxlqs2miuh3Cws7H+
N6OU7Bmfu2GZovz/OE9cCX/Tk/m4KGAv59LbZo7W5JsjC5Z45UHCUSHu62xSvu4OI8A+pI6n174U
H8ayajZ8w+NmnHqL+803hX1b1q8/7CH+Eg49YWAcUkHkbTm5OpIL9E4BGo1LYv2WKW4FSWoI8GpU
dRt893Sohi015udNZj40YFB+4v+ULodbkJ8nUi2E+c6CyxVcrAMZz/bcE/wvH2m2JOvSq8PtTn5c
BgKP4M/Lu9Lawv4AkJBEHbyWQJIfNclWrESxT2H1Mm+//ONVvqZOMuk3JrV8/sbiBo2OqwRhoGie
kHPsMlNRgpvKWPJO+mYCl6tnGkK29IwN2gUKVhzKwQRtL/SduQueP8SkxDFOpeEwjNPUM8i9XV+R
7eIbbjSBI8QBQFPlLS0GVYF1oEPks4tnhmhdq0Te8NHZfi1gg/Tk0L7qFQJU2N9nmF7Umhducbsv
FK6uUNo7rP5py+rH/vpaTHR1uCWbqJWtaJnW9oTO0i1+6OYXgcab/RSYh9y80pkmsSYE/7Lglmvx
2VgJeqyuG2cIn+cMfG3BbGFgKH5IsL3i6uMkc1Y50rDBkrBLV+r61qyaCYXretl/TGTi7Tr4eXMj
4wYysY4eTMsAOz0sixu5GuJ1we/4pyJMjQji1BnhmHHvSouvits5Sc2Yd2Of+0aKJxRzhmQ/nXON
YPsUyIRTh2bJIo1gZH/697gLaYCYbCq1JpXWiDuASaKKojo1qzhjHanhSyIpxzEcGADquPk3GVhy
zfwq1PN5S41RHUK3qIpmtrkTOYTvTsvtGwuio1egHx668nHzsobAMbwyO2tV11bIfHimruu3pCjd
IcdHcnC4gwLDxd/AZsrW3dRvJxvvTsWztc4JPoRtjsBh/ShjItsv6gLROL53WnvbSidQxhtfODMf
jeNj3hJecXKUjvNFQ42IF6rj0Ve5A27J5W28pYSa0b76p8BCAszBkp7zL4olDe1sFiNcop4B7rV4
nnADrL9vXjWUucUt4ukU0xOHOa0mtGmnDitYYvfPv32MAbLUzFhkEHeCeiynZcQQFXgE0iIbBqVC
d3eyl77HAsyOPpJIsvYhjhCq1hJS3+VUAcW3kKdUJwbpu9Wj4rzeZ5hNuSbUa84HlfOBHcSG8iAf
aOypNtmaBWft6tDpIxHFRDgVLdb+2wejB+DFA+Bt5g0XBAvnJn3uZKO0KMOfVuFLaJCPq/j5Gh2n
UOFdV8b23eCk/NSZ/9t5Yjyo5tcqpTMUlflNoJ2DXs1pEmtdT6D2AhhvJBCeqPNjpjByeza4oUc4
IJbShBfV9Tl85xHLhMKj47dUuEd+goibHgKTmFoFbVq3Hmkgyta3sodIApuKcCIxeP1n8unrcH4Q
F40kwkYQwaFmMFvsO61cwsw7XN9acs357ykdNVOMeINpg9ePMRzpR3EWBz+08u1pxuD/6m82Wgoe
qBs5hHYQFsMPe2oA3MMDK3ByYbu1Zq+WnyM4hWf8OqT05x5KOm4RWaXDLMXQyOmFXIpcGpMCc++W
wZoi+0Qjp+7uFZlFaw0IR7hALR5p3UKjd++FTWwuxQUZux2h/V5bku09HwuP2OpCLnul8Fp1mtNY
2hVqFUI1NbpEh8pR0/DRX7dE0Ah/luW16U0kI2dPawRGM4UOv6fu0C2f0Yb31djnO748o8b23UYB
O6VfKG5DZc0w8KCeUyjG/fdRU6YcCHJcsAWf9KaX3icLZtKYmI754i5gZ+fMG3nSCLxsXqv2BdUB
XU9iaQ9csRAAR7EOcU0AhP7qGNtCcRiME5JjEfY2u1+0vLnqa9KyeXARQXrvKCewm2IAusWbpYyJ
Rt/hjv42IkAxpCRJQfs9mBw0xnYMhBzlofBOyjdQxyBRxe1xMB4VCmzRgvrkSRNpMULl5pv/XKfJ
J6dhIiREN5jQlAwZlVrEr/VWwmmNkLa2WZ9eGicSthj5ylQXpFfFbNiL/G8ZNqIQSJQpQgd6XHrr
0gNOdddYC3QyuTwlmOgp3Zl2BWmzIpoBUCsg38zUck56yXZpEYYJUdJaXnmAcj7CG6SpmR2eG+sY
akIErSBu1P1IMcRjd5/Qcjj92yZeX6WAdtWAkGiHL8Z4Asg2lzslK/ngeSlc6VIa0hOxpfBEZaf5
oV2ThERLP/xYIqpHoL4eliM2sYZyh1pGK9VZAjRqhMZNZeuOJxM9Hjlaoqmgshh3btBYETnT4kkz
ijILOj+AgS3Nu58sVsut9Fmv4O8FrDpoaeJO225ty3G0cHaOYTfaA6wRRvwgPLpXUYvAGZPfvoA9
vOYTZnr0P6oX9QTkK6SZv3wnZViN4tPqLmw2KkOC4SVBK90l+ipzmgNoS0YZKCpVV3xCZhhPPETV
Pq1EGdAk/LaoHKz8hOIsBa42DeWCuIU7/nwitqKAjEuly1u+Gh4D7yDSgd29N1QgxuvZv+BR97C9
FNFnTcsiPmFD8dsTCaa+kvf9C0DVV1crhJ8JgxfbCvZ4XPP4ULPt45tJ7ojnDZdZyaubdxYf2WiH
j4XK0zn4TFP0j/aW1TCTjjCBOpUBnFBQAdVd06uH9eRAIk9D/l3X5A4HiD+kc0nr0+IzAO93XO98
YUzFHKtTd61HhX97Os0Iucw6oZ5my2Qgm1JKWdHFbY3K8x3r0regmIzqc1w7weHU16hQaXnoeyBr
qnQJoIeS35UTnzYmW809yareZjzrOsBgWJlT9bUos58La+cZZ/kCYoLxv7R6mE2/Ydlagfgjy4ju
oX3NyuAgT4i4byCvzhHFEKaMoMrmh+gH413llZNoMDTuBkaBlXNWlbYaPjooF2pg8fbZijdBlPZ1
61KGMiYp6fQluDr9AJ3Xqdqj6kZDOSpghgJv3szPXcgtAjChFP23CHFWeOdkh6Xd+34xKf1LvG5T
K0zdX2XEgp/VYDjQT1sttlJN3JH9h+zUAUA0TW5qvWE+idZafXLu0jl3Ns97wFXbc5z4nqGvAlu0
Hfr909W7ELSSO7c8lGAaS9nO595GhL/fnEB0G50NsQOCbJJcrFh/s19bGkXkZOG+KdV7H3R68GuK
VrPhkQi75gOBYC90NBs7ohyjiK19CwgFLrgdzX9U9Gul2xWiUabLq3hFxNXvWeGp9tfe0++SnSD4
hWjkteT0mYv5g4iVBF+jghJF7KJ9Ob6KmFeNlcYXmBU6k1ToH+8o5Qg7diPmwRVsl8Q6qG1WI7+J
QZCH/yHA1R1aSgNGYmZLgAninnxuBKdQlgsVN6FWkYWYWTmAdPLSj0dgajYXlU3ysh7KYv1ZHUQZ
T+tcYxZJbXhq6VQmSD8q8F0CZMpi3U8pLV1UHESnjnKiPW4+6AVLjjNWPCF1iwEe3n9ktMhGUk4J
UCVmrzzQRJatNAZoGy5j13Dmip8tvMfccqRjtFn+wSCr/Ok8j7KJZlTo1m6mnp/r8E/73kTjg9L8
UW8YOVD06YtNimBkXCaw1OSxOkka+TJ5Tff8KGcvtEZ/PjAIXw+NjVkfWvYpq5CZu7goh8fDIfI7
qIv5YtTDWvTjIzLlLvZ5zaNvqLdk+8AcCP3daTYtj4W+XTnC7yOWIAEHgHI2+aLKEtgXPe6TZJAF
/IWrhnCxbScXbadB1672kjxi1nkBzOrq0lFyUnLN74iXJBJ7JYPxAkh5a8J+7SDEZXY69UxcofJB
kztPykLFEF3Sc5QVex/KX4RheKAjskNGZI4KNyFL8M78MrjU6Z5yTF15d2Yjdx9aDCBjvimRjxrE
YUzwJcSeSG5EfyPArAU1RNcr4NC+5D9NtexX+7SFHKXr6arYnLQBiO59EjiWkQIu09eUt2bndWJR
VO71LTERwXoOOpVbZgi1qmIHhcp6Rhn5LY0XAU5f+OncTHU+i7iTKXeuYLyaVuG+RgG/dqjoeZX/
p8g9c51YaqwQJkAglixM3DqZ+M/8zWbbFSeGCRqsm6KO/Z0a4ro4En+qqM7ip0aL+6LLBSztxASo
zEFFb0qp11lz+eXc0lanNjcRl1nTjmvtO4wXpZqRz9cig2aZfW+2x/RBVy1RVAEr/5hbs981DPQe
hd3FPLsqs3BQAAHJwyl7pbG5HlgBQCzUJ9jorzgWnuryJQSqc0qW/08fLXYOQn7ENIHl5FOnKuiS
VKHAeC1M7IB0dct7zLJdI5N4l24G+/+kXoct8HURa0lgAVrtUlXsaNHVwk1C0DOdwS4RFRXsK8rV
SoBAekWnD1o9vNMAHlvQvoipH51hC4auj7pOnuwu4hf7x5N7MeXazCrEBHZpIriWevgMVq7XvFjV
GemkwwFXY4ZVSmr2yRxRUFg6DcFgHoX2Mkh+tE9L0Ervx1fGBhkwIPbT+xMl7CJHDjMQ5mRezpuT
SK75RHSxl/UAyt6V4LbX06AA6Qeff1JESrTEf2T4l4d5Jb2aqRCFv43F//khW6Pzeb00uxypeMhd
FESU6DfyMAAjoSxEieYy2Qh9B5OR/jkTngHble2XHPgkOPKwnxze/RfYzO2KSSx0ZGwlz5VUc7ja
d2DKOqTgEKFvWvGwuV9krTJSNSdfPYmxpMZgO+bhAj3OAfBhpTmzf2MkwXYXs+PHQRrpvX/RZVMR
GhLhorsGtsiKb7OWZL7zJ7xJLHsGVbO387Gn7flEtNbWf3Ey1yVFfIHFu5OrKUdkeN8U3xso80Ai
xKFBWKpt2UFDTHYBtCXNN9lNrB+Zz/te9P7hxvzMoswHEGE9vuODi0OVP6q/19yCQsYQlAvSnaps
ZXnJaStsDMWgmrkP/piclEsTVXnYaPXrEB6DNW6XbD5N5OQyajKsoMm/iiPlhGOGCM1ldoFE7aVy
Oni337YTz/sa19/xvkPC9NzussBzspgjKb4UJlPuUyq3EW+ctKdnVkDpQAtd5PK7mrFxv4Qi6qJC
aPWg1y+uXJGfpGAjme3ZRHJMkgCMwow3ATtxo1XVcmEFYpgIwILpDg75Q3rsOv8ys+rMMZ8DU7lI
AaUknWrAS6+xMyEYqha1mFTEPfyRZddfIAgvy2eluOx3fKaQUrNuDs5gF/boi3iMVaeiQrNibMib
JigKp8WKJ/ORedQo+VbvIMmnvjBTyUEePjPJ2/U9L6gyF90kVoUmoKFBaGKySTm273qlvZLoIlng
nyz6vu6kLWvlYFZmm6BnBIX9tJcGC7pytUimipSqz8jrZ5QLMnjqglZPIkvSbwTGykyX/IezL7FE
ueLm8XzAR0isCprajlFMheGZPp10mrOwfYpy3CV21/rvB8zAxWS3TUBe0jnD1KAoEsMvC/JZkXig
spH3C24KrdzHNEqW97TYy8xmcoRVPzDH3a7IG7PSNtVPSKDNmwfmoiC+4XN63i/B52Jg99WuQ4ps
/btVuomoPkQJv+s7wA4NtQwSi9aILyWTLRHV6GDk7ymCogvFuH1Y2LXbAEOI2gVM9wJDxpECQJYp
f4svcD/lPT8kwHGNy4qiBkK47z6Gtf7qi6Jo1eH2/1KEW+qYwiGrygulZVr9Giu4lT+isdRFVXQx
hQthrUl6usYM2mBqcYd4FdUd+7LZsZnntfbHWXDhF/LNqV/goVPxRn+zaaoXnKEZtzPBlpb1B3bD
mtCve7msbAAld7E/f6kmg02qt2Xp+J87BInCrTOzZ6jXvzZkzfGIkE2vkKvw/oQXBTj1Gl3BbBXD
PbeUgsPA0OfmXKOtZQCY0tk64CeV+QibVRQd2RTPu7JS+0lZEtklhixZ7IVUn68c0R5MjDeIbmpM
3H4Mr1bRhxuA8C1WdUV/m+9cDKm5rt46qeqJe6pXGTjE5FJEKW6veEm5rbmURC0T5c+P9wU1qvFB
oGFPJYikcl5UMGevqOiinoo1ZZxktYTle9lmZ2jTthWOmi1aKn5lgN58Lxk0mX6NSTmI73uCPtpQ
sFsagEzvefURFzr8scz1WxlhnryEJf6A2GKMZS872z8HrZl4QfHu3veSBcZsTQ3HGR6M+iqCgLBC
LcUIv/0hyGzIJV9X1YNwiXDas4lwZEeEHy4fs3UOAiSKNsBD+vTG/DWUd5y6W6AJg9Ml5/moTPry
BHKIAPdW47BF9lzWvtkYivNR7OkgvN85H2Vnn/zfjgIuf7xDHjk4WFaLokHMEgKJgrQknjpJm2Js
6GPpAVKIGA7JE9TYoBswOq6GNyWcS1sQucnfv+2aKw3cybuj/2kWZFXfnSdzX/97AWrsayWVvsDA
OfwU/BBrOr8a5JeaDTUSXqmbAq8U9vwrYdFpxklrnPy5DDXGSpgNI+/JVvteR0IxmJJt6luTHb6d
DLe3HZDqqbI0r8xIfQyb/npXnZjbs5Mr5UZBhxupzZWqedG3O/59dqIRAF3HWOTV/OQ1DUIwvk52
exrikVpfz8dUlK5sBDK9Tm5M6twtv10eJkFWBFzyV6q0Pbqr1OBRDG3ZV3v2erBCMHfrkvmOJI6S
KhmTbiZaFLmuPaEhi9LIzHr7YKdKeaksq+Kj0zSmZ2Y0DzM7va+krmkUZat84LtjSVfbKh2zyqI1
pQok/k/d2b5kSeO19mivNCPK5C2m0OlsPEyyQYE9zLKhiThXaUTL4GJPno+PDXzWHZzi2PSDHjW1
ey9+cq2dy5m/S7im3fkkrVXId2CWuQQ93Q23WxaMBIYZr7iabjTD1bnkHa/+KPUE7w+5hYy+xb10
A2gB4qP3OSoXGi3pk2wzq0BSMS4C04YS1F6AzU5LQLChLlgac8cTgLao6/8KH5eA4Ef7Qnc/mFI2
XldeYsmsZfJAbeaQyY9ojs6JEj/sG+Zvcf5GfZ7K4NiAo/y9rKQulUrAcuWc2QB9XxNfmfzUafpR
eFksisY0XbRN7yLx0+S6mhD0vQ9MxPLRzB3y+e7Ln2cQqBkCyifOn1NBY/C8c7xTiSfi2v1ngSt6
VQUZF5oDWBKp7QFENYIa4LSL0tH363V0PwvjYJ4Jl1+R8Wd8OpI6APtGGIPN82NVyK6EISl7Mnqj
+iJGtvbOpHKhj5OMzYCiAExCCwG1M3nID8ZYCdoR20KbWt5RwaGQ+VXhXCU5y6AvY7EhBq8iuJvf
HB6vvekR8zFGf0h5SI98fXDaipLxOIwO495hMJPBcOl3NnB+DO6rzUqzzD353kh1oIy4XC+y66Zy
SQt8r3dbz6blIBTZebe84dwkrTJKXWJifhykVYqOwCeLl8MUwYoadtrF+grg6fiS7wgLIbtd3Wm5
yADd+ct9snvGD47ukUbM7eF2s2MVQB/+OOHhwby1IlUz8tmCGgs3hA8XjvI/aRyklWXTRWALwMBx
GBll4clinC4aQ1vOp9dxTzWzrQw5UWsFDM44eeq5epsBBKIfLtUDrdpXkVyBLurz+7YOQzJ8aZGm
PzV0S7aO+h4qZ3pFAZ3u/zkLZ9tARyJA3qTAvqC1ewG4cn/XMh9+NNgjnhSrDBazsXZNj9c130kd
J6tbyVfZy2HCS61Nz060/aMEGBKrarfWeVFHcYR+02vwoF0HEL7uTLQ0d4Oqb+DmHcCIco8AOqMt
f8jheIAlTksT7GSE1JN6EL9TwIm12dxLQHRVXXFbTdc3aZxMXFdnsEUqZoiNd4w5WcWA9M6O0HoQ
kGklKZcyhy+azCjhYX/7GCps/arp7f1SYGCojp5KjdkLfmit8ttgDOqxkeYWakl0WzvFSxJSDrjp
UagjJssj/HB3s47GKuwtRJ1TjB6/pfNjtPHTpvN0T3WUin53rAxnVC5wlJslKj0NMpwbdldy90Le
rER8/+aRn24w6awt3/XzoDhYIOcAVO1FNXQDzf1gg+keNNJ4kx/L3fti7O5wnNuVCpXudT+otHSG
sPUmO5dRz21SslHTLMtwc2kLDR0fgJc0mYEzhDQoMQw35b2o9z/hQPbS7Sz+pO9A1jUZ3FFrIbWK
F3J7HprN5xgiJjliCEhplynraVJ4tYlRrnDRFz4Q31UTJKW5FNqUPOYUR/uNLGBx24jk91GRwKDN
JWQgLV3GDS5AF2CXOSncjerNckNO0oQ58vDi/tR8/3DnX6plfI5SGRbeY4hUp3TKWnbLNCBtFPk0
l1JLU5Ssd1BsvWR7exaOYwkzm4NTGQbxV7RRmKbooMZ4sy8ifG0paiQxvQ+OItvbq4yMwEJ91L5R
BgE38l/ngfdv69z9G+JIhrkO+zNy29FzJSw63cuPD5S2oU4Jeiy/OJPuE9rTZV/n3wxhoRr/mFXv
o+4xvBlsDORacIGJC0pL9dNE9VSLG046EXKTao9ZIns+Xd99g12p3eQ0xI1VcJVb6UnJc+S4oWad
6fLOuzZn+3iiDsCMpsJcIWoajWrMvSs1815L73uVv9KJtGkZb8Q0t9Jmgch/462baNnfPtHwwwmr
PJjU38HrSwQ7q6Zi5a55ABes7zoK3Tk4PDx8WurJopgG/QZ0bHf1iTMWc10eR9DyX1z0fld+2JEP
I/FrcVExjBVFMiiKg6zhwkdDHy+9rRO9gqQdmxeRydETNu6t2VYcYyiAwRX8Ay6gMz41tp47nLrm
+KySqnNuFCkPgbcg3Z0ImXSND5c6jDuVE5BWikHNA5N700lJL4GMMHKUM0t1RMnM9SJBrrm0x4mE
GFCUajhP3wtJPQGUqxUw61S1MOsCkR3RokkTFTddX8rjHEq4o/D+bu2gDhasJG9i1Z3md8L3wByb
tYE9IXu4vMgR/dinK+ZtRt3Mzuus4LJL8lcNxADkYX+W89FjEIV4HG3DrRWVvK7qjaLtV+jYUjll
o5LrjYifS/imI8UztX4NVM5hxmrss6hvJtbqnO1uiofRXoF4k2MGQjnaWFdfhIphO0/oIcSl1QRS
anSzrGhkhxF0dcxOFFZ+jd1aT25vBTM2QJPkQqo5cR4hklOWOFVljFBfBGKrgitYY1EIDbyz6NKk
C9BEER2AKs2CIPkVPV3NaGUQv90f3t4Zf/gHnJvVDRWx4YNTZgRJHzDcmOpCdAiAyLH2SWEm+mcy
Mar5o8GD1CpgXlhmrM8/EHjliaD2Ftx5M65nd8Sy0/AYbHE/mpflR9RekyFnL4vGQ2lehsPrTROA
QisL4xOQDkUpv08j6F2KW56KbI+1XMrh7+UEWJBgTNyFShDszaDx1euLXbNzDxx/OVePKbrEsmeY
wbffIakzHZpUmv5bKA+PD5G9RhMIhoKbvx1cjavI0Fel9fOIwkBGBb8FC/GQqEnqFsAreslE15qT
EmCbmUAriiop0Ml2Bl5XiWINl0Espx9vbLPSn6dpFSVSu119CHzAWxFxrEUHjwiXLR3250X1IjnP
M6AkofqjWnEYmY/C1xXAwLUK/fQM5cKA+LmMFeIt36RZkyifh3mx+6QK51nifRDREmtDKt6XQA23
+2Ccxmq90S7bbmM2Cjdo/cS0Jf3C5a5c19iU86k+Wso2X2gQMvCxro2ylG42Vqp5iNz0jQCz9w17
E4HIzkemjJ8UBqtqo1XVZ+qfIo2zUZqEGRLeTGIKgY42+NFtyrR3ulzKa+CTLbz0xPy+S0Q/7OT1
amTHyAPWoOB8gaoGSfpFdfCHrJdZvBkvxXw36Njf9mwYw7Y3wGQDj1IovM1iJrI6UPH6tFAB7xEJ
xzoaAy1/xyf373XdjZpTnKUKhbsIENGXQlQYJPB+J0Vtg9WbG8nxLPS2owKXH1Q5ps0J+pWIZsVo
tY7kmU56RAgb16Cfqt4wUGQCpSpKIRP+5fbkT8cvEM2mg9yRZeixJAkurisCLWNhcSl3PHPu9+uX
CtR6J2P6d909x16HX1SOhc18ra0dRls/+HECkYwn3RbvOURcD+pL8BJTuZSCfVYWQywSqj5g4yAq
/MCqTXo/dF/oxEFiH+q+QaX+ImWNwUpEKRKT1T6YznSU+90Okcn2f+FPmVve2oB4GXI9TMq7iJiN
VOC7sU+fPFfYjG85vVXCHaplqcOZhqLt9NGyTt7t/qFPkFmdpBp4xM7BEKlTnkK15rNwvJMkSG8p
xFwq/GvVtkKCJELMDXbIQg/LNVCbEyNETEyATmZfxBjM4WO4OyDrExFZxJP8A2PVC/IGucs0Z2Bk
Pdsc+SAMQhYDVBZf/WvsSBJ+I7FbJ0Iaf395t0EQaxCqhTaYQNsgrJM+kHRz1jRBh7M/C870nwwf
Z5VWwECi5Jp8cYyG1XV/RTMjH/fF7PpwpHmLGDKiwbGs35V43xZ8LYO1y8avtLTbbFLbYmXt8gcC
JSSkz4rcZLMgPrONSybaNZGLFoaZrP9hYEB3VKsmTF6jGkbIVOLgjG56sYDXAoh6Y1DIvVka1Uvq
aO0SrAzJQVBOCKiYL/57UQXgfZByFqHek/6CPoAmXywvVHnRPw14Ycx3u/UE75lzKZ07AZo+rfL0
gKK+sC3U2sPduObO+qFEE/VWNik/Ynkc13FKDL5Endv8KgB9tfFuKzuHm0DOdVOacjjLAtMyDFak
+lzEhQvaPHzKiKS7aVbQBfD9MdFCy0iufEhSiVvRDKtk6MUs9dkIAkWMMaa6Hh8hQ+LnBnUtRq/0
sNrmwg1b9hkhImWBhePau0HyfT/5+XYqYUXmaV5Yv0EyQ/BQZzeOTQPLhkgUeaW4TgZvUoU2ZuRE
2zP3NdAakrIl4twTH3cKP8MEm0ECdBm11zCcAxiHyzxufW86ZDezX0rhHiFd25T1sC2QjEO9LW08
IkmhhIe2OJeCixqdchSN0LVUvu6OnyEGuJiNuyCkqawL7X9zfE3V0vzRLiA0WHjxVct4xQxt5csY
u7OmupOXzbo51mPDwaLGaFzo3ZJcRyewNANM0djRAXW/riMkJH0E0XgnUAQwDirFrTJz8NFID/vv
Xqb+G49Mu4+kJ8jnfwnrrEmZAvdR/TUYspoh7e+tq3oStR0wpnztH7D9P6VJulnlZJhdSjGiL/23
jGCE9/Cle6+TnMWqGlgruIPiGa5E2Ve32DSzjFBFdJ+pcuwjLQ3+h9qqccY/4PLw01anOqWojNHP
SRf+qzPnlg4+tugJRK4pcbLWrtmfZuQjLachyffF1qQh4w622rw4hbsSmnff8yrXYMHHEiTazegJ
ftUzp0NtWMTZdXxupQHtA4PtupQSqbKoWkLe4ufBl5H3Va3fJX0jr0wOSyObzWV51jMPXEmNaio5
1XNLhhnc4nvgWwyIe+AoTNI0t/ZgNyN8y0NEJKRXrvQGhYrbROmlzzRCOhRyoVDsadj/YYypgSKO
xKvq9cXQW6cr2BUGqOKdHOO5bIEg3uSwDrHSGRsP7PvnVdQxprepGNGYrQ9pclfp6FC6Ct3FZmZY
W+6ClTb+vVibair2R/p6WnX0O6vMUPOo2dQQC+gLBN86ho46NC9CmvW5QVEbm8wiYtHfmVKc+E27
Z1vX3XTdzCRLViTvNsovhMZR1TPyL1ZOiYBYzfolhtdeBfR0Zyz9ACubCK9BwmVUzLkedQi545bN
TmZdAPxKa0e0IDRDfJij9pGrhwTlBETPaJcJuqlKxjBV4iQiVBXGULjideLh0prx/dBoTUOSqDHf
fcxjDV6k+skLg4hmuSjhqEiM0DU7KafyjDJPSPKzFwwC4vw0/RD4cvoUMwYnVv0wOwde8tte7oa7
8x51OTdq2BUcFhvQ8DzffLOZZ/YOYrjy6Iw2Z0VY32Rmwy1SOXSx3+XPWCwhvx7GSWNm1PbGTC6k
bRv4sunUzix5Y0hIOw+pn+n6f17BihXm8y6kmuc67WWafqjvuZLBJh54yd/+9FuQiAMNW7dtCRO3
ifYZ7NObdaTiYyoJ4Sn6a32wKBfnem6r097t2F38CqEdi4lLwMqL3TpE+dleSZbkjvaWRSgp8UUQ
nCj2vuDcRvrvLHiYJxNJK2SGUsxUQhM3k5Fief3f3Lud4FNhkgjjffrGac7MSV6VCQ2RDsbn49M8
cgFUPbABnutJmGFpnTYxDnp/7LAEsClfbrRNYfhwhc5M5gPUISjq77q+vh6GzMYBReb0cuiuG6Q2
AP7q6uTKqYZMoLNz69IfUYuFMUDJKWAn0QeJI82QBZilenVSgr3cCoI2TXSO/wSs5CHPkTjjT0g6
Bjjgch8A8i+I7CWDUxMtmXRT1HzpQ/WD0g1/LUy0pOrvHyG7jwzfhk/VA8HYGW02odN4ug8urNKr
xWDvDHchu/x7r7eDmTmlD1HUiLkMJ1VUv1EDucSXicel7LXoJHbzrM4rlUnHGsyOQbkMKae02dKN
DPwvaA4WZhU0SZYPbQZ037erUpJbvO0ZXyGW9MrkzlDarqZxesvgUo1quAA+yfS6yqOhVjGdwqQq
1jNlcSWC4hqoXJBrAZcyhoalpZQj/9FsbHqa22zD9s4WFJ3Cj1I6oY7A2igxWjyNfoNi9yI7jslM
s0pQig0t6BE76H2zQN4hmf2f9/AkTsVZkRyBfqaL5mGMePO/S+rLXRrvzarfo5OAk8ZYii8gr4yj
4ZnVxH4kOvuml4AWZyJxiHdDSVUOhBdzvHKhpxqQRul7QJsArMpgPlWOirgQudmkhon96XJUK4wU
niMtoZuqc9NjmnUzkxh8AfT815LsHYlAaHnhAnT4DXihVVO+5hJskg8SRUYPoIYkXDu5lbAkPuK7
0zFppknqi99mbfcfMpfSJWPV0EcrILDp+KqHx6mzgCNfF4vzTW7BRhlIZOqcd23BtViWKY+xWKQY
t0h5erXsdya7AhNc5cHWMc/47aqrBVANK2VbvwS3YqHJqh8TsuvL4S0TNseJw9x82eGpcCoFS1R2
mg8JOW+/a8qtGZoN31BgrB4hPRjwrKBxJ10+t88afdqGuOV9GXZBz/Uj/MhaCjqAWUUXAPxishPq
kF3lOdtf+cKTHy+g6f5E6RcA8rbYYMJj/NxCiHz/lXzJPVTXFGVk6GZ+8Q2ztYIitvarebJLCrY+
Yhj5uhuAsHquBym7IN9eYygrTf5SlBWlZzqKyQ2ZLwUS2wCCI1+VvJXRzKOlMNFKaTibICJG3//8
Li2Pa7HJoETFy0xpIu3SaLzcmRoc4wwi/qQPKzR/lqcL78TJ+TK9buB8LqO3FSNWM+atBNmnRZ2/
Xbp4aPVof4oMaoCoess6zbxOz3LoJknE/5nCJ10fEBgH1y3OcpwEndEYj5ECdN8Kbqwjp+HKTOCy
sn7b8+a216JP4eus7dJnL3KrwndGxEmWhbDT6gWb6n+B9nuXLmO+E0fCbxqTbNv50UOPrVlF6qyw
vfCsaibbgy37ASQE9/Y56mkCYUXeYQdSPwGKVF4bm4yMfFqOLLPJ1DuHiGhOgB6fcWZywB9Ch/Jd
tjbp9gqGY+TSR5qt1DwZyoh77MTBLwF2L8cSZj/FhKeT5ITxxHJK0M50jmihwEQLlQwtrjxsTeWq
TKe6gmLRk0r/26BZfH5tL7dTY5I5I5mAtgSoKO/tTmPkJTmdyfwnbAgyp+IxR6gOVr9iX/n30VB3
3bQoEYZzD+C2w3hRayy7DzmSCd66DA0mh+Rfarp+1p5giBfHqTsN9jF/+ixvHHqSXFInZlV49KxH
rY9fn6jj+pEZQIr1278Tq3QNdk25NcmJD+e/Hs58EubOmrAPsfroKmU+lAfoHHhAFM3XaTSQ8Fri
AQ4Ebu07J4LfHWFBVsl43kOnti2qUTzwq5FuCDEjG1/k+NzUS8P2wqNQD00AS/A/k3lhh5LUgERS
qT+1lG2GD4PzdOdOHGl6qu9L0Vz+T5bMpC32b7QobbGVXHfvNexO8DcH9j86+RiwJKwcuwXYmy/x
//rOficUrfXRHBtJnfN2OgixI1g9chn+WTrnP9aGqiBk5Byx+0sGbHHDYl78m58vXZz6UpWWct1c
ci3glrqEQ0DrJMZw2jwbb7mm6dA8AqRSaFs1L/hZR1wErA6yN253VxTeuREej4WdUGRT4S634gWT
qm9BMfQrU3bGM4MsIYATWR949/Z/MlGprhK88eDq2vTSxYXO8C3NwqcVZ7jgHbDgyhAgyDx6TJOX
ppbzYFR9cLi+z4Qg2G2IoHu/SCPySbWzabYTGU1VJGKyCt1hVHhuzioGRrWPQUFp9v8VxpafFW8o
b6NqzFBhcPiPRo6uiTAbrQmdYYEbzUpaSXiPCAoaK38Jf4zUcfI+YYAf0ZWFbYfGNlEwDtTDb2vf
+W/HRS0zZcFAriXL3qWhnLO8fb1rDVKMEb525b/NDgLJBhTMHELi2RmaZ1YZURn6RfazHNwRbd49
I2EytM1p0AplVkkmVoDnx0f2Z1Npi6ytYr6a6Q/Iw/lTbWAMTJmXlci2pYIAdlfd9qgLsfacPLRg
QwiibWkBlBaIOhFr80/qmZO/+DorW5uJ/UA9ME20sa0UtLyOzb8ku9WvDinwUfBd/+aUTqRWdVMY
6lmb5D1QaOB0VanjIWLdSWERMLYWCe87k0wtImtmo7mnO/dWXZ/zABykAWI3mqgYH0hh2zYnfxOk
eUbNji5kMujjAZeFFn9XUTova06YtV+f9WwDmqaeOrpHW/5kyEiM/mkYpl0391D4Zow3DPMicTES
BSZx5ppZ9H69bG8GkwkbWvWYAQVm88tauNrF6/B0amI3fFD7R2rNS6G2lnKU9Wp4l8Npd4CGXsim
/QUJ6zd7aq8o3OKU36/SLPOhGIyaNFjcmmZ7JVGCXZ95SXgFAMh3vbdNSH+eMEYXZ2B2l+0YCH4m
VzUAZAq9Fk2D6S47jibyRq9Yj7qfJI6oeOnjgqSrgZ/mEhmGsP1lF8uRQK9SYnHLidTOyMjXusKV
UV+epi3JteHp2NrkrOMcgmDSUiRnMdI4hFCow5bpzIby1k/H28BQQ1mFyHzlLhYMnzGsl1tudVUL
F/MF1W5U8nwXA5H7w824W1pWfS/lXFUrnaKJAA9wIx2rRJ7ia9meTHk+9XSRNT6/gTIoNHBWZ5qj
YbnN/Owp7VC4QIkXfHPaeFBmhdD1JosPNBrJBW+8R9ARaC+14xgnE7g9z+CGGRSBpEtOBlA5bq9E
Wri4cT5mq5CDxEys1UM7Yhvej5KXEMoscCgtWGtHanOUdS9Jyqscy6psS3hJqLBiQUaGLxT1AVDN
7ZMMulYsS1CgZFVj8nSIG2yg3PaEMQTgtKIvQjU75+7aECF5aW48Bn6jpCd+HqKb0hvnL29pslcJ
+2byigRryXeoacLWRUXOZNSoGZRjcvHMVVMDKC304hFlZi9V/vNXzOGgSDKDESeiI2/xwBQ+R+j4
ZpG4jhJcsTFg3qQxo3e7iEIJWmE1Sw42YhTec1dbJkUeE8DfaZpfPVzHswcCzZ5VAaWn44jhESX1
qU8SJdFWnw3tmIqbXFLheX+lcI4MTWAj3gggQEFTkZVl1Y1QARcLU3lvJUil4gQcglD0gDkA2z5n
/1sWbxfQpM11YMhgt1oYTK3iWiSt2Rhvg+48m2ZDxAVfqeLUhg3Nj7FBMossP15EKQAT0zB3RtGF
BgTmBBXYIWs28F7DJ5uffyYJgNg1S4XZMYqa3HjDScZ1xZ9fvoWZWwou9rGBq9eO4dXqtuQsNrjy
0y/DSCpxzQtdGt8u25tYWEwWlZCNCXPWooKWjhIPdys+eY1Tf+cHKqaXAKKh0o5AZBXrCT/qhumS
GzkWJb+nGpK3gNIKXcuf3plgAHSQvE+xLrqvA0ndGagaEXkriuk567w4Ex9FseFfv3bLLRx8+F1F
l9MVxBbmIFPGyHqSTzCL+RBLOwnhQBTKMW9TM1KO1HriPRfH0bBR1U06N0JtQ5lwD25Eq0MYaBOI
1UW4yDxvLhkVLTMhjTZSo0B6NKFbyNgp1UaHWOudiSTWk1W16zjMJtyhSiwFvNSvBqPA7LeukOsl
yykdqKnSJDWnRMKHAZbHld1ng8mm8yIrw/0y67uy1ojy8EKySXzPRhcJjnD9yIExmBC8+Y0dNJAG
dVFY29rLZHHlg5Yaebq6ZSOALYZtc4K8/jOlJAzYFVnyGsTUJNtxEAVDKhtUpTxAx/Y0f0tmFPCg
JD0mHt0hx1FP94CF8mY05hRk+GiU4GabE2u3hqHjOOSsIEFhwRspjDkFHuj7EhgZZCuobNFwHApW
sUAwH55A7uMW3TzQ51jUZ4YmCHyWcR7xIlPd+avyBKaN4PoazVgBOjCqmfl4u48HfyuxjpvWgxo8
FMjMJquF0qNQ3y13TX4iY0IoxB+d+DBgODfHoPlEqR3M+p+2Y/SFP26IEWwLdWP6bQVR6uqWliqi
SRW1+9Yg40lnJYVAMKQDovJRL855i9OMn8Hk4Ho19Z5z38uIBP1UtblPwcoWjcnwKg0/cixiFKeg
OGWsoN1Igchup1schKlfEtUcZ2pPXKHe4KeLJ8joKIkMIs76W93OWB4FEwsnZVWJ5+aQAVHDdnFN
L/kuX+qQNKsb0xAaG35aA/uvLDo7AfXqiX+hZ2skl337tuaJ5PNLQ9z+2poAjjdJI0Ea0Otik50N
mVFB6yP6stuxy5Mjp5JxBrUQ2UdXXohU/paHtGduM+uPEKzmq23J54vTr/OotyGSCdnDYMFdJuzF
F0cl2eh6jmd8PAReBZdnUBfHni4nn1RqZ4pqPj+SLi9dGdZlOaYbSSy+SzT1S4O3u+HQzobOA0gZ
uQhK0dhx0gccVxLgVdBZSbE70RJH0rh38jykffFd0OxeRf5hXZQ6rXf0Qy2vfdn3eyast38zFPS5
FgFVSJ+l471rQj2Cu+UmmdLhd7T95FCmIgdysv/f3NpZgzm9ZE8BmcG4qTX7Rk3GIUtSzBdPsa7a
rj7bwKEKxf9pe45RG6vn/gssQz+9Cetijl2w0nubd9NCJ2Fhau/vI7pCdorFjK14T0REzbn0jz6/
70n+zABIxevaBBkWMTIPIi5fMQKC5DoJqP+fR2BGtXlqQsIr/BtYb4fvSsr2JbwNBWxOIJGhlEsX
v17ppf2AbmWRwn2OdphoysXaA9p2JhTM0KFyvc531RmR4d6TU7URU6bkVfwS3U5CBUwpq5XYtl3X
yrKItQ6vgkp87negRNyNzBSOYerQRWXr7+oGb94ZUoq8Uv9iVBAw+PBgzr+ln7asRBgBlXKD3E4E
/PWW62/KZHf7+PYEB//V604Py5L91+5v2A3bRiEvlvDX9m5mqK+Ws+cZQC9NuO7N07Wc6qH5pdSI
Posb7aKzvv1cjzGF9G/R/UOMfxdwNZKeIQ1fcN7PpB3aprCNfVh4/TcqPu1IkDzQCBv7q8gh3mEr
EbruQoL8d0cqxOm5wSsDqeeQoIu867lS6+Xq/MaavSE42EuLMc1d5c2+T/ivZHSxwWWjen+YFTir
zlv9IutZe4fXY2sUSA+Tsky/v7t2QT/yNRRgm3TjH15V/EzP8jVOSVbkLxlt9A3iJaGwEi8aJiqW
c2LBGOvGcAeBLsywDMZDb+jtt4uz3h3YYVhbv05/DIOFYGuVEBKtQSZ2QRqyaBdThudO1gVSXbb2
3+9U4m0jhll5gWhDq+urMZ2kJQT29Us/nw2K6VMRR1/BMOEIr8/pNoKJfA5Gi5Et2bWm9jS9FfH/
PM9YRSFTYZEHfQdcf0T2SljYYTo2f1iwen7rwm2BRrB94i5EaeGom73u1ZB5eWVFPRoM82VWSs7z
8ZTUFdfJx5e2l3NzD51Nq85np9tZ4SycCNWUz/wQ6/RFCrjH+/uTNOS2AjtqZ66+EB+uirqbOnkb
/dnwIw4m6dssyYIO1vjn8JixrytKIMRm0LubVkHbovERhF4jL43qLfVVFY+abm0yCNCZhwQjVvOe
M7W3888Bmpel18Zotu5mSR7Vdpzw/tjpJ5Z7jqsYwVW4ol2A6of1IcHz0rF/lDYxvF3zfEzJ1d6l
9zitivGZTnvIu8wrBLmoNQoXYEfp89zg/mYOvmIaKA/D/CLO7Pe8UWnSOBuoZWyIJhdpl6vVS7FQ
ovksmybfy+3VILPnLflAlklctlTUq2Ik7U933HW3ta1Gz+3JbIXt7hQKQ1TM1iaFNMstawkb26WO
9y3xAK3Lgpoo8AzMIPUIaMvsZn5Mj6858KsZrSe5PS27nozyy8TU2pcdcSjznKN1PhPBHFClTpev
D/6fTmoSwidHKHHXbHUvMbxbVymvLMJ3iL4PWUYWy3Tj7PKXkTNevhvu6Frx+lqO0qOHPxV2jcDG
uCk0ZrO0vAkfrvx8IFOi+9o2rEgZe+QlTB3tu+VpHHJKDUwOv73s0VY7w748ooxuntFqjb8ON/rG
rby1xWvduLDPRQnNhTp/mb8NyCRw4VDLZMnUCEL7I+7FzqIj9Y/QgcvniAUqVu/8LAZ2NL8akGXS
5jgBBmgDKyDhRncwMeafyAu3xILJaDcoNgeU6Y0gIJ1rStag34HxiOz1K/W27rKSjaHjsIvL8tMb
CgW9GJxr5BXY43OKfHToUH0YDaj4iv1JI6RGCZNEqeaVcwzjuDolngMrUFPYuKBvDSV5BzuVBQJN
2ATPe/gJyAQpTmetr4gKo3BWzQGE8o8IgLW8fFCM0WWXa6wf1WaxesSqpCXMo2+s8GgHmi0mcuzI
JmZtHHXByX9ivlacYlxMdEaPEP3LvYi2GdvuLEChG7KN2j61HS4qsm0cXvDioOxJdFfDBWAi8K5j
J9KdneUApYc55vQBafdZzO1BZ8HAgHovGh59rf3yIBtrZbcjzuYhrEQNEhntyb5yMKj5bItfjNyw
iMOizfz9ReMaaW5AI/1EFMFCklkD4vGo3eCG4pbwQ46uxRACFmzDX7jJYpXNoj14UEuCcZWfnAgc
ynH2yBHc0mBN9va/uSY1QjEuwLvy0WTJxyxAYUnhhCCu7XdthvfXcQzu/DeFc4qbv6Qrl9cy6yFv
r9gq6E0hsibNcayoS3IiuidZTIIow+naNJ5HRS5/eCceMGRkzpqQfL9uNoR1OCPIqFIQVUjl6qfo
yuLQkECUeo8qs6Nmxgzp4H2ygmrCzXwpsn9jiz7z+wN9x62DwEtuwNCTEvD480N5Y++hhhSYJEB+
94DmaGkyVX1cL7qG17EJ6QHhk3p3LAlI9i8P/W2vJ/eppoHAtHgBb5iFsvVR2+MY8NvQfQ0pBDS/
CkAw+p4c8v2sQRIcWwNMw+fsobY+h3g6BdcWG/wjDzBeAQx5ggwzNYgrqFWuhLER3lR+NlNejTam
8sqhprfPsu0DkDXDP3ctHV+GzVIOaCaTpxWjXZ0MGiL3Re+l192lrm4GMRYt1ggIldE2lWUKv2Qr
u6p9egukLGcLfufgGzMNRtqDBOru9SDoS7fC54V81ptmZBnUJAWDFuDmjGwES8wAsT1VIR5rqqhB
XmJC/Oz8dm8CpK7grJD0XedSgWoPhgbAxsrSBuMWAhYtub9XKMysB4wvu0AmlEjG7NKz4ceaPF5J
Xhl9eVuBocdD280uT0u1kVYkQo/IKuPwk2I40QNY1J76+ZFNESa6w7MdHrs03y4EPypvYliBszUn
SmTaktGh5vl6XTt/Ccx95xi/TOXcS+d7d81x+ZWFIv4yNZURq1XSvHT70VASfGSTO1cWES9uU+VG
GNNIpr9uDeEGHuin2ya17aUHNAQ75OvwJvtKB7lXtmEWV4jbXBr5hMdWMfrGMwwvnO+6N/D/6R70
geuqaJbJ3Vpj60iqkL0gYXNBEIFt8jDztUV2erLOgV8R6UGDpBwju/yEd4Gnn/AdFagU6rNEMdSg
PCEDFfB/c76Oa8LnH7dUvOywz1QffUKmoSq3WLbMdUpzSyhJ1zwqpovIfC8efiTfjqNoVGcz0XWz
CUds7o5LQNZrhGfqBiRMxCqDJlZ4CSavNjdDNnL8DrWNZVsNM4FPRfrjFScKBz1mEo6SwlFPQvvb
GbAgwuZMHgBwIhYHcS2hAVqewUcC9+016PIXHgSNdlF/VKRUIj3KL4hDcHotRh8AxlMfqGRj1ot1
ziIHlvN9qA/+5Y4hG+QKTLMspUKXDvh6KxsNhQjvpyf0nhBG3WqeNtE+iYZUneMTP4onoNm+70fu
mnWkOPkEOICVyrAcwH9Zub8aXKCigRFXoRAyepnSFR5q2NGKUdyN2UtNwy1Mfjc37P0zpKGKSw0W
6p0rPpCBMxTqywQ24X0bIrR7fAo7EP/4m0bLcUvbeR2VpKsINw9o+8BYE83wBHMXjCiZbM/eLUq1
0UwDiW5DKqwIBh6AvCUFfEBjPSrrvj6WKJZ+JxMvZ7n89QtdRnLoJB57vGrn1Dzje7YjFFAfnE8a
NuWyuJo0V+TC50na4G/gFw88Ehn+mZ8ZfcB7Rx1i+uQ6E8WFzQGC5SvlZiAusPFaC0l8QfBtm5Ih
4kvOFX7ujIliqdFdXH3TcE7P/wQNmM97tcGAvAMosL8vtHj5DuBUaC+Dw2p8ffBB+uk+qrQskIZw
hyElHBxp4PIxvMgHN3G4Roi/ZU2fcmvcsB8SWjbdzxnlH0FJXguX+UgweffHqFEWpcpj3ZIN3Z3w
g22FR5TNwpIvXwLGg92PjsNr5Linibk0bTm4nGiZNaAEEYxR4AgGykkOHE+NNjiPzdZ8kjUa/waK
7R4m0lT5NMTAQzWyc/2VYLWVnoDwHPFsOPpF0JVz0PXvjs0fGDbkHj67LTe+2g1uNtbhdF4qCE7Z
U65sBZqsvNlhgrnjj6Mwp44G5fBZO8fMl5g9HCFboVSOyJbtgA9hyth/OIBbXiRnEhP0t81VwoAj
IXeNc607WxxCX0xJp7vrFCPQO9CYFBCaZa59WFutxll/Bb8Otk2/RERNZrr8Byv/86FVmuI5Ux1C
0xZRe+/WJK3+xJsKkhTK1LNzQ/uzDSs+PGygWDZfszkHCT1xm7qll5prHT5zpg18DYAdoMnnNBLz
Yk40c1avEcJFJMWi5n3ACfsP54ILE4RF8DCkmtGcydc2c9XhZxLurxtuKF4VzVzlcWbKu22Ta3+N
8n29FtqsH0wW0B1/4ay5/ztd3fe0MHmWcH+qh2i5pV/QtQJq9QutDjQztl0BbjtOoXbC0eTtZEUe
fYkJSuDxmhfjQ8Wk9GtZHNMIqD0MdfkIIwIV7AdGU5Sk4skPNzUM7TfRyIKk3JjK3RK15u8wmRJH
AlnBvekBZnLdpU8jRsqPRY8VTwBEkP2OJFLn0BNAnifK1S3uAKiTY5ejx8ejSXvsxy6u7xt4voR6
nfZKM6iV4/QW4cVXTPxr2ZxlmYoqPUC33T8KnNl7klACAVtieQk9HDoq+ivb9qufKnqw7X/qZkdn
MGpC08wvdWE3lcRKlbMJQp8KFfX1Coml2ioFD7lwx1nY1LGCiNh43LjX8A8/SAzS4yJVN7Uui1eV
fkvZHtqv4n7plwIoiDQPQj8WJzPdELdpaSSp4hpvRTO7D6r0I13w+7i2O9HPJx7UZeZxA3cfZGmw
/k7xwcXn5+AuNLPUkc4U2of2MIP9C5UmSqCcP5qQ0Eefno+vpZAzoVcV5WbscFZreAKDBTxAMsL3
dhdI4bb+fKW48yvPpsnKktdAzlVs9aZ3ZWu9n5oW930yTsJx/c8yiSj1ztMKU93d4mTgRGrPtsn6
tB6X36qBb6z5ZKZXTBm5OuJDJMwfEUNSL8R0e5XXTuDNaxI8pYD/HJfbIZ7BWOnQmyRLYRn56y2O
U0+t66Y92JTB8Eig0tyiPBBrhgydCRJjeHH8B9ELaj7DE0gVMo0JKFpmXMAjKyDYTScQSjUxbrOJ
ipl9mpRCzHg2Cn1jG3R8K67kXexkwmO0KgbAXrPCF6hvrDha4btQk6/wvERG/bZzudkhMKGXjvom
lclf8StlTvOwUm8Spk5NlE8f/Twe11dGFGLdhVQS6i3hZY4Vbpx1yB0ErwNvvTxIDgxx/wAu1mhr
a3+0gwbu8Y2JtBwzIq0L4JtNhn6Y4z0cSiuUflNb78dWqJZXlFAkiSrg81/gubQigXTFaYsw5xx6
Xo1S2mt+0kgvN1hXDgnR7yopARETXbLUK6uMZGO7QlBp6N5o8bYBl1SvavvPwD2n8mMYjAdDlxvZ
y3Qpdqs1uPiuGRrf0NOircpORkLb/793QjYCbUMYJxbJ1+I4lOSQJfkSc9M7OM/5U0hw5KCMQTF8
34tWsOirP9DR1xO0i/NnYdATvVTMOiK2Itvz7/KLJtCSUbgT0Hu5eD4PVbAbHMiQTnIZKQ9sjeJY
krjQg6XUo3VbPg3jE+W8+2nIXI1SgBBEURRkclX7lOyIZEr1E6pJTTiJe5bI7V8LFD7qNppDPCT0
KW2p8C8F6f8QD+9cNaO8p8Ds+ggzIOnDEDOtHB+gY7bINX+0DqbovZ5iTfD7gkPdeicK20mYACeX
2rgIxKCN0gZkYHZudzUcQ4sowB6hy0FeQ1RuezWS3AFWM91BFSivWhDwJQmDj+u4LcxIyxWeSZ0r
30kJdqbeQzWaj8ayhBlOf6iYywrPdZTOJoj0/vJ+lXqnJ7KPVI2dqa9xkCqqmYkqmaTDo7b9/pTz
/ZOaDtus0F2vugd7Tn5vxSQigEH55fR0O80fKu55HnVOtuTsM109ZvXbFPXpReagzc3Ez4rsODme
ZMl8QQmrrXzR98/f88/PHSRz/r21HBxZufN1VYusE/HHS5mOXoChb2Y5YjT9Se9iJQoKS1xnxL+P
gFVAKM2ZQD+s3purHAvzP9n+J582xvG7mAZasCCZAZmvZx1ctBCqEjGtjxY8I/lODdufAgkdRTK9
Yxee0Ykaz1WLa3gcSr25kSOhzWts/93/Ns3SIU4A8LegGr2tDXCSkEpw2TXcn6NnNpFAAYGYc+JS
83DB9Lg7sRir1Ms1OoLH4v8CaROy2X60EtczCmMwqRclWz05pkvSt0n3AQrY3c/nxbutjWDz8DRA
2kacyCcPkB7k6CfFeTsvwxTbZGuszYqEanseWpV/cfagkrd1lMgTdBGyzu+Xhg9lyIIfBC6XXCwW
KLKRSWmTaCqguo1e2bC51a99muWo1AJ6hjgeHskzxHMeOObpitADYhzyy5YzYUre3u5vJeRbKhYv
jJjg4opj9+V+YNd16E/opoSmyigIBGJ8sn6qiBxUj/o8jXWcrGSRC5cOLj68j3p6OaqGCdUwihzh
RZXGHsn9NReboI3UL4PLPTkYx1wRpP4E3xjEhD7jZESMno5lBcIU+PU1kFp4EJpzEVSI22tMKO2V
KG+DLhCs4JH35OrMedsoueBhnbZYWFBVCYq0VO/3emsJruoGtvlUQT1y98/ZeDT5wr3A3QILRwqa
PWK7JoqLhD/qJ0BINVo86r4Em3eD10YgDPwuwFA8fEL2Zs3oirJEJX73wBrY7DI70FIYgxe6PBTA
+g/7iebJMYoqi5SyuF5soNIX3x02uu5uuxdqIG2dYTeVn/KSW4xnrAsAMMXpUSITl8LD8cktsGjh
GweCSKVpFVAOds6XgoSviTNQB8p+zZOSgrRnd0NC1Ls1E6Z7thOtS97EV6R8VZP3JvTbw8Fy1eaa
plHALOEmbG7e2PKmVOlQFareGb+zluLRsRspPQfuZD4zgZWUlQPzI9Sra29fJ/50wnWnYyrUSi59
oas5t8lO6sxZ/Lm3d81JkWwWr8dwQjDcpo8MEfAoIAg6+qDMN8uNqUdW6gdfBkAw81mitF24cEsI
jZhQHTSRi380omas4LvQ+yz4PJJNTwLkVcTADIfRpA3qBAJEOVd1Ukxo+2O959GA2JFAhj9y+Nsx
ZHjLyfMx+IqyBdsxxC5JI4FuTOL73ybgpXrmnyVvW/XU/LvmXBNdph226MCV0OXEkDtUyDXS0kyq
8Ayu1O+z1YOvGRdrsIpH6JD8uq+OZFkvC+PBCMrmSNYlN8Sp1iQFHXT2ZlrS90D35wqb4AuUaQA/
aDl80jC4uv4V0ZmvML63DpJ54ZpAAxMraU2bBPAM5lwKInmLkurbvm+mKlB5p3sunBK31Jl61jQ4
fX3L9kjmVazTweOzgpdm/LofeFij58tFLI+Gn6A2CSsE7s7VcO+9gRyrsWRLKe08o7jldkHYIgeg
kw/BrDzsZ3oP1a4Wy9/IEm6mIKsuCUHvMVhRPhmeiSeFqCsB45FnU/+rPbO6S6tu2uVIRvbE75EH
GQ7IROlIG4GG3uI55mNUKpgeWq6hP7I4yKdFOybxE5IUqJpjkO5j2gRCrMFsUUWS3D07RK9/DcCc
DyuT8/pqSv67x6yeofNK9iphF787EVGcJLYW+4NnWV2zCkdJEt+9LOIS45oLR/h1b4bkZS6cotju
gyk90TP7zn6xz+/gOQ60IfGcSJtd2jsMyiufPHoLsLIuT+sqOISMWdo8dfyHr+MHU/mxaQYGeRVc
fXsHrkwH+CWTQBj0xFeEPkfe1oA7G95dsTUW8yYeXn2wti3xeMszpFGqtBdxY8QsABQynjYdIlEJ
dS/DngANN+fagc6Y1Swl1DmJEb9ZqAqcKeP7ZkuhMAVqiD1mjcu9nmS0MbHShxw3fml1hoZ8Xv76
DM3W0Q0pw66lvNXTukUTz+jk5UipfM216KD8dqGi9dIZMyp0k87lhv833oXNkph9zYq8K+WcEqUj
j8wCO42Aez+In4y+A6/1MVW2EEuxdIMRXTAoqt/GVw+owzlgeDN+guo6kODmJssZQEdvGMfVFGDj
ADmx86W5JDToBy4mawzTx4CTfraOWS0VNmyhnye+E+4ZilnnaS7u2xajBjoRcfNWUsscqKO71zRt
FI7O4GSZez6ZP1egD3rCfH5ADhF5ncSE5NijlW94sbnoDRNOFFxw3xY2qK5+fUafldBJImCQ5uYn
CxEYumUp1Hq5IKd0xG3VvKjzOU2xhGr6NuDC+9R5TT7cG+kwG8WlQoxm/wgLuphfZ9mHGkCquUco
pKzeJbrVTVqwqpyFGJIGaFk6Ee/qoVbJ/BI99csVMmxFyzNVgLhEM6jv5TVswnvPopeTf9FMQAvn
JnnCD52B3xItJl4n1Mh7aDHCZ1cospN2EqzwfL0v4BkqtHrr8LOGpXi0bmDA/MKY7YK6Mcs5akT3
3HDEPIBuVhjF5jleNF6aQ4cMglkUDg4JsiqaZxGo8Or+u7oawY2pmJK/iDASgSBJILQ4jmGpkg93
GFAVF+0b3fF2gXf9o0FFKI4O80JS3jNgqPOTuiuvWuM6ZFSZ50/Tel3HeLQ4EA4Gko/KbHiXfH/1
2krvqDP2rwgrt9VCbXND+lhKzhtWFAfQvDp1CGuEkRo70yFn5qBKlfMXaJS76WMtWAl0l2KZkmGI
V++pkA6GS3UCp670+AtsaoQeTVLaeaF4+EoDAHTN7Nr3waarTIHXnpbgeTOUEB/746Kwk3RUh1yC
vPUbRup5KHBNyNR4gr+ym1Myv/2aBqTNusrEmPUr6PSHdaUijZUX3hxQFLV6tJ2f8A+wWqmjn9H0
b1izPb+LlCIitHGerknBddbXS4F2HbR2DJCZeEwPNQi1Cik2YeMzN757PfmKZ1x5cxl+vkugao66
48sewKd0VBFI7FutUMjPNNr5XPMQDzRXX2MvFFPxONa53jyesQw2a7WgzZPCrsbIrikgpiGRhO8d
kkbkr4Bk4BbqPv8L9/ixOp8Tq+hOr4vbPDVInYx6CPEdJW6H1WfHdwGDuWD9EjOlpf6kmuQ/co+B
z+6uh/u6TNFaZuCxfAPqDr8wD3cJ68cwaRWuX81cnjnc0qV5uBlDJnu+wsTdNaOQArbJO7jurze0
zhEr/5apV30Rha8C6p1o2LAnYQ00WVD1UeM8VLPfk2UwejMB9K+K+bha0twVO+By4mI9HotGEuKf
hDxppMzfPCcWXTZG6dTfbyF8fw36v1U1h75U9NqDuw7tfy9+N8ribUDaPZCAOwhpoL61V7PdJabj
pINWC1RGawYA8c2L6ENQMl8O6mfMw4n47NGQRq9rs8gp8QSbvldJGWxms9dpuiyqMYP74sMrEpxp
3DkzjBhpyLNclHnJSkehgIMGMrU/rJvrLOCaSQzfnrNGSMYNmEiGdmR7G+mMOVlWP9u8+CsKKfft
UgHdgOJYTO/us3feA2mtYdlsYEPSQNAq0dIbD8WJ2cw4h0F/SX1nwhg21tdW4gT7Pjczdx6DIRAo
XAHRD9pXAagxmmrpwI1sABVUiXYX/tsSXS0rKoTNep6YBDLXhhLO4Zuj7E82jZi0jiYyFRNPzx9y
27y5iob3Kh7mrrP2wK5q7BbMpNM3hsFKwqnG+xmec22U0PI0KvZOepZOJqcsix2SyR9Tp+rF6odP
0VvGF0q+c/3NffAs6EtJKzmV/DKzMg9KjNm/1bp5DvM1dkhoF0imgvNCUTJGqS1zBmFAStP3yP8j
EfdZjugECNLaC6O86qMgMP1/19aXllBWY6K4Z+bjewXcdh5dm3GvMdOU5ZN4V+T3cXx0j/SkrLtY
GX///ZM0+mBnBuQw/l3qk4ysu39fuJ84ojj+rOZawaS/x2zcpzw3uDQJu0i725DaNCHWZTVlzvrO
qvMZ5aEqlVScOprUnkxUmX0wMMPmABn1EXPvQXoUOpBjpuQfc0oxgsMzCCQakxxW0XByzH8sROY7
MOROwN4HAP90bLuLov/V/92gPNUIvgLz0Mr4ULsGEgcfNMoS+1+sXY8Tc+rmb1RnMbKEO/hZo5i7
NRe3fE9QbilHvXBeAD+36mk906jGUEtCl3Sv/2KTNW5LDF+VaT/0DOwjcAHxknQiI7kz9+oMDd+e
X2WZxKF+M+9s+IV+QgoIP4DYlV+5/tHI45+HEmKguSwNAg5OZcSxOZax+/Y61Rf6FEfCjnXzFHt6
Axkyri3vIOb5B2fZmyZI10CXaKTReX8c5M9jhZLyHhWTjvyzRI3b3kDy8JNx2PmP/udZEmo2XwJE
FpbQ0CEoKsz0erig1E8+3z5iQIux8BOiz3695DAi6XNXEo0Qt5o8x4EbVbj93kbU+Sl3jfPJSXdo
RCCdA6WneDZ+ovKjv8hLh6B/IOwtY51B9rE5grzKNDEPWhGgGqnR4FYOML5KKXhXQE8KTwrai4oS
nppQiPqXo028Tto9dm9jMJMdWb9abSPilK+fpGpCGS3eWI7tukakOWiF4K/cHu+HAl9mehcR/ih5
sQH4qIxrzrqTiDdi37xC7tNZTxqQJVVP7P+MZzIlTRxir9d079LhJ0Rr0i2ojASiYJ1BpKLJ6W7u
svEaycRia1g7LKeu6ID2rVXR0HmCq89NvRFJgDy2H3+BPmqc56X3mi53erxXjvmzSRcgPHtYX2a5
MRYxRgrV0YBPDLRrv9M4v3fwm+HsGuyuzZtNpFhGlx6HriMiqSs080w1qnPxFT0U5x0wsjg+x86L
S8F4ZV6c3oSliVITeXruoz/FU+tv+bwAC9LXriBj2A0rQ3KyofhNS1EM2HVtw/sJvCV9052vIbrm
bkXWWhWFMgvBl/B41myTYjvZAODoX1zFLLiBQDZc8j0Vbk7qAbGVz5+ldIMzlWQo+HBkyNT1Iwf4
xAA17cWGyuSnMEd4z5U7fA33Wb/K+cuzVyO2LIpWveOhzAoN3oYb2599P0/tvZuQCVnf1psPcDgY
iAKOplIj/8JB+cquusK/Q9CCziIiCwhQTr0QAOoGi91bpvnM+cxyIhuq4iUCdrspb6/RKIPMR8fn
vn+nGgzcUbzZ+zutCGajf1Kz9OEUdyQy3d0w9nrIQnx6bqiZj7j0FVHZkMYRPUTRoN5bJerXUn7B
RNq8xyBOGsPIM98hNnTrZTrAHRRbF8szGOwtUPvMhOH2OS2Zsx7y5Ucjdxsy4qgH2UO2em4gJcpr
QsBtmao3M9MfN5sivn2DL9AaYYwgeKkiPE6nMvBtaySJ1N++3cbnDdL1IDgoD/G1EGdOzb1xxcWQ
cYc2EzVOj7AJNkAiEvMIoKd5hILh36c9wtw/vs87NYCwWITwPb3S0WtmQWhD7d/QMC5/SUPWSQsu
hH38PjFCK3+WgJ0dHg6wpae2r4WstxHo6x5P+R85DjALmFqtp+aCc/UIj4flvB+NaZpG/f2++d0/
T4r+pfZq5kBIIiJPE34U9nSywlIXJEKhIa7Dz56aOaDELThm77BYjL549wSUni01DJ4WHN3ZKM3Z
59t22KcfOeqs2dNDWRrOnJqMoayXz8rBZ6AAtoKcRcCxfcgQFBargRgxSWMejar7Ia00yl+TK6Nq
Mm75GU21qCJPTHlf/KnhzYCmxS8OV/9WkFIB4nAPaBQdFTL2ADbHjAv/d8AyfZFDINv/0UdNJmuI
jdd+NywItvCbU1mLHWCVcbaxAuLETuY5Ba6qxHoqA3qC8vuz3Q371z6IpXSRAztVyBKGX6CV3l5L
u7PyM8sHLILD/vYRxEwEWXZ4VNfwjAwXU8FmVNbmfXcMRvJMypzN/aqnnmfGhLH5o5Jb8g9ZMuDY
G7XbEOSevcFhahjPgrx44+LH8OJIMGGGeIohhIsfyLpB13w7ZLB2D/LSXcviZZlPR/lTSAFHSIf/
rI1iyK2j8ieYg7eiDa5ieuN5QOjluflG7+g44ayT2a6kIMNYWxb/AlFPkD7hLSvDhclYp0ALzA0R
0LGwPcgAlnJ+krsTLZuiJQS8WrasP8rIfhH9tnMsB1jD3nNszuwYLmyfk5ondOWfHRF2Tfu+0/r7
L6WMCHdBQ1BJwiInKbxalSbXsnf8KrNnqWJJlarbXplYID9xaSi0xZwkwjA6AazZnyepq6XBL3Jv
IYXyjg+f32gmjmIA2YEMLXjf2Z92UiVkU3CLE+NJ5bi04VR5MdrNx7Pf2Bu0C9H4KBjeRGMA9vtb
4jwxqBPvyYs/cUyUbQ53qU2zqSG6ln4i12akiai8kasPawDNQ++QzVlTRC+S7skkL79f15noTsuQ
hZ8Qjv7O4b45yAfEJqlhvLoHR4W7gJNPehpHQjBwYSTZJqHSPUDOfGV7uiMN2rsCbmsNrFmefXWY
8yOK/lgzcwyfTpTgM9V+UZd3Unf5pH8wN2WtIHaHGtRjdoxzJeAKxznNCfOETNAEmer2L5Dd/Gb9
8pafD+FWYXO3m03I4LKhRRXwJ5US5RuHSzDOndNjiznhZN8511vA3nmm+stXwMDpkKmEB3gcE1wL
AyABjxDj2171fWoxtYt761Iw96Q1JhOeBUyQNi8GecfIBJ25xgL5aT+l0n93be3/zWlLFsRztPS6
ixHsZTZVN8wzxjsFMpzZxZ2ccsk0kzM7qVTsjEwrj5fGmisi0iOzcxirRku3rf3qI/l9XNZ/s55t
Rfp/d8XdLCu2Qj6Xcer4WPizbIcyWGEuB5ZRU3hhILRPjl7OEpyBZMuPLsvO/DDp+tMUigYwVRfQ
dXcnss8nrhrjvS9TL3VTQ1PrDTfOgNxE3cuBpC2BOfVcnO3Uhqf5sc/7LTfZOVFw8t4AsA6pAT90
mDJjCUbVhLeqPg8q4sqD6tS978PL5ySj7mVS9hZjEECik5XSWH98Qunsvuybtcn83ECgN9EExaue
KstWrAtNZpB0Df93gM8lPJDfUwoutHq+9f6iS67Wy+MRxadpniQ6S8axSsBvRECsc2+LMkkf8jee
DHJ8bEH5oS13CmpPuAkEnnxd3pR5h522uStNbBNBx+ESR7+orX4quIJK9EOtkepdtylMkyhbSuoH
rZsa2WrATHZK9tRMURLWqODrACHbOEJxPkw7MWC65fOlBZ5BjgoeR3JNMymYx6PExJgIxuGG+tRI
+h7YIGICFaB3GtbaI1atfuz9+Ogw5AP2j4sFMGAFUDJq4kqTRc7h/t2UWY+CRY3aMG06DapJ+s0f
eH0aB2jfLGsZhmgD+5T42Fx0NpcH0erK8nhDz9E6ibkz+5ikKPXZhi/BxN0tv8z8UdVOvZkkcH//
CLXSRcf6zJiVoMLKJC6qlvQo5VN3yCz5FQPbGcwNbUum4kenoRWv4UD+sKqTKzfSIBTY3Jv/oEH+
RVzJ5bu/2Qy4xXb8mXgnW5UyTa4OuiNyWKaHQ+F58hZRij8a8CyxvEuxJ3QLJYvRevlKZznhzB6i
T4zKU6DPq889+QoLWb5XsJQoFbFTa2plLATLwJH+lf5AKXKulTG95cXeHCMonrvGomWTs0ZqEG8w
UBfb9OXH/1NxjbHNLO/yfJM4AR53Oy1GM5qjG6je+RQJBXnSKmiMa6geNP9NhVr/CmucbYmsg8Dr
K5Q+cDmYeCfjdO0CNgyMs39NS8myzaFWgFaOxWF/CvbkTdnJjozAxDkPE+QHimdn6a+mUkqT1s6h
OQ/YcYywChtfs8/R3pHGQ6jQWub7SY5Zo5vD4aKdbKqiM3lMqIHNJKt+imaRStrCDMr1rxzk9lJG
vKHziNKkHtBoMezR/qNJnp1a+DAfG5pCgxS7evRIVtQ71na/ZoEwjROQ7qqiaL7/x3hvJRvqgnL0
UkM/l+wRTaSIb6aEyXG4G53lrFrobIhldV4iRHetqXrVGmuE802q9LyBBFkSuT9+79KfJ+iPEI1x
yxfMtv5RrRc7CSpPv4T8te9LlDuz9NVDR5ojUsPPUhpfLCc1H5Pt0hcrVMwtxovEp3Xhw/72Rriv
YWsapqPQiTSdEt2bB8pWbU9/FQ1ZH+vvMVa66GkStdYTBr0HTDnFkpwP3WkS4bvOCACANlChsi8K
08r9HjdTHCofRrUfs241ykfaydqTwAk+vrBVHJyLkkwAJxWqfLe0ygtvYmzfigxuA49LQNzfdmZ4
+WFaQf3jogXurzVcf5N+zO5kUFa7VYA3SqI1/M/3C09zOdFvzcasdAYFLxlAT+G2SpnYwa7WPFlS
oSFnFi/E6cfHhKGk5krFrVWTrDnJ0mkKgX9rodt15EMjMMPlx66lBMV4tRqKkN5XGgL1Ofj29E4Z
Y71J+dZUzBig3I1NKAAUUaMT+IieUTSgDupqxr6dqSyaOLQro6c0LeeLZhb4SpA2RRSsRN4rxR3g
l9yHT4oLFsNvxi/G0k2qhIN4/ST8O/9F4eOVpZ+csx116ZdnugjgyLqKiu7/HlX1RI5tXBQnkJ7f
+wbOOBS/s5KGb/RycI+x096UAyYd1GGNEQh9nDcFNrZvZTM4Y9i/2ukRpunXC+mXrdUbTgjvZXty
/x6TrkVSUnqs6WH3eolo+ny7V6YWIoUfyqlmaI1qcFv59hHdGOosOwQuIhkbbAvjqZumTV5irKOs
CwwZnLyNNzvn7xNmbTBSq30cyjs8OHKhNOvBd0iLWQwKfNlgqXd8qlwjONKUrh6eXHGHXmhHxkQE
hjOvhiUo+RwMyNUAHfcdSvsMwIivL3ODqaOUSM9OxrKGebiXB46VHEGuBzEzJcI7qvDCtZKf6kLx
udT64jgcd8oMCfIG+exmNkNha8zjANsJpMVJhY0gF9ZhhtZ8rG+kbuoUC56EyQybWV/Y9ZxjNXNk
RHlFNKHcspSXvTVT0BY4oqHiLR1nqarLO86s3T6ndSMiQnpvpMYymC2RnCZ6Sp0rW5MUSk6L3vAn
XobellbsF3CDdoPjWM1Ip+iawzg0x4ugjPMsiWyCIrR8TfHAOGyhvSbpTIqbF1t9eM0Mj7mYatd2
4YmVIIwTt/rnjPdRnsepRr9Zp2MuNw1WXkBt9oxzjvI6iIozPoJwP1FivHrBQzQJyM4mxtqcD89w
2o6LAnlKzr4BZBP4TFowd38x6GW2R5qVjf938OKmSmW4oD8MwBvO5ptRJwKqpWPCTL/F8MhaIcFV
10/PIPL7QkC0We6wGTFaXGaq9XM/WZNE+CLiLgylsQZfWnRxI1NTy0ODr/OjQM7U/Mjc/O2ktR7V
xj9ni11G8IIqO9uag9KQrpKi+7RBEAjsqEtZtgHBM3MoYkwSxRokeAVH6mCWNVlweOqzrm35OisB
HxxtVB3/mJOyO7PbLn2i/AhsLJEN6wsPaRNJmOz2QqQiVStfAYkvZLXH57iSy0To1g0/dllOpark
dP92igBQtt6ny2o5fTddHDc7cohOszCUXdhQQfhGj4qjzjgJULVqa0sX0chQb6CjH7Uf8udil88h
/JkIvGkL2/bUGOFhmeOpd2dTfTu16+9M/mn3uVr66pMNnUeFtDkp4dx43TmM6u0FT8kw0h2ZWsZY
5O3N8r6qIIuWhSDZrOsvhJW7x8OeON0EQDbsm6sicBtfL1p9tNzrAaUj/Sm1T25l+Vnc8srIPiEA
GYJzDBJ+yamULzVxSGABIhi2+1hR1mG33PM4wbxFYpa8bvevs6fn6MVVOJ4xXdTMvQjr89PvG4VU
4d1NrYPNQdRhvKZ8Yruo9Y1YTS67yKxo8gwHaI5/fr+znkWNsDzuNSIFWsPDEPxapLPvjCWaO8X5
wvDPCyca6NcxZJDPDT1TO2c7+WQ9UKWPvtKf6SayF0/NQMl0oFUeIrjO1zNbAxGeprGuUsSi1cWj
tMV3KchLuLrOclJGYUJZoYWgaGgBJfyr0Vw8KtQK3+yFok4Mtko5bu0L/DqFKeGF3+oKJ4Wd7dry
gyjNJ1PLqsc8eSMS/GZvZ+S78mLMQdd8GrhwzDMh1vMojXXR5l0NbzGxvsrk5QzxA2FZf1VpRhrr
Mm3SoURBydXM5oEX09TvrRoJ+g/vWfOtdevM/NrzOkuf8Wh2hYXutTIwjP8SEngn8I0eOBuWrNgI
rSQiXEV4Uwoi8hTiDjYTBgHTKhn7BWiBt52go+dlVSZSMytzeKfT4ghNjirGQgQj8pGMqCoaYWz/
fLr7Vr5UfCnpCKHOa+/2JVMZ4m3zVGJPtpYQab9UGbdOeZV0AGe9Hn10MKEqzCwZ3ZO8cbU/dfcP
KObOln51O2vHLZIddIYQ/ox2U1qZoTteTm/KgFaSC/TC9t19+Bs+GqSMVttXBgwdf/cau98BHNCZ
z5RfiKeky+/Dw3y9/2Bf4iaNr02KeT0sG2+PNsRZT30mHmKaZ/JUzJjmROJPbnjVXEmF4LHLKvUp
YN/tdvrSaqaTSTe/NVUCZKWaaNqXjqa2C6koCmdcFj/BRUoqUClbdwKqUIRJcBNCoHlBWvqf/QyK
igHIG9t91wsYllQ6DOAtJD54jiv3j2K6C3U37X8ZHiRNpD8ffQMgt71UZggyntufBQ/73ZCrO3ix
aAcOdHtr1DPp2XoWNq3LDOTMxUh/EktMNe5gj1vam6DnXwuM5T4ZPWPdcWBTCYOiOFoE2sFSfYF7
FDGriwOdJr4yk+7al8gtaPBGkkjE9XVNJpb6jnHeHt92iCcCh3gBw8i+vU/kP0BO3rLrgepAHY5r
w7fB4fW2R0jxvnA378yVkANpz4kAvWsrpDbT8fmc70qM60U6U8aNHXtJkJwroP7/7IgtHRUDQWyI
ICbP9L71vh+LwQO6tz3wRGWOBpAQ5WcLyA1cjtQ5Vh24uIsb2DOWCV0FmhoB7abwbO9EznUoaN+L
8zjB4wxTLLoF6ANEVcrwnKG2hU1DXGzX5q5/SR+lOC9q6P+rzNNRaCo4Kw3bDBOepB2Lx2r8aHvi
qQhF/5PVG18TH+64b1pdi3Ix3/+lYyNM1hESfFuJ0+LUcImMbqICYmPOVPsc9UMFVNThCZ9IDryH
ieKXLKkRYGP0fyC+9XjpSH8nSmv/8TEnweM6gDU5r3tQxibFK2V/MYL5URPM+jZkWJ6LsQUzJ2/d
GdmolhUCHNhJRu86hfxcu8IaeHeK4jtmR9LnL1sO9Qh0EK/ii/wwTBHKUpUIQNOMQhC3NnFHuHP7
pUfJo1oMrSkiv7uPPOVH8YQUPD54rVvRdMYxJryQIAJPWul1WHyRfcTGTlJ8W/e+vCg/KN8Tlt2y
tEx+vzDwAxBMB1J2LZL1LDrTPUYNaGWhyxYhP48nROs+3WHiTIFw8b2d+iZUQvLVxX4CgOWffdiY
s2GoCfnlkEwmNTHOQxlP3FpegzhXRq3pU9RRrIiguiGAESRWUXp3cqknZMyFwKZw0QasWgj4eiKJ
Xy/qeqnmDuWt+MWUA0QpexsaDIkKPEBFHPCTGU43xZqjayrjGrc2VNbfrnF2l2j6+N45CE7rxamC
sdsvDV8hJBmBj4GFeF77O5swzZOxJSBIwa1W5KEyDqDVAVJgHbefKxwEoH42GEKYWDDDAuw5/dDk
IGH/kDJSlRpG6ZKao9oWtdgVBVTVZGXmUMCXxUcwd0sbUq0lrJvLfH+OrwC7nUZTszG2KH+k9zrp
pK7QEHCRWA52dMxXVPWUJZZL1oIrL6vZ8pkoZ3Huy6u9KcPDtsICDY0dN51bqsyma3b969bPJJVj
sP5bcyM4L/Z/vvQLohEgk5J0Ng8Tobuju9kcHgqDMxbIP3SF/nPaMQJjVHGsJOFtXKAtaNq5ufUs
gw/+M7IILkxjIdNxYwd4hcpKGIMwC7SPRV1D83pRRiwjM0dDcyy4VTJMBPzThWsBYbSJ9Iiep2L1
eAZXVjx7GUM4/ToC6vQWBWe82W/JanFvHQhZU39sCOfTuwXEtrBJBjw9dLbZz3p3uIaEGTKM112c
EfUVjozRfDb/LLjkRPPxuEyjOJDY525gX597EGBwx+h/e9NmJOeCSqjqTfHh78wx9p7CWlHjSyRY
YqvTUW3vzuZ+PyNkZZVOoZvlxsMH2unFnwxi09Rn+7vJgWjTyFYD0RP9TzfwTNna1PlPTXCdWN9y
fvT4wOPMAo85q6MGYQqFv+q25B4soI/KVO0K7PRX6HOnkHdC09JHVAEIik9KghOau5tq04wgBzPU
OJ+RM4a2LnM1e9QL5PqUaWDaHVXjnOG/uWhuYbaoqGgnDtkFqXAvc2xeOu7UE+sD1CDsRp5Cda1c
jC95GxufWPnFBHoh++gwjbBJse+lNVal3gRpIoFZT3289pK9LUVBOLK/URkw7LYed6Z438r/CKE0
yG+XI7jIOzP5EH8TbC/fbJmeF0UReIJuECw8dNbrt703wzRcmEobUmXQTDyYCybQh1rHWRq0w7+x
kFTHGNXd8LbVhSkIt4nn2RI2Lr8WYK9A0WM7v3NEVoXcea+ESCl2h8ZGUJkQD4nSRqTahm4GK2R4
2G7qZV9godewzPX3O0azKY0NLQhBvBqdwrpZwKwEd6oAa9nV3JQHw6e/X+q7oSIdYVCylyG3BxCL
GlJSbLgJJ3yRIih6vbJt5+JwRNmgxK79oX3emwR3gAaQJatygzUkkqxvpe1flivxzHUio9Bt6WE6
3ltYDgMhuJjo16PQKkljC7uDox/mgdK+tav9Xaqv8Dj1KuC+XxgPvLofQs5d8QbYtXLGLTxTWK7H
nDOaMxE+ti7wqCk0/ngeOFfNy1ib3JT8oIOn63RrgIXSHaG5c5caQ7mf9Lzij/dHlOg6Sazcl18y
nkidbrEY9xn1JJpjKRonxvKPVL95kGCcINUlRnpL7mlSuu2XgHGuYP6RBWsFEOrUvvreJelFBYNz
59L0jdj1lWPISichrszckMQA/gf5ugsgR4M1K95JGn2LPqT7AykLMPJ7beL2/yyr3VJp6XtL0dvw
pkafT3XIeZGkb197wYs1jvO54bkTvbwr/r5Juhzpg+41OAMSG+IVTb867jdw+J/g+1kWhR2yfyzu
UlOhYER8blp442vI2oeNNXkUGzXJHPJ4ts9+e/c/8dES4DgAd7pAYj+zmb2sPSQsqBd8GJRuagJ/
KPXqyvedU9gR6le/R+vgopk2jOxDSTYsLJ6sAF+1wUZkVucmqwj6F1Dw33qHVuWlf6dryTUCOmvn
eAr9olkirxD0X8e7u5m8sLYQgJZr7YyLsdRtl1ChZIpHlkK3UnSgBsfGBPn6GyzL7XVYDNQqejLH
ik9snaXXkhQAfkbR5OR/fMMJxLmTGvDUzIJo9UkqsAGQt9zqPmsUE0PqQWuBuPHjr4Fw8LWOUig1
HcBlmgfwF5nt02HbBvuepBKFbR12nfy/4beUosJ4i/2d8Rc123cr6JohZHjRiE9MZ4MmuN0zoTHn
pkZUrLUJfdfGi68OsO/YLealnczd1vV5cJos9auSmHH+iqQimxIJwdB0nO2WmrDm04n+yh6/Q9U7
ciFme8ebgh1RXnt/1DWrnJNNbbDrjjNhinwjWqQIcEQlijBwW7GD0GUZYsWebdzCie48ccXUW4n5
XMAKPU7PIy7IM90l+qYB1A59aeKT7OEcHqsrRvmVZ6BO93gOra2/wan8iF7YHs5QtLyg1xKoUk0B
/ti699JH289QMjYCsEnQavxbFZGWJusW8YtzCR2PcvHSN6bz+HWhOsq/zuIW6UzGr/AaVers3mmY
sKpz8adCE6EYg+RVXC5JZl28Jq57Z7PIoigDbbCFPz1F8VGGQVBB4KrJ3jUwmL3aUJiiyEsT3cyW
Muwi18aHutJ1ZDDU09/p3O90nHidePIeZXYyWqDuqfQ5SjWdYZtMjH+OPg3hZAjrzVlKRlVHEhak
GN2ukwm8UKgWxeFHSnnO0bRCBhlG9gTBQB9BdsUdkOv1+fIFYTckVRkJUvTEsrdOsqKqzxiIL7u6
XMPUtRZuWpdDOcvXChfptOCOveapH1OCGC2Mkrs7eHPet88mYk7DUURBI27XEC5AOLwa3e/kY+vb
RSEz2K2VYlDyMPQ2viRKL+rPL8Wjg5DqglpXaI92d46u7KmnxSjMaDcMrgtYkBlrZcUA2+mWAUU2
RzgYAqcd3ei+nwaTc6f+3WKwRiWeQtvfXB97FVCCy8kP1QCSVXwFafGnk0+mb8NDNVFxZIaJl5RE
hdCB+Z/40Sr5L36E2JtyCI5mnYEXvvAKSGmrBA7ei6ISyLlmiVl5We0V/OtPH3P1qyYjINN3MsM2
MXLf1I0gPq7gra1dDKyNu/TfUyvEHCJkgIDVWcdmI1ZDlXSBxPAQeBZvFT+wZioLUqaMV/aNJJkV
u4xCPAo7XizHZw2xvyBq66gs8imPtJkYksY9DjdE36pI4kNhtlTHPjFrbYtIqbNuj3EZdzsp5WZX
evEmDZVSgRK9Uv/LQ62xcAXG2eF5vD/sadWxuFpc4FFblG3eGxcaQAJADUhxRCe+QrnPeqqhOAMU
BcWDlXo2tnWgxYBnQVaD09cTV3ZpIIJJhYOx2dTgSm/AMx3lcXQ07knEx83+RrtwoBrm8hJi+Fvf
GqcJcRJBUUJXhxqQKMrx6jwoWoh51JTr14S2O4IeE2Nvb1qJUbSXw6lJ6208l1YgScxroUCzndw4
U6pHPnkYW27JuSB8KlCxD+n9NUq3YTGrz0G+Q5DCrm/fGu8oEMEXgBaiaoRyNb7W3zwaMZ5ET1eX
uUmehl8sUzTmPT3X9ITPz2Dmlq8wVh+GR9XJOOIJIB+b8nE7uPofpRAbndy/BHMzHSNW1D1uySov
Cjr8HuygrOfgL+VjbcvLLDhRwDl0QC0Or7equradVmGWdxa/kDfFknWuTUT1lFUfAphUL/5RxNP3
H4Nu+T8nxubDYoPJN3TKTo1uCTTG/RLMMMUOscykuo/3NwQHJB67C//Zzf1m9vz+fUeocskFqzUR
mJbStTmJeb3NVD3c/2RF+zbG0lG2XHjojOnPXBq8ucX4RgRNvimZ0pGsLClpHjqf4p0FpWmbLIs1
ksD/dXfYvOMKmHQEaVjRfpgrtT7BJeoF/twDwV3ETTPH/GVn75RKmsDj6FT4Ecz7NO3mgXZdG8kA
IQRmCaqhRZF26Q1xIXFcI2f6xZSnGNFJxuDi5DXx2gQkmTRV2VSSa1O8PVZjubaEBFqpE7bFdTIb
r6kLizIVTWWVxWZPqgWt2NbbJNQT3jFecIGLbO+al90E47QSZdvQ1UJMOjGcxplBbtkouYfAXOoQ
GLpOwXnT3QeaOVzz+QDhOQjc6pLmxCMdrCNq8MNv4Ql/tkmCxcjVq1zvmDI3sTmxLO16eO4eZSjP
6mLro92REKxI32aB72j0WXi5Woru59egxlI1rKhDKbG+NAdEL29iYc5sHu2pE++cfdYQh7Qxg9GV
rRzpeFFEVjugwK+wwi2ABdXmuOO8cwBDw4LBf4TWoMarMoTsXUI8bqxthO5tlNS3B6LpipKUN9zO
FL9b+fMtFKZZfUFjGr7fgABa6w0mycDeWh0bfft7lsiJwz7I7LpvMgVMaXw9tfsiqgYNRxGGYxCT
7rhK8QccoiCB3p6H5PPYVH6rJXVyBjXU0ELThXI5/rr18cpXkKLxYu4nTv03MfgxBfegV406OG3k
KMS93uFyaKeuQx/DzxVomvcxeLyUXtbN5qmwwi9jhM2rgOpFQVZhaEycgf/Bh+WJ7qair+wqfx7l
SREe4ybLj/N1qMi/HEdpzRcOYXz1DzjSkWxZ284s8GnJY1ywMi66WLieBysRhNuZr6qR03Tep61v
TPWw5WD46xhriAzGd7p7aO+9Kir2E2V3sBgyYD592Uge8UCgDBSZN4hO2z0t5px5+4nbojyN7PeJ
/FHDTczTbAR264FvqJ1SiuT3sd2cQtL7PT9PuVuIDy2p1b5MUnvlZr5WblKGB33jirPjZ1FrOAGU
g3QzuMo2dkSpsYiQzTwDWD4btOKOoRq52p3rzcKkCjs8/jXMjHTdDlz3bT2l1CtcucjPswysF4gm
7ozvK0vyatpSpRL+Stfmj/z9EAdN0Zu8pr0+0BWm9vyuvvy134ZMPmEFJYOjhu9+a3aV0qnvxVjm
WvIEjsAB0v249TWay6RPE5Oi/785i2gq7pXaIhN/eaFh/3awzp9mEUPLH+HYil/jh+R6Ni2AshBp
YzYFb2mS/9NSLMmL46ZfhXNotGVeJF/h5Cwhc21Tzm07xjmNT7TcJ5ldV+RtyURm2bh92/2jmTPs
F97IM1Dc5ll/mZNKq1JtV9f02j9UksG9MxlIdnCLSh8OGf3A1/zgbYXxVQagONs9jWiolDOali+v
22ZjpQ1lWsXDelDhKJf6JOaUFiupjwzmlZ1Uag4MBKyThpi83mEG5q1sY7aROswSYHfxugXCkXEn
ODCy7IASW2JNqBq7nywpX7VZ5mvqq3zWf5CFgfbfibsUFeNO1N1NKVrRjzjqgE9UjZEivwOBtiok
2uUDs4O8uCE3wOwz6tX9tGhRX/pL/JGM1Wy8rl1ha+tMka1owUT/XTuHQcOFmSD0hndpOSTV2baS
Hxg1Joq6xE6TKN7qRxC4wAz3pXz+VO3IhvdnJBf/1tXdZdlEagIexn1TZKdJTd3pKBehuFXwiYeI
/CSS9Li6XPU0qpigmbuRGjCUhnTmbleh6ejVdLXjdpRgLOve9kFsMowPXk9QbfbV6eW+ejR0sno+
hedzJTQ5hHvpsQNVsJwmP+FY8kKMfLfU3CkRk3KuQ027vYrM5eosuQi0jMCvC/Tr+ePlJTmqHlJJ
s39FyNtOAG406K7SwtKu4laGP1ivIO9JWnWzU48E7/z4xqlNKPQ+145iD36iIkpoPM+XVQJ0mNeF
hFezcqNJjgpDMEbRMQft88kAJeogVGy1Ye1Z7NYBbpsrpOGJ3KoqWKd0u/04rVLSnm1FuWve1DZ/
VzyvDTwxgysaBBiyZ/SQ2TiRImzlreyOR+DN0QQoCl3yOT2a5a9IQy+bNrIUSoYYcjrIB4aO4CxV
ji441UtBbbWIthodxItPkv9XtyAFyZN7IaFvYwODNIPlXqGcJw19Qetu9GU2lHbAUqZ7dHSqmum2
K2YgY39qKuVojH0st9sAOfz6LBYqNIwu+G9xQ+zTN4vTBhy2+vozxvUonLbUhrl1MH0VxtungYzh
eO851QJJ+XDIvAwJU4CIZIOwC1USKsqUx2mpv9JjrvcnNxME21IUNBJwEqBBCJ1tk3dJ+0T00BB4
QH+ceddP6L4S40MaDlzJgG0AgJwnvqbEBnN0GtFwep+csefRKzEChmw34FP0LAdy0yZQrVS+J7Px
yo85jVwgguULf2yVikMKHKCT2BhHTfB7vD4HgFeVJgg++d6kBdnJYdIHv9FYuAuknwN72fEnqqTj
6Po95nbFlhrTvqs30DX4wfAATyA4E2I0TqEmdi0Zrg5VmrO7fNT76rwLDRV992Q4KqZJwxhsOBoJ
eMa4ZJEvdxpMSIyejirnu5xaSDfLhX3jFzu2Mg4MGjGiXOZ/Vev4SMFDTGCU28SwSTFalT8tmum2
ZveWU5E7BZCu1op725N1S/gWPZZbbboofwEEQfxztmQyP+fPH0rpS40OtD0JIaIC/9odXUt5/ekN
pk0i3pTndCDOtq5lv5DWRUjG6vcc5yE5TImJiAzlbBzQ6GKe7UUQvHp9Qk6JMabOTZYjlacIYiVy
2jV7/nlT9nNQYUoPTTm3aqOzkfj5wbcJy41lLFxTMYMK4B2TbW/7YDazMTn0c6I3SyDYNc3RGYLp
ngBV+zL0A4bNB7v80sU2CHc8GoHDz1ZqP4RGFeBdsUFifjnAGwBPiN6Rp4GT60KwaWkizcZBa23o
9KaBSZP4JrOPq7YvE2NPPk2GJjtlHpwZzQYLHqJHa9iBkcYZ09JvG2vmAnvenZEvxQnpKIUyiSPf
G4372e+iYW/DAH8746PE6ILuFYeGwwuy7GXVQr6MeQQOU+OWTTFFWoUzJsYWhafxNJTVHkjXgzYd
zvPoMgU69Uitd+79hW2ADohGy6/2cXGGQ+andLUzugbg04xBK7S2yr9khhi7pTQEQdMcH7/KnfLm
JLNyYPQrd8rtiHj2SHOa3O/7mdpGOuo2wuSfhiUvnDWWTXtHEvHTQueDWxZYexsk8aOoeGd1ZGUl
TgdzGDa9WsaT3Uzu99CZ440xRdR/XNVff1EJyyfnhd8g5frWgWQj7NlXeOK21Uif7KYXuc61wjUG
8MipmnxiHWbvbtTgcmMe0sSx7CWvwpFIUwbTvKzRaa5rCoXZZLeXg6TE+7Ol6/XBALWmi8U74cLB
AKEbJBakT8OdQV0LN54cehYmZscmE07aBrS5Hf+eimeTBl3tivP0kyYUpl83RA56ogo74bL3FDdd
DqAY2ZQoMQbEltO9QJBcYYYHzJk5RSzX5KGHrleND754RZazeuRfiPmhCZFNyR7DvSRnXKvsg1hK
Bp4gTSUEWw21Mp0VbT5UJ8ghEi1dMm+i/SrHNYeM3yu6sWcPuyfBgC92sbmY56aH0ZH1/iaD70af
fEj7xW0idpKNlYhHpHjOjBH+QytvWZLW0i85KWm5Mv+Ljn02GwVI/ffW44Tvo20u/yoVcajeDsDs
0BUJwQeTPPslo1eTdFwPSl1P0n2ZOvYlbL+zaaHQ0KIf0rnLHEufNzUkbetNZfjYM7BfZdiGqLVu
fWb07M+Iigp4f4tWm5uw+nYut+YUQlQsju7Lzn80rctUcEWGkWW/MGZm2Ad9EJ4XnNsmJmAihKYB
Ym69IBqYHz+/T8hVfbsF1hPu5xJ7k5LVUCbW0uRN8lzE9QVf9ixC8I/iZoh6ZED3LCcorXJIonFB
PBuNTQhdx6DzbivIDygT14vEu+RVwckoMvZ0W3+rWeMv7QSM5HICaiaTwXnRG0kjKSP0KKFGrAwg
UxfeOo5lwhNBo049f+cJIIJha1O+RrJKM3Qoii2SVOZ9KHDeINBVqDL3aLxZDZc5xw+VmhWjVEO8
jMpiignwnhDhjmdzDKxzLUiohanboJV/dAAa1ooXtOBC0EfJHFdR/JYP9DIX0x02d+TkhfabT31E
0if0ynbIRrCM9GhB2V/jZdkZW+3pZWOXPdgYMFochcGu4YgujoqT/YwRhAWNWU8R9uiLpDV6yenA
kcDfajOdYUmzKzd2v14EdppY5ka7cWZEUksjtksgwC6Eb76UUwoY8elBeFTsPiSF1GZ8UisfS0JQ
ZmUAU9CvD8wuIJuAUC9Vrtq4AzTQAvFB4g5BOMSi4D+3NF6XsnWUM9CO86KwZKj69jIseicVEEyV
d9W5vDhDvmEAdfLh+RVqKnpfubn1eHmRa4VzsIVVRmZ6sAKCgz01gSMtDY7v53GljhRNn4t7Gvqg
E3pDyCHbDibILhI2x/JSl8BSFp5ieeakltkNGtDnKsdD4YMy2yUJdgIQLgWNF7QNT8FUUCSHMwnf
Ygnp9uK8/Shv7ZWnAbY+/Tq5v3g1zvnBF+NrNxi4PMmB5Q2+Lhc+HBV7xtuOSgOJK3CDciNEEA8m
fUlz7PONx88v/HAqiH4VYLwsxmuNK/on/waAKE1Mm624HFs4iQFf1pt3DA4NnwO7LR1RMboUKmya
VcU+s/CHeLbai7rD/QsMuwLpnRzYGiFJc67lSSY7aer8j8KKA75r9zdTvpwQi2QphPrFlH7agXMz
N2zhas5HMf23/qC5Aeu3NCzN/ZOEruq/2UY9F6r5ZXFe2rto18IXtlRT0ujb5T4PmJCRCBKM2bBU
wcnjULTvf76tu2/TAmQpcGIKOcofGrlGicz0KY9n17IljNIZvL2Mrj9dh3jJuX5VXXzCQOXBM58Y
xfHxbNFkJVucvCUloxS+CSTalhJxkshWioK1+DbN/DIXRgRBx35S2oZsliijMA8AaiE4M8Aq1z6U
Y8cetr3sn+QqTMno4oAJXENVWAlsHOWkKhNGmMZrRE1GztiulzGUhqJnnwUhNR6CuNwft0DDk5gV
OO0QKtdvH4F6+Uda5KJX65zPtWKDSFNO1H46kgz+C7nKC1mk45kDBPLtrf09PEw6NFsHFxsmlQsh
i29mRV25BnkOrsKJslbpJfom74xHUqmS6RKnbKM3/g4/oZqYwzC79aSD1Ny3YbAO2PYpeOBWnecH
XcOuvGoEabceREx3pVEhNE+M25F1FdKjCW4yL8HokKUxE6KOVxDU89mrEOoX3Uy/45KT/9ygUXRK
bEyA8obAdOiku3ZVlxQJ9zNUHghdGeWvfnRjdmdCP8Z2uozgbXjAWdBypHWgpoSvvnYFE+XLlW64
KWbXwN34n9t0Yt0qxbSbGW6LX9jtuQfBF0LKd2w4D9lOKds41HQ4kvm0hTEi9SO+z6dlYaJkdaIx
1p6u69PgwysCuLYaHeGsaHzIw4uxP0YuTBWGrdqU3GOdhnLQpnZJjkJ9huGrZv9ZI4ZplNqgmH1P
xPmQTtYCgFg0qUOgNf1SSypSQRgQBAAQRcvqzUhyAD5Uxpfg1wMojJdZFhkHtOiwQx6Vv5NOyd50
O2r86DRSsDRjqP+wt0rfAKTk/c0L1+XZ5SZXwn0kODKPm9oPZnB8ML/mIMGF3xSD03aZgFxkobsx
lKNYx7Krua4onMtmYI0DRJXcS0XzGX2A+uXOvTf21ULBXu9mI9IzcMqAnKcyWBcxOexvyXqh34X9
50B6Q1kKUV6tkf9K+Cb6qrMAD6XNCYo6ZvrqxtSRGmgEbUC1SZddS/5gNtt6/lgniJ0P32cwidh4
CDyfLhJbpV5VkvCgi8UXC87xf9vcVLV7RZnMO1Pbfq5hgtl5QipCD6Czs7ECfQSP0diJBSyGK+Sk
RPul1WTZquamVcCT/VMjCGYLFTtfSV/off3urA+zdPPfETVTLgU2iEFAqUrMrY6PMtyGvsYDrsmV
H31h3fCro4d57DC35H4x1Zaxc+KEkXLr2b4wfTp90gxGwOalpc4dnJuIt2D3LiUin5oDSJNO/BIK
l/L+6IoN8loFdF40ygA1qRd2sXIE407VJPTXyHdKb1uk4qUxBhTRg+LscaLPSrBlOWnq3L4+sV31
ea+Cx2X+bt4vmkwiptGfnjbB4Bz5DKTdXix62xPzz6+rzz9zB7CJwvEn3CPqExA9jkXKXI2YpUUT
cz24VGZ/rOkjIafPs3nLBaRxWLjgHu04R9Cw4ZMEtbBpGQs8YRnVOrk+tRP0eJ4qSx/mcwZ8MaK/
YZ9MCBm+FiVKGzYpIJyOWz7inXZi7eEo/k8jeoMvzJQ52Xk9Oc35Z6iR639l3EoPcGGGc8KQ1IpP
2t1ZnwlYOb814FR4JBszbKFb+NGftsrfyoKB9aYWTW0ojjet0uVaspd0M5Nm9nGzMhvNdmSc7Rq1
3iAUaGVDhUwpkWwz6FnKUu6LRWs/mjdCYHcpzyZJilZSbRAbHtkf88Xm/Sjomuvoeu0HxkIlBiAG
Z/t4ycJq0z93V7nkOfNSmG57ed7AXZjWSgMgPCy9DFRNk9JYZ5UbuZWU5fJeCVBTLbXsXcjx75la
NWvTbOQfBFx5JT9IsCfmVZRcOcE0EhQI1sWkCyE6dfnIxzoZRAmQbbLC1GxunOqN8xYGbARZzy49
FaPFlIQsfCkjeLfMo20+OeHBJNxEq5pfyLEIEzBhPVjgJGiVtc4oPt6bEQywXn/AtSck4a7dpnnQ
7lyL2KjHBwlmIiSn9SVUN1TtWuqGhddrNMWItV6b/swCtclG3puOtAxFGpHNk1xYYH4wtarr4QYt
hNsjuEVXdJRe2FVHjuZpbI2bA91vYs6qIeQN2mt/3t93BAWlhv9ZcDE7m1HJVLsPG8O+AZYTYzd4
CYD8n51lHGUDVUnFZNR3rAqgjJH7xN9/q/vlS78pdVqEFyBFyJsDL1xi0svZs2HiGsgIdDRSqmqe
mriT2vxha6l5ZLHln75vxJBMkuPw4yMgFNDoJqJo+4i2YOLB664nKCuMeSo2DxExrRKGEQ20oQcc
q9q7qFde1s4EaCJJdmaIY3EVdA6WJ0A8BFtdncCRXlC40y7uCXhGrffGpbT/lwAgRz3+LcysKGyU
Erusy+Z53O1EmMn70IaxVQn9sBwqtif+JYjQUA1FNl6j7lDCylqTOiizmbfMQqPvfdsM4pR/ttNl
Dhp1sieVOdk/Fm737qa5I5pOG582XjyAJeXhOagmpnfhkw62zIf1cjupgamYnn40YvC0K3AlYbRD
IzwzDm4KdkQr3g+VNUKgfu7auzZIJD6o2RD19iSEz+mHZmvym4ZFX93sCeQ4Hl8S1FetfqtktDRd
q7q31RBA4mQwjPufWGgO2uwHRRv0WBvcnvTPqgv+JnUD8ze5OrpVU1a+dCollco1gmATM9wLmiJ5
LcJ7+3P8XsSa5llaT91pq2s7UhxWvtkG58KjsS78u34pUbIi0mis5CzSMplHCxB46iiiCEGLJcYZ
xLQRwg/VxGQk26pkmEtdenyq0Pc691J7xfPcUNSlCwCPp67qKELNTUQ8lD/UllocdU8gNwXfj0qb
iFV2PqlRgIaLbB5UwIPpLA5ocTNntnaJUt/U4PreTVn7q0gW8S631zvCelcqWelbhGF0ou9sMmtE
cCLqMQsn5jt9Sz66I9rNcjIsxifB2ue5e6Deub+1+pdeRe3ycIdPJtZsCpDoA7fVZbLM7VNetFly
h1n3bgUUhX/kg8ETYC53ZdzjsxBbBXnuXze+vao4VBMqI8Yg67TNuENk5n2d4KGZxws/XJtu1eK7
WXFn7HHz69NAXN2sh92OmafcWCq21dkfUgnsZ2C+ub9pAskubr7ON6m2CHJ18fuD8fSeUus6d57T
yrWwz5f5DJmDrONXJniNdqQ/0KkRaeq3iLkmnUTUK3AhfWSBrpAM4DXXqzYY32INtPLwpYAksyD2
oJM1gReJwrYbF9Zc71zz1m3XhiAJ/WzUYaFvzw3NQawSgWb0QK4KLMMMtNGmRU5yaTWTFiYzsFuh
ejqjWhr1VJ7RR0Cvcmyh6agOySRbf9c/5i9w3xLKLvgTMbZLqT6JCA2+W6KOH8faq8X5heEStTwl
rgKhYTOkE9HyRSJHo0mz5/huolLN1BDyD03vDR+cqxOv1k6o3EiZ33HGyVgQVsalOEU9nwBggRxv
KLttNTQ6k67SsSo7vKisTwG0MSbcTuSy5Y2AEmhUNJ5X4vkDcXOxmd4UCHauN8xMhTBc6bjkO63B
1wlE7bQ75W6DcFhGFHOCCvGVAwfepnpbDb+CHsl/HjnHyngVVisU64MXxmnvHQvJQOUaYyMaeHBm
GZDlcR332die5QVbHyhWwK+nUEt+Zd3wGEA54jUwRAaKpYI2GSYcHRD2lXMgKlrNe4HIrzT5tyQF
d/dyKOtqLaPHk0Jp0kfNGP5TyZbq8elp7F+EhBz+X3De2uM+cuYlck+I4s82Q2YzShz2hKCmpVXb
Gyi5Kn3WKIQ/gU2j5oyMpHQgmSkdzt6gYgv2WkILFurh6cDYmcM6idA0GrNx37sEGsaHmwUXWcIO
/FzUe7euYaIKYQ25y0jYfv2LUmGJTfzjaRCaAyk1A8PqOtpB7N0gOPQyW06yUrd/HaEgCvNdKQBJ
QTYEtaMfvzTcZOoY4O9SMkErt/BBSLEMo4hg3vv8jq7jRd0+EijJwkFazcWrmCvfLopu3fsi7Lqe
B+GQOBbWuGsV7AMVmjANj0ct8kiODVZ4G9TWOSB1MzYzKfMWx2yoOJuOuU5agLTlb7+VQKLiSp1v
g53sRpTtwuqQaw/CWeknwvZ3NOZFYpt/Ct/BpVNqGdyKoRxLwn1gXJ3vXXr7C8W6rn83F4SQUrGv
fwfUyfb2Njo1RYKuEE1x8ZYuhIfI5c5exEosQGihqncstWLM2YI3P2po+wFNDERaabdEBTcCCbjg
sskMduAYYnDxH6zsKADIoQuyDMP4mLsf/lej+zWFIGWGozNpZFuqUgj1SSTsY9BxUFtwjpkfYEd2
jlXc2fhuOyuCOFHkdnL4TCx6DwdgM5nu0LgtYRbc+jkDSh2HAoQvUGvvu9uYt8rfOGpdpf26OK/Q
OS6XM0DcluIrvcrcF0GaQ2uRFbKPGrME3sSxXw+RZJxNX1aNGRsRMdHrMP08Jf2wtc/5qDhQ7pve
mzYRQoEQBZHItGDdAV6+8YHoncK97tQrDMEQJklPcxzuCMt/Yiee4zQE5OuviDZUbG2oDHRrTLTZ
/btQMwODQ/weNfFvHdCG3MHr1ZitGFTlun1LhnRqr04mQ0yDdKnaxEMZhRErGEWeKpdGtMxdiTbF
nA3jeGfXQJpxLtXzQHnftrESlItfx2wxLRB2S0375kOZsNGFYmEks7cWXQj/nVtgueR8O7YG6slx
yhC+M7rntXBYFMuPG2gUR73O7Zi/51bh66fnh1l58bbJonpVdVeHOPhmQrC6iEOm7oucm/Emac+l
PwYBNAMwv21gABoKFeRO0l3JNQsZOmXtpaL7ILV/MYgY9PrIFKahbu97UIrycQutKcjFD/CEnAM+
uRq5zoKh9pBxTKKviWSgkU4XBspHzSKp5zmTwHjlLpzrupBHsD6bJ1dERTzTyo0aj98Li3ObTOCr
ZmzEe6vA00592tBeK4CVMomwgaPYCiOgvuevNSbpWLdJqGFqEOxMpA8/QcefHquIm14xV4kwbZy5
jc2VdYgfm6Sn4DO/QlQDYRf0KTeAAYwTMuSzGymL21OTmK2ivWG6DGYVIhYfz7l8Zj+u/tlnA9pb
OAc5Za/ZJEHgquk3BAQnt1OiX4DrD9kuXpRhVbHDD9/5KYF1aebJfrFHVqHr58o80ds4247tMifz
e7BdITmVKezO9SQplEHn5UO32DY+nHyKQCGvbfDRNu6aVqKkhcVd2AHY73g2aWyYMJCyK9dd7RQS
CSk/kPWMs4qmb3j9/hBDRr6mtnekdPKikgWGFWx+lUxlspvTKi6l2avqJIzWRfV7ro12nQ/ZuzUN
IDrFM32jNqQaayz3Pu1c7ILMskxSjI47c9TSGWSRcZf9OJgGD3O7pmcI/Wrt0CtHDwYUNgDrM30h
LNmRCQicYkoFHxVj7c74o9blBsMR0IrU7CcigbJo/BUnk32En3bwtMgB1HjHbpdRRDm88h5HaoSO
rrQAkXPWX4R7+JJVm68vnBGNsC36FJCSyIq+Qd5RnZ/+iOJNbCfjZxoMOusxrpnW9Ht7o/QESDSE
lfNVMaRL//C+loBtD7ZwecbnjFyvHI9v1+iFEQ68kNkiabI6ErLyDhNuNaa3Xd7sZbQ5m7AvF+X0
UMSSLX7TfZjDpsCAivNhZ/RwV8v+z2tJGaSWZ6PcaWxuwihMGen7qmDCNf8+2tbhtLzZgu42JH6h
cwxbNsMUms25Bw3ZMkU1ZNf0fdgDMFHenD8rRrL56gg1XzQ/1ArApBwcVprSEbbRCdKwdgkwXqPg
rpsahtG57lKWtTUo+8Wlf0T+HjxomRpDzRbOfvXIdnGCTqLnRERW8vj6GcdLbBWEf/qIPFpWD4u0
klNL3t2IDzSFvuqo+v0bYsDVf/VXMDFfudJhqralUPJi/6eMMsuXrrIdZcFMgFC5y3A6IRYMxebW
toeEkA74kVIRsz65XqGUIm1RgcxjHBSuNhMzJVd3ZXTJApYuUutIJJh+kCoh5MMRbtm3LEOVAdVn
6nfd5v7qNMxURThzcvSyV7PSxX6mT5WlGwNgr8jyexinsNnsAyoGD9XcR670z4ENIU/9oVZTFkTZ
Y87swa4kNMFwj4b6VxVQ/sM7hQS8seOYDaHb3A5E+i4kHZ0rF6KFVSNyR1sz+F+CYvY2VuhAt71x
sCvh98FNN0kfRJ0g9jMQx3PdA2ATkI4st1rOZdjrt0/9CLOEfHeD3GVbPQ7jKGbjL/K87G+rVUT9
iIpuZV0MkCmzDdJ7hw+lKkSRQw4wo9j6NIORBZqx4Bzkg63yl3n91xMAq8HiCrMjC8FkgNZlbJpg
n9mkuvs5tR4P6vHB77I+UVB/kpTKJFsG4GvJYi/pGqrTnY4QVjQ5DRW0LJqKBcqBlBDCco3iTsAs
Hj5KuzrbQ/i+MwyRjkRrdLGR4WVyXKcmYn2LD3oq3943osuedfamkyo9fU1SFb8wJfBoc7Qf1Atq
g18uh9kCR+qyicZuAQcxmcznpIoqVwYjI/EfMezoNARXtRekE/d1QAT21GHT9dOsi7+zosNccLOd
C7qHcVd+awhoeSn8xmsqWqJZlKtogsDkCDfvOpu3BF7htNmdvpQ0K5ywp3K7UYpB+QGM4hXn92qe
5TUj8cs2DRjUozTGWNSKiFsKis+vTbKFyfkq9LUEVnFYfcSzmgRkOIZIiY6MPSThS8LZwLUwQFMw
N24PIr7kZMPE5jyd1D2+2pT6IEUAkzRFkncmkcakRIE7W2VYR+rU+jxPidxt54FMLLAjO8GKln5f
UowVwCuoyVTEBuwGDhQqtVljAR8kZnmTWQ57e5EZQSCzrZk6v5QS1PMvAaFUREWtGgpM8kVSAxP/
k8DmMoyEcoc3GLC0puOAbaUMJ1kJtQq1WncLGWTJ8g4TkFjr9iMBk5f9dbARF6AnLNAqnZDTZjkh
rPIDvKA8/JF/sWzQ1uYaljY0Yh5yctv6dkW6fOypDNok0pq+cKbJkFq6NIHj8NiQV5iPkWVRAciZ
hyJCEUUUk55xQQQw9JicefG5gfExDPaUcskSrgf9J3lLSIOFBX6AmIgPA0cFApAv1E6VHUPhk3FN
nSmJjxHa0aafnGcprdC7LA6O5AtQa+PQF4IoJXrkTiGAKqF3xfjIuWLiLjCE3A6TPPEBifGjuq2U
puk221nkugcLSeRKWHbtUCgEQzcZciGD3PkyGqJ/vBrFNC3mC6fp4aTxckdpFEAc2KZx1LimRs1p
RQs2Wwq5jPTpZ7m7WuaXytnToMgR4muUI/PNekkBGhfa7mCt6PwWf8go9WdEvs9a+UjLoBl8GwKg
eb8dUyxWOLPYy4VCaW2J0aTHMcKu0rPs+iBt8hsCmR7oV0K4y8wOGq6yoRIw2BfEKJ94EUBvwc2S
sXQAHwCPzH2OxRFtHoP7C8+rAgXhI6xRJh0pC0raJFszBu2GoOuqfChzYW01xKMJ2ZmaoC8SzrZS
ccalRFXtEc9xYIob5T4WQazmXfmPV3T2DAwptMw2hI3tkBglb1G6+uDRVubJG7egbfyIIkYMVaDv
TRPDqDUAD2R8OiAPZmel2kFOJJr2E+5DTSYGcOL09lRlDObZS364rs5FrrVgYvAAx2osMW/qPsSX
NKxgMwdC3oubAFGaMw/tG2K+IwI1pPs6OVaMSshZ50+R/tMWUU8AGrC+kE+ue1ONRomUgcE681WG
1+9kAah/9kv6V7YQgjeg2ZYUDhdTVlzM2vUl+Yi8BrEpbUyg0142Zkawpkfz0fsVccEBD+9qOQ1V
i782PucUFofUAqZiPbnF5cMa3fPQmnFw1FvVymAvI9qxkiFB3jLRCAHmR8N7057/bOYbXAEXf366
eoPcqRJGUC+DEgKTpp2BIgvSKmThedRkzdi5kGiZGwB4wxFnMUnhnWdAoqa0gSwPpktt+BvrSX2/
W5JfHqjFD8an5UuT0MlV/Cogu8AtYYu8v7fFLlLMX/Vy1Fxc8LKwDtmR91ANj/lcRzQTV97GMBXG
PGa2J/FEKCWY1epHAwUqF3u05n6uZn18KUTfnNWRB9Q1UkCEYy0QYfGLfBZq50VoQFuEOvC32PQX
PFO54Qt91ArOLGxFUXTd80mK4bbZU5OA2NfpYve077QwFClXkhyQr/DwOu1/OfEqnQdMweIlY1uS
D99NwEUxbHti77fpduw4/u185D0voQ9mbbEMedlMztUQKpUgdcgALWQnXbRQuuBkonuhAGv24pz6
O4G090ee4sSGwqc8iQVfDYpMvUlVS4OdUydmJQwJwxwPek/QEV+CWLkFOfiddwYJ/P+XXZaa2OxC
KT0ezeCgrH1uG4W8MsdaeakFwvB3nHlAeeNmWdZAyfk4r2IEgJ3rl302dHQuWAi4dzHYQwDfLf0q
H7JqyhGNBBf4bbQyB+9iUtnPjqNqF1LibGwI7BLqjowcm0lLI7KD7bgYII+IIpT1iIxCX0Bn51JS
ejrXzLZWtABNl5ts5ohxgoreMn0Ml/ZDd9AsecnEWZJP765huWM4ATODP0E0vw4cBfCq95jd/pQV
eoy/n5erUQwbjSKt/jYj5E9gy9Q6ZrDbtS4RNqJ4kVR/QkWjUVj+BqvPU9kNPum5Xzj9waZg9LlB
hZ+htuaG+3XuvwNnPDtgIllm1618CLwyMYyP3aCE1LLQ5eEXn0gG79Ul71gCK0KEup8FTzEGbvLP
+bj61Jh5T/pVtQwIpOEs/zKUekVi5hpjjGBjiAdRQiW0eh8GXME1GK6N4MJgGxRaqIWcQyRI8dlc
k4Ct13VexpfSrkvzUNoibvNa9B4y2T3AdbLtyW/z1sR4wKPZ3jJ2t7YJ+F/oPdjqw260+T/uqRsu
z5m+akaPmc2X9sXZEeoVZkRAObXmTjW0XCPLj/NRE4vZ9EXWY8iWA9wTYTdMYLdwzkiia+kcnenw
61+MPNEMyShlE74a14bR9xOo1UpyT9ZI0mBmFjSBaQsyz9z+G6AKm63B4ybaqPbeb0L4Ra18cKsQ
1t9b/HslYmOqd29+sukUH577WQmoiERh+qoZ48kADUUzDShystNoTqEhMJy12xhtnyVXLiCpEyeq
28I80+u5YN8lwHZDnIbDClyRCmUjHh1ZA46yzqIpFCS+DQn+lfH28DekW0SVo8Rd5wSHSCgq6APF
tmvc1YOV9h1UNxZ6htcb4Su9IWomVp4NgeW2pNFcL8vEkeX9WCarlq6t0GzgHjg6LyWYIOQxPZy5
AOEKkOTFRwyrq7kMWtNVKbDz1O3xiPKLSqmOPwRgMq64oc8BzzYT9/IdcU3rMJpeTeERnUxFMZpX
DKXU23xmHw0zQlHjC6cKjxR/Gv6Ybcv2umd5HNyBtz8t6s9KymK6AI+J+bDydbd+97olW61aX67M
EeGUFSg8IpH0uo2ZLDwAL9yLY6nA5abbLvVZgsXjyOYFbe2dvgeUWFrwS+lJ+apRJx4th/mibhzl
1c9Q0S6I0XPodE4Okvumm3pVpY/lob5HMAXQZNUt6Zko1iNHrb4bZx0dA2cjwoAt55QenhkMCQ+V
/E/8OZEX4OFX+kDXUm4BtQrpDmc8t+h8itkJRtrfD3y7a4NSRNzXDsZV3hvegIHozTtbUnxpRSGt
BlYTHcmy6zuzAx+7tAlhvoeoiZYUEoNE1X5Cnf90uGydvHa4ewVfDkjWbl8FBVpnzRCPil5i8MH7
wXDkWe4FnA86Xv3G2HRtS4RvISjN5vFwXed+P0hAh9/EHB2DDRkwAhsL6ltRDCQ7M7nH+/rKiw7O
lksuu6ek8zDh9oe1ML/QUXhQpjQbH1drbDD9F2FkvcrIYRmwp6Oqm5xYbSAtWS6Ea/i9DLZcsH1m
jwSDb9CddKXrNwe2ogcJgFXPalxdMGW+hToP6QnJiHFtm5CpKq/4+TijgJyVFp+FlStl9dXAkqGX
9AxmteN/oKFetUlyooNn2JaNb9QIhTmhhabWqlfSd+EFjV9/ztrAJjMgAWAsQgWqSzjMQ5rdB3Fp
HhitVUtOwjCoVTvGC3nvX5rKEApPOfwkHXB3yC43GSKCLJ+4p9quea5HTdfNfQbIU0p4p2pWWKSj
WqsHSy9kJQJWT9IUQN2RQtU2qyg0tpoTFgaKiQvCeQBem2rtLjSjzxTdSboF+YGMm19O0xAmUPgc
r4Qz0FAdpPB4/0YSECN48Yh+IEXwNlGeKqd+xYaySrKrX3KgyGw0twwIrhkf/p+UZVc62a5AqFPT
Q6EoLRgt737FM0x95snikjkrLnAjHKaxS+pBWc6wtLs3xPqzTMEn6qeKn4Z1GnqBodKxer6oZEtp
3e3UBBUUDbFMVPqFs4cIi1GLV0HMhpcGF9PilIBlV+yDrsPC8iWS2uUcmYTTEKv/z6akzTWGDH5Z
ZG5rV3xvpY1Y1tyV4IPt/Lr8zCiDFbO6tsl38yQMKGf0imVNWQxFvCNZQDPrGauAdfJJE6JDMgzY
zRmBUMU+630qpwGnuJEGtPKclcbSyHamEXAtEVSjTgsAQSt97HMWOa9aBi0/6JvXbGtf5Suouj2A
CoeG7IneGN1vlMWLJt7CaEM1PQXXQhqXQyvntBIqEyd3cdwi3QP1Q3dPqUuBFXJXOKFEkaqeCvsu
ukczl4El4qLeRCDqlLOdxxJZ0keimRcMM5FJ+pUcyGk1F/O7LvdxoJVwZdVR6AcMUJLWWXxjX7lM
E5r25DH5rldIP/kaSZIEkjtrB+XD0B2O6d7lKfSefuewPFA8WJ/QdyM9PFLLrAaD1CS4huYRzZRS
NGI+q4bvIGtRsmDZszJ/yOlpnbmjOaqJ86B4jjECtGZR8+76KHhuAiFr152qW9BBFgPq73+rhHUv
XtFz20TZuiylOXGZlkxjT/wx2/4UmTcibVaJ5hrR0NyIV06TUtl2RhNvkF7YEWJBECP4UAgbbNKt
GiS7hm7meLrT8yaF+d9ySX27su3EQzvSzfFR7Q6zEBNsrfgPxq/D47LqHoKfvVViYYBpje5JfQhz
+uFry75/Cig+5xZcX2zuki+H2gwEtBYipeJkr5foXzQlScQi4dwBt4kr6+d27LcAPN/cmS3v/cPN
JEhEvrCRu8TkQfnai871mLGaOM9sTgDxG1G+VF/WvTmriOhQh5WFN4YeE7yCrZ2yYq7aNerdRKwF
JPImYYWn+8K7se/i+7f/aAiUKoH3Se0ir+bbBathJsP5OgQl2u6mk3XHdkAedW81mfAbh61I/2ls
At9cWTrgCWWaxLOxlFo9N1i8F6kFao7SovsSaFRN7aSmagowk2zMp7sxHcoi9sjeR10MHpFryL+4
OPjX2QgTh3J9xQ3eeLfLxexffd9lngSctg8jfZ+fuialQA8qq9NSZQkmBMcVLux691rJO4s1M5eU
MsKMsppSTc2MbjVlqZWi/t1PBWY/RXsHTvINYh7T/P5am9XQCU1Y8H+sdK8jobDhHRvWTMlNIcta
CJcLyuyOO29yaXU7VsYZyIYr5p9R8IFTGKOWx/Uk1rVo6K2rKiC/aB2qV6TLqyHKuvM3sxn4MTR0
joURwLCmP6I/R1LZ13UsdqFnnmWrz8LJUw8lUs9Yto7xDkwtXM8JPdV7Tf2uMkSo9ACS2j/Kk5bC
ddAsgDigLpS893hMYzxTVMb3rVkNd4UAQwd+k+tlDJ+GdKeDhBB6ihqkT5iJbxr/+oJyHr5Nsdye
PdG9jq9Yp8GLaq5WpPecKc5vds0HQpLnvIck+NFgB2gW6c8YL8SDWo3cN/YT//ZLfHlMpcvVOqdo
5dX5d2WfDlsHU9pKkD8FrRlK+MJVL78vbexGdpgFEqsVXL/lElxVYaRICN/5Sqb+Qc1/p36V6mT+
h4j+ahaGWwniCDR0lNpIU2G06NjYVBBpYxDFxaJZHL26A/LNAqcoP4U/63LJfXMHMR6Q62WoUmfe
/zr/8lqCrW/4gHIPa2zOzyFjTXSdoN/QtWTXOIueC1wb4i+MDgcSgsurcwaRcaOQhaNqmC8B8AKc
Wisn1iq+Dmgi6gbLvv6mNDAn8LqiXXW3VGEIm8HGAvCblrzwdQ1TmG3Jf2+9xYlXGiEQk8k53ltH
LK96qPOf4d1akKoIiEL/YEyt3ZlQ4EgvvITj7JS8Vr9/8G0IpBmVfj6UbS4kCd3KaYgBUrk5dskm
6Syzq0QBTmU0oc5HgYWzyt/ePqoMvBKXJCDao4u9GjAaqNJ4KhDAo4+41L4I9pIsXIzLe+YoTh7m
BMXM2hZ48DKrLIPNv8OzoXC01Hz5wJ962EO3pqBNvh6fZsqp+b+ZaKeDG/GWQ4ZHe5qNHwPdy/NB
1e9PNOvInOt3NwgI7yBxzaOFxeg3DFBftLxWyTJw8upKirJwcGZmT33dY5GbnL85YqJO3Luw6VVp
vBJFtM7kZImMCZ9WTCvQvik6NsquDfDOeSrdIQgqUOFxCDwHpLTj+2s385KOBXk379PMGKV7HaHB
wGSILxzQrI1bPeTdohWJXBILlTIbo6Ow4tyadNBU1UHmncjyqes7dYM60nbiivMpGKBg4x+V/HWT
eOOrJfNuWhz+3TT7MEg0cnRBUJ9Jw3GqZcnnEy7f1qWPAv3pxVCKjDR82/3Ibaeur/2T3eT7hVDz
rp59IQ9XA9NdY9pwbYBr4NN+kZGlqmt5JwPdssLoXmP+toMfv0rJ0aJ8o109Ame7uYGuQRY2cbwG
Xzn0gYvprrCal5b4ZZl59TyMNhMlhuZUcyVPWpjEUAGn95BnS9J7Q7yVX8ZKuJja87Lu2QDes/aa
xusRRBrxbDqa6pgCfWTNBvS3GIBQ0p5fhfQ75T2/XnOPZ9zb9DWUm61lAJRA52vRiCxb9uTg+qGA
JMCIZ7UhWS7T5FAB7w9o4ykRjsLE+SAebTr2t78LeSHE4A3kGW7oaNAOowMy74LdHL1FDPQ8sKGH
VwaQ5/bXh2i2v/pV0o0H/CvyfJ6dU016FIfT1E8cY1w0FGfW2DJToyYQ0aTsrDUIq8wM0yLYACQI
Ahz++vAOAavLG/lukfJ/EG/k4qvCLC1O6b5+pqFya2a+kivUg0DOlvi0vH4BjRaCmnAhIv3AMwGZ
Sgcm5gi6tJj8l+QMZdsexpyoCDeVevZmnlkPz+qWiCKbJTamI7QNc9Qvea/5/jT6g49fZJBzqC6J
gLfVJaFItAViYtXx/r3C3IMo4ZFoB1PNpINLj1ZiPTfipTkT3Ub9qmtsjMqWxqMfE91dTPC0xOr9
AtlJ5D96KsdDrXg7ZQp5HnN2RhbW0wqfG2L+mdUdcpFhHPczgJrwcIA1ZDFxfzbmpZ/koXKGiKKN
Ldp0nkUWTqmdN138cagyIJldveq/HdZltxIDbqJuMpRQ+MIO4ypX1uIFbI1JnCIZ7J0ZBKBWUzdD
F/YTjfykDdBT1byj0YCQv68IKTcTzdAFzertQ+M3awZzOx1e9uMy7H86KtHk1ojM8muu4MCnTTgC
roHdxzZ/cEBIzRpFA6IwlgWLS4P2n438g8uX9nood/AKsjSOv4g1NOzLedAPrW2tTpC1wwBZg5AI
T+lyMh4o31ROWEn3c+etk9O/17+VWgJPXM03MyHA18YIOqulGOSEDlPXdAvs8zOWq2Rl3q3tADEJ
qS36zM4fmEmnJJu1w//WTo8lUVh2XC0pjQKPuNhBL7OT0Kzsl13MgZb770ItzHEr80IvBXY/N4f3
iLsE5fQZjUhkm5vxJZglros5zm+1aTBYkyXXcH8/1KzrxL3ELMY1kWiOZOawwmWjnFe02VolwqCi
hqcAp+ST+RFOKRbQuYESnwWMlNeYIuQ3Vz7mlTGfXfIDO03d1aJjE6Ip4qih8pssMbM9SENjv2mN
rAZVxMvuD9JJPxxUSDA/V26v6DDwwFXiNYQ58nRWylr3WEy280T/mpDHw9UG92346PeuPZfFmkzx
FUUdIw0Pz1jLxRtysDnjCH0xJ5Doph8NWLVUlFBb/5Yx9+U8r5nJiuWwu6oJqy5DtAaFnPoB8Ib7
tPd+27BHbP0g3Wn4Qd7BSGlauESmZYnPyADHo61g8buibpfiGFsQ7Z++O8NnQu5rWQRmcjCNjWUF
MJsI7rNW0I8QyAP6u2izGz1B3LO1E0lfpaZmTqg62SIcYpGYJKrbltxtc98VSEcyXWdI3Nk+fUMk
qzgUzmo5xVBq3/GVLr1IV8f60GhGx/oGc+0TCSqTzcImx+uTG8W3dITXAwz3eTdQFRdX/lUjfkmD
xgoxuC8CIdcJHlCPil0ZUcvLHfy1wES3UWt/DkC0nD39h5+jXzH2JsTnY2X8HoUiljuXlfoMtfvX
4/tqIX9EeUuH0EuWPr3T+9dqJK1QaJlfoKXfrkHbWjoBUXhggt3Oh8KC7fEBl6J++8VN06wCJA48
XS6Em/YI0UlaYzRldRq52Pke6Ux7vDKah6c1aCLYQjcnlJourFrRei4KkZx+IlhN1+Dh0cgsEugU
4lIiGoacH5wXXkoAhKzxf/PDWEnj9XSjghJlJ+UByBeQz39MyWgIGtN9OIOZSASxPcISZnAisgt3
wQfRHkYHwDfiVkCiRYKEEjYwaD0JwtSiYUsyhsuDAQTtZX1yQAiUy2TsgyOmPPBsxCA03Dh6k8Ys
oAimsdBvXkKARrmaO5TSWsnEO3LPg677518dzg7aiOEzg1Dfa8zqRda2V3uUFH+iml8ouwqaScHL
HJrB5IT+kQlH/ZItXmUU4YK1QfYJCVfPVvpUckr+k9Mr0gliQx3IrhgEF2fiwTLqgzmsBtiNBMGJ
Mz+VvMMa8MuPc3dSXitBx43Quf5Ih6pYCxfHtR5B9XwNnXdiQ57dspnU62Zm+TDljvOm/XBZfuKM
tPRECCpjExN5aCAVFrjQ7jsObznmqXG8CFQkdff5XDsIIeXiMiRfItPLeqLXtLSk947M5nYmNYQn
eW8dgMj87mrn9la8qn6+4EjIlSqNXt9aUjn8jQcXsp4PjgMbFN8XBiZYwWTIeollEYFiuP3UWgQq
J11TWGBATyGbV601vx34u8dGAyvnuIqefYRnLl3U4fLW3edp682TZe7gDHsgx9c2Wrr9UFT5zgvm
5kySg7BsXHZx73duzsq2PytkwhAwotZkIm4vkBJGZLJz43WEp3tlgJllQtJw2fy0sAQsWfIL7RCg
aXfb5skn4zlhv/Z/2iwYdnouy23yZWXAPA0F+9h5B2pBrzvoyMKQaZSxQNCCubPteTWfZZJQ1blS
RZ/bMN3S7TZG88oVvVSgIFZ378OBadOam/s+5PVY0m+C+l4acpktqcVodaV48BtAmEzlQFi2SEa4
7DXUnP5BjhetwJgP7no6dKKpPtafPdBuqfp0QYbfiaZGzhqg1tnAn3pbBMxTQ3FpWwoVVePad57w
XJA8PUMQ/V5Y/0qof80thw7e3PHl4TOOmjQxM/77WmjzKGaeEEM7DUyouXEDV1H7xYS3H20oOvtv
u+a7SJnKDnjayHtJoPgP9tcZHlCRUinO204GdjHV+vpehVQ4xYf8pSd+V8PxdPHeKg+SVQBqQqg0
mPA1k+AYckhe7DBnZT4TaJWZZko+W9XDfdy874StJLSsEwQrOyaWtgUg0QVU/nxl7Sp0r2d31OuS
J9feg0UictAbEBWUYmnGAz62eOVkhr5hHp1FV7R/Ts2KEQAsyl1yIU6UIBQUwKlPzVt5Vf/PFsnf
/18W3ZsIkSxAjnVmqR971Pz5Dl5vlrfU42gh3YRTaklj4Tfv1V7GxZt4VjM9w72yFrAEGPjB2CbP
dQ281SUxRTLps1KJpLB34cgYxA1T0OceZQREBMojqK7/jNYkDwa/Agm82NJNpQ565+8uLubO/czg
7+zjEcLjHjqyBUpGiy7Er86L/nQWzbSa5DpPXla/qV88wnQpMgoi8R8IREjJmODoxznZPP1ZO10y
iaeytxydkP6lFDnShWi+XqGZsmnJZwf+LG6ZaUXq69gyd8iC/hVwK/YpZcLF1vSYCZ3tTiFKyP1i
rAwuVEQ/nIUrLXNdGgKzoNNeY1qbNvQmQu9MLcLmZ77M3rM9Jv8/uQ2C+4le9R71p7jJBH12nPoi
jTXggUbpp0AOeQUss2Ut/jtr2o891Cly5PDpfEi1uZWwB0ILfmivGShKBQdlpz8bnnD93ft06gXs
g073NEsubvF6qsnlBKKqAVv9RTuiKgfhRYf8uGzm9nMVn3Jz3uV74K23PO/KvKJg8R70CvUxCJL9
UcAYhb7QchBGDKn2+j7kVBMMthkLAXaGXYaosAuqSz18ZzvDgW+Rcofs1qIAfv44zyZmHQN+oOQl
cKxKzyP3nxg9eUnSuPC/ND7mALgFNS/MC92SxXW6UttuP4pfRlvXlao91/0aMApjW57hi+QeGqI5
7rbeST2I2LVGbkAZ8tNwFOJ7u9r0g3ClHUIKdlz/+ovZnIUl3kjxoAI3Zx0mAJvrLm5BLdpJR8QP
7WlsD+aWBttoBNaoPUsIOX6TXUd6wl1nSmUFmgp4a/BjZuse4DAPK9tTthUk2zUxQUIFrcw+WJpb
KqGZJkGkKcsYguErgOEnemhKr27+AtTc8eIBfcF0IrVm8fPQnRJBfntKh+1hgRV1Nj9McnXtVMdZ
wMUvLRcimAGDOEl0E5zGFRFvqiTjVEns4TMKUGKvItT1pdsRZe13GGI5XZUdMWmoO73mKT4MZ6V5
/1ifIplkwkDNX4R1PcqLNQUbeZozvqv5U9y1N1JsM6i4z3gzhR02SFDO9ZRj82HbzhXZZKettetW
nOL648XzmvzrCr/6IXshLvaD7MjTrwyeFAlgK4QcJlN9OkTQW8YZszhmKZL63QZWBBDOYWMlfIeE
L3AXA+lKTRTpkNrUy/1S0VRY6QsduHr1hx5S5M8sfPtN1e+x7nnBZI+udLJRJAGZukVvT3iCKdCr
+s8esW4Ud4+f1WAnNUfCwaiJS75bG3qjVYS9eOCCoIrbLvpEJCuHSnGbwIu9OIfIOLCF7AQwloC7
dCBV95uxLLfsoEPObWzj7ioHOKoTsPcVr+hVcoXKwioggslEdPcmLytan8ajc1GwijyFzCxq0fFT
5H4WDlqv9/2yEaEBefiqECSytoHiZuLaTKXF+dCtz0oBglI9CrvbyT8TjpdA13RlzjTtszN2Yx72
V6jnO8dp9fy9iZMIYD/XaH/mOjyXagGrxyEm1vwqw6TK4tCYXtJJoz46cPRSv18Q0QMQajuupl5K
EBtsODrGg7dp3d5aAvqqGNsCCw0bJztdjkuM7wm5pka8AxsMSDgX1FGQ8sRYBEbFM1F5rbWKpkxJ
YPPnSNyLS2oFqL0hy+lDhyrByWRUIODzzwPE7XYuRY0xmS+AljrwR8w/oOj28OgfMf+CzROiP+5U
FcgqerBWzhiBmxqXxSbPfYxYNS4tlvni/qKpi0U8ibXhlAIhaExmlu/dSJ4EOmb1z6ceKH52p1gJ
nFOriVcY17HKiz93nzpl7F4GBwPsVL7BVDmMt3UrjvWZ2PHs4BIxdfZaaafrP+Wlt4n/rDIrCcv5
cQafJ9NjukDADk+VNSZfmNHRZ1UAzAlUSpRc971SdTiLPkrwxaP87OUF2KrfxrDi0Ik2qnEnpT92
c/M3YWc/2ItagXYVAWY+kBKgxA2b4s78QaGiBENBXZKXV5h578fwVSN50ey19BZgWGsgbb//eg+f
IbY9O9J7cu/a1PyIgRKY6MTsjpp982vV1e8mFEYHMW6YRbv17LAtFNTJT8keJ/Ejf+gF8NsygpnD
h2X0Zmmr1bFFl/7sFhnjbzLOx0ELMq95eYCnXRjDnjP56dUpur6JHoU0G4r75hvqBcjFOFXPThq+
5S+bYbKM2w+P102WXC34ueSZ3C0wBJi4O18S+5of7nVcuK8WYPDDuIuJqZOXd7Ck7jyAWLY5lVec
UAMFJXd9S9Bb6lMND02k06BYU43tltgeaejMH8pQ4iRpmfLdMXw3OlBN2AsrbTuulBKpfQY6iul5
bxG0bkpLGc4+m2OifxGjNI6g073iy9VWlP5cxJupWOEqO9Qx4+u0lZitghSNu1Eub657hoFFnpWu
VsqDooTAiki3Jh1KC/L0+RZYEiPsye6jMYLGLqoITaX7ghcdsvLwVLHuJUvtC/lEEdkkosyr8XGe
4xJDmeSWW9jEajq/vjSwBEVdcS5/i0eFU+zy7SksoN6fQW1keIoSxT1npQygv3dUhwoY+Q1CKw8M
7eIJ85w81sPRXKYtOnoJcPg3XwL1Bip7+HYnR/hbDn3GIg40o2woNrrsmxArXGnrpmTx9C0hMycu
lz5/9eMAJmQJSeQb4WvwzGwKL4dpXPXHLXEhI1h87Gyf18h0a0q0UeiCq3kqO7Mo0zm8jZxfOHhc
uPfXTWh0NxUlMHDtW7Pa57/bJtICqdhX6v9c9W9oVkpaRYb+gNwIduiCKq+14JMO9RJ8Ugsj/PMu
V+HUpcD+wbeco+jkSHA87tgXCi8XcOXu7Ayg7IfPX93WD5A+hb3jcOZKoBu6jCQiusondQrnfxEE
vvc5q6XY/1bL+iUtiiKEl9ho6aQC5SEXCAX8V8mXkYa8ct6xHaZie04VFEkeExd0kvv+jo6VdJRo
l5/aKOVdushaH/6k+WNpdSlQ90VYOjnE6TMHieqCtLMa5g6GY4VX4x6ZAZsBW/J3ImgK8ZYgfnkB
e5Dox67l0PnBUJe2z3emx6UiUxCeD0qw6XihaQA+94Fv0mDGuJlVHqxTWBVdCvdAI6i0YC2rCiEB
LUyhtk7HBszMHnw9IhTu8mX3yLVRaPYavhOq0ErFM4CHxdugy6amQgo2Z7+Dcu7OJ0eWw90mv5Zw
gxiPNYwQmtw0M8NsYWZuW41VzrrMKQlgNp9cqcELC09Iyjgbk4Ko0jcmt0fkxf1SOx2/uNNy8AXj
o31vgYv7AaVnFFUpfuaGk9UTkdXfBTsoBUIsHqbW8W0kTuVBt+G/sehY8wuoDKGcubiMzA2Kdya7
sMWK4p64bcvycbt4KX7XaZSMLufNz0vQF0Nx1oIFI4NTe4H6G/PXW5NMY6TFmntLEpKSXy5R6y/V
skDT6HX13Qn1EhNALXu8rrwLIBFDS74CoxepbMhL5sitdwGk0c1I6IBdNl78KryDP+pJxDFztspf
xWE+HBwFSlq8LKLOuSxF84NrG/MAIR5d8B7wwT5Wj2WE5Ul0fAJfu9mKfjWAMIh1njen45wxcKTZ
+IJebwS1ZtzWZ3Dy+ZNiBazAFfEAo7nTXsTNTKzzM6z/xth85E6lh2MgTUE+EkKV8b5+SW/6DFgY
+jlTNksDOuwA8kAnM4V23OSdVbAYYyjoodJ396ahwRm2rF5rDwS8jcbyX6xULJeX7MPgpmtYdSPv
noPSfd4v4JttZZMkXc/TQbcx4VPoVN1gXoQ2oJ2LGLqD8YsACd+GgMbXwCQom2L/4fs5RyoRAZRv
1gLM8w7mPC9I5L11N8xUn4JvgDrB7qojT+5K4tq7aOi3bLuM65GPHoW9rDAjTfRsRQhNMK4BEdBc
xyhPBJkUQTr6DXw1d1jGYuwxo2tC2uurntrgmncdXpeV/jLEYiyO/oOtLwsunUQBVxwXMIZNgh5Y
o2wBF0/kYA7zf+vi7U8TjbVKDI9eg5FS23Wd/NljVuzpizvtYXmUxLKu9dkj0GqZnpYWhhL4f/sd
6Xwz1ca0GfZpGRKdNZnJLhrWqtSeNwDT2A/U9CxrJqbCmwWV7XjpQzyTxwicSU8SJYtLM2nUfKbV
eMYwUitIK9CUjRHXJ3/puq+lRmIDMmUij8BkPo+gTRLLP/GWPSPH5RoUnDdqwhNRWosBc1r7edBx
xpB9MVC4tvDczBTJ8jlQGYaxqWtl6FYLfMNJQbiGh9g3MKfV0gfrcZe0l2w7k1F7+LZzK8Lm6dBq
UklGUrSMMjBQ9kW+ZVkUDyyvW923JrrHXkfHA3aKedw/2bGmJL1eDUA/ds9IkEMiQ4ghe18Kp7EW
Jm879Kt75/FGR3cHRSDGN0UjNu5++XTYWQQlU/67zoSzLpAW9iUyeOVB+R2wpoV2FS/PysFIboQy
1CXApWXnDRuDD/gyTomzWQ7gqUgTlYQUINUvvDCSJCH3JLZjHgYX7/j566Y26hOPWxMEHvuFvnxi
ZQNq43LGIUOK84z+ew0AWy54VYqvR9do2FtmtAixXuqSZCNXQaSHrvI2yKzBXNZWp6tsGih7cV1G
ZjDhWI/a5R5LnPEBNV3HNIHw11/lAvMHvOx0PYEKXuAnObJucgTGISdwDTHxhwO84TCHEm3bJHxo
p1jzo6ml+4IwXslNj2fV1vkExX04Jg9qQ2kv+YttKaBVqT2YVmvpAdTbd8MUhgxfak1plshFadp0
BUiWo/y/ytOstZD+WuJhTRuHUxEvap/UDNncEsB+nkdOoJbXKYniydLZivkEGR8LUNnAgSnWScA8
NxITNKFs9WI5DABrw3trebUsQt1PqGrT2wOtNELMZI+D/o35sVbm++zzDzYNCl3++EkQVmCNBFYY
xbTGYE4EwKNp4BWOXWsdLx53AZ3mfRvKt0JgNZ5MoMEa3N/OECnlX8DP0HQhs/k4NeQDrWQZfu3r
GzLXUcxbKEGlD6/b4uEUhk+iJsWmSZJJbQ8HJtmxbgIgo9VTlGLOGBq9jzLSaj787bu4IM/PmeiI
qB8ADPbG85I610E7iwZnDZuVJHaxoOb4xwBEBK0VHcj7+XSnoNtQ2A9GQCI2cEOtxwIquzy1v49Y
o1gqdCAZ37wPBQujv8Ba86qVRWcMLmK2Zzj5EHeoyx3fm6Gq9lfRNGoLKB6gpHCr75X5a2jozIgP
9hVKyZwzDC73T/wBOktyEEQKAm1Z+AtnZo8002MLpfIDOb1fu/ePf334jIGUaGFhkdL2t3GXnP1V
gV8ock4O8QJezRuuZSDxFTtpAwQwWe2QAdMicJsk9BlVDNS8v1rfZEG9+BVSBG4oFdvdavrFlr6N
hnmGcT1Vp9PJkQ+GQck2H0sFpqLq7/iNBevVNd+RCcz9ytJjs70/ox4/TDNhbvr93cBOmmqm39Mu
9YNMMDMLOzkuRo9u7L52fZJxFhQB1qBUUZIRBiJJEY5LIyNRrLZtyPvjo2EPSjO2e+dmgawVgrho
KDduYTkNJ3j6sQoLQtGQgnVoBMuwYZAYL85SydljIqg360p8PnPepsLEVVXWiDZZicNMObJ8b7Jl
+hqjOJoe0TZu9lMsja742mkLF9iusXE+S/vWSeV+O+N8i+q9WWPjQmAThUCU+laIL7gecBp+vEAy
rj37CaStc2+rTw/uSdXJ3jbllbzC4++mvlYLKJLAlWnHVJDID3+wxwolqtbD4/btAqezPhTlavNM
Osmea4Bk1i2ifj8c49mX5DaPiOOU8zlusFvfPXt9llXpJ09WoJSi9dAV9iVmm9YfA2i6VVUNOpki
UGactsSaexfqh9Lob49oXN8C8+a6SkAvi93tNTeIVZTKjGlQhdGcEuIqZbs5ULbTFfvvtfyZc+ks
HgxfoL/nY3tNxxKHinp46+ykdVDEZ/8/FoEVGSxBxqpGakOWbvGHtx7mFKBBwp/FchyvTLWVJOJp
uXHy56S/14JD0uBLK33ACVHJcamYKlec1gBeIQ9J3yrRtqLcjdkXnYVutlvr9PRvE9FjMcN5iUdl
UT+rDpFtswe8lrCFbSfxZDq9ACYHs8FhfX1NqrZJHtqdBz6vCCQnHxA5DrnB1GDB3JoELWbK6E+v
DEIZsLPUpjR9aEX3pjgsWirDMo6VCYlOXvPA1WkVyjLOMkEqPIJ9vxITpy+uPoK9JitPaT/9RqdZ
rAHqNQGbRZUmK0WlnXNcQCClBZp01Pq8U98p5oqqXLk67PSezKB8SfiLfTniWv+Tq1YLkD0i9Nb2
ylINkAMJiwrdDd/K9BFLlBg6eFTcxJuBxySd7qjOvY9Dvr5Pz0nlDC9aFYqu0uYoioyq9c+05rkA
xGgtm48t0487rG7RGdzNOMySeKIsYaOYeRjtOK+dsqFYB2JGmUuxY9Gf1yGMnjO6KMmQYEIJF2lQ
UfV21OprHPFdKBQD+C19hqUWO7tlWVjGPaKs8rOkPIf2WGAill0M0sHrGM6c7Q5UT/xpB0crQvd4
UkCZkYkFQQZJV/kyzP0ch/qXT1o4l5oCkwus1OYKu1+vhckLTCCvEUhQdYZrvHTUvGr9t/sveV+7
oSVvpH22Rlpr0avuVO4XcetEFaggaST5U4MFhixyqE3l9gJPL3HmC+lnv64Qc4Urw21dyPLPtIcs
tcpWPyo8TsPjFBue9uzfe2WfiXTaa4Pfw+W5xrVArL+IkdUfU4qudxfDFYvf8Ci6ro/1w5reFGdy
kJZIGeYXeeE+km/AXOLn2AeqVBeV1CDL+BiTEdKrN/1gV5jVYEQOLZxAA8VlCkZw/UTLFlrMwwyv
rx+yAh8fLvTqDrHQocGufn55+BZdVr2dlFeJd6QWvCvJ6JhUBqVxj3MjU4qX1jr9wRoDeI510jSE
Pfr9GNyH5tbSECTZo5C3+n5cz6mPutFrSMgD7usOfnJlRub92ujpLjBbVzE35+8MlBnUel+iaFWo
Y8/CN+IwlouLYJT3qKH2ZwoP6LShGv+Amr/erRIQWJTslSiRCCeBEGEeNR4LSDo9QHVzqZdclU0p
XCmN17y9a6urd6Lf9oDRFxSxAakzQb7GzPFNUYdt/PWg6l7NwR5GihICwEHw9PxOFk+rKBz+8v10
X6fodeo6ONZJ4XSYXFSwNcpZMUIcOlrT6W9vLWtoYhR93fRMXekMYKAoi6vm3tllJzmSCOUysCME
NwuwvHf80j5f0H2hu3DwmjYK6pu4+BvL0bmcTVpm0MUspD2DMfcn+6n31Ve1upkGzt2kZJJUVAjb
16o8LonR9Rc5h6Q/Edd1V4BS8BaBTgnGR/g8YRwyYdlNGdhrrTfFtBQhDS9LEHJbdqW/B137N0dy
+Ixlg1N6zLg6orNrWd9zW6t+ulBfDKM/xeRQgdgrwNzf+f6NLLK7F7RSRYFrf9uipBtlEoPbycP5
ZkQoESbSAB+7uAON6qCF8jtJ/z1X/2appk4BYgBzrXhq2lweFWR0Ev8cZP+NH+h6HeDKOePqV2hu
7+qbvRBmB0bJiYeZDpHXTi/8Cb1GiuV8zRqDOHxxu0ixnc5szNm3JIk7Am8TUed4AVKj8OUSfk0C
UI7bmzxyfbVE+GKbusGljZWFY0qz+BeOnyb0E/gsnRx4l823J8CVjhMfap4RlF6GRTN027163nBT
2mXf7dgXArv60qQGQ/ZhUpOtiQ4msGcdvy3GjUG4s1dnzGzvrQv/AjDc09i72XW5QsI6TsvjaJp+
NDD3ddug2sFtppRf1PcHC9kyb2bkH8yCoLHGVJKtvrwBGW9tXe0CxX97uMfwiKDUCo4WUL77yYOJ
hNU49bPis58EolkmvFHFlq11Us9iEyF7cvdVoYt3UKCeJ9Y/JJWfKqJpc0u5wKbavuSOn/Ew90nI
AFuv1Fqixxsqx8teHRagcVjEi2D771WRfJ5DjC0z532Kar+ZiHawmX82QBSULVivNHTMrnhOqGK3
NiFkuqLEyPV2G8mImtHkJTym3r6i/XdrAhgPHDGGcJWYzgN/wZbgnTEAbKpilcCdlAEcL9lHt2yk
emxpMfRrikRYlEuAFLtVwK2vgKCiaHO5IkGdKy0dk8Nq4V+sXKf+HYKukEzcnKJEe+MSLoptugdR
/1PDqNCmPTfQsmHZbkxuLqMaV+NLzdfKD+/V9StwziPPbYS7wXp7GGo/yBrVb99w6sW/RYqDiP13
RadVeViFR2BxekNGyN6MxNvOXQfrs8bPW0EGYbQpD5hgNk5oY+KPD4kUp2zT7t3oxnGZvPQxuclh
rxP0vUvwFZ5jsDFET70srm5BvLCMgu9xnScMxtgIWo0bJk5Uom+Eif/Ddy0hdBluHODj+gXUf0pb
klId6nyGn2kaLGltZU/aEm7D1xnxk5rjYEPwGFHVH7QKVW6wWP/IRj4W0xToGw3iynXyO6aLoeZM
s/IvYFtIZ/3k0vVLHTXgUBPd1C0hkVhNAd9frzaM5Ulf/qWTtqlm9h68xRgllCTnZQQccN8w0d6O
vSyHDQ90sDqgdGiRbSEcfZA2OMVwi5fa6M39pk124qPK4MGB+xBGZ9iQ6fUxtxkuMrZp2nlu4hVn
pbnwJKfdpDjrcxaWn+3o0r70PFH0e3pO3ywUSfizUOWmIG4oW9/80T5nwruWfqDiBVn4vRgmLxve
uKdxMZBJgb1rZ0df3k9/jRSlYQyajeU6iRNCelBw2dyRoeC0rKfzedCmJkPl5AY2XnPRyNNAcTYC
3V171FD23B/X1KM2iFgT1T+2ok7OwLhrHIV2wQiHlyVmPHENs3WtJcPi1DqqR7djxXGmnNCgriHH
oJDozNGG2heH+3ry3nljeMqr5Bt0xw/XabCaAwaNOl6/LZTXlC55Br9oxtWhm3ynf5+/D/GjAty/
Ombx2121OLlHgWXGXkraH9JPUElRGL13y31TRG9Jh4Jsn07ln3UbzET7MRw3TNkj8CT62zZfTZ6q
J6s13/2PF8gDdSve0wtxv3eX2tOgDu4tqXaSAFUIy3zAJP5PONf9UsmAaWNm+CjPphQCV74NONR5
YaiafHywCiOujP4AuZNwAPXdSB9Tx54JC0OJCo2LtEpCARVahRNq/xwjGwf7LTAwJNiagZ2v3S/O
hhsiXEp5poE6yDzJ1w1aXMYHYpIOoAeqlZvzE4A1En4rq8a6ZYHMcSwK88Za5aCfmBrUpjBocuYL
/x/1xx7XB1DzX2mqdkd+1z+rnbgJS1sNFlXdXtWJaYwcprTYORDvv2/Yzhv0DACVXa/XaNq020WX
AnKxSlmKh/cPdIW+cUYNjqXJsnwbMUIn8nZS+aqwf/W+9lUDukoQv3fph8BeLnRLdfbjSwbwpUxw
aiHuSdS/4jBYmt/ZSMFgKoHA4Xq+HbQbg2ahUZc3U7psDSkG7q09MYU7BOaXCGQVkG24NyT26R91
L6F25ARlRVVFV3j4afjpH8xR4y1/sw+Yq3eiQ6aaV1D76d8LLaMdnto3twsJkYgHc2KOJgpeq1e/
nZc7eDwn5glHU2ipp0oZ9cIRqbbmCJDiAKXXYtdqPZZs75iQLOQaUj8udYovJPMRYITHmftZpLQ5
qLbgP7RStAlMPvxMbVCPsJ/T1JPct92PACn4R4O8+BFKT2DfTzCrg9T/ICpbIU7e7zep6sQzZUQx
nAvOY4Utqv+DUavdd+4KgpB9MWybdj8OicbyAUKKi1CVh00CIUCMlO/6mHCcOis1qwXaewFzqgwW
kW2lPgHwrMj2vZpIcWkGZYEZikweWFsROxchM6unVGPwdem6grqRupkCahnfvy0I2vw8mLMFTqqP
QjOJsAcexzHqy8u98VRacnvVB3bnK61Iva6SBkvGj9JhDhPfzaS9N0GFxLcm1x6ug9UBi/p7gz9F
+UJ5Ox+ROj/ntiGTODHVMXM3LPFtJxSU5Glul3vgkfhIHBJAb2piraNYuwQF7n37plbILunf0sWb
2qrzGVyH1ieZUXteD1Hmg3S+6DAoXoBqD4gzqFCh8IfahXsA8E7xtu27U1XsRwgFwNCJawaWJ9ny
tIKAjq0WmRTXgSl+gxDByxXO8lIOo+6Ps1NmIV6d4ITDnXdTYs6MGinEjMn+D5M0dL4AUFSsl3dI
O8Qp0qk1Mup5QsuEki/Kl6MO3Qy3Dm3bLfYVaUmTDAcF44Vj3cxB/E97WfCCCHhyae8BwCplcNax
BtsKoGEuoYY0UhuXP8KM8gvNDXiviXAELEiWSJmpGMpfn9sh0g744ypckwiuxcA7XYMRThsttmjb
dai9sCAMzHhRU+96Y+ljpSNHVC9sJgQDwrpPAY+N6rSAAHW0a+BTRQWyYs7jkbIVkBC9wCmyityQ
BrW6GWdnIyuNZqN4Rct7KU5pt8j8WNT4cUN2CSUSo6RnioHYP/faJbOj6BYXL7MR0FTdK7T1RQ0P
+Tt61UtLEZ11fZLgne+TDEFXrXjps0iTAfqMziFaZRWPpcxonc/fZYCaigBtwZ8lTvQAhTZCybeL
7lGfRfMCwffKhspgB6NsZzDSgMCelV6YRec4UED/6r/0YblnhNQlpEJNe76gQZoeQRgiRd3ETKtt
lh5cxkWS9skjKeYqqavmKZyUZ2OM/0xAF3OZcJx6XSV+9xW7GCozVmPw6n9U+XPN9eKbN58WSzgb
43gyfNdLJll/RJbmzAEkTgfBhxF9WhrHmUR6gfw1Dt63FhvsiNF6Jz9Qq+Jp0tOwaw76HLwUArJF
gCBAa0Bu/JBS9ToG4b7dVTBmgG4tamJn9tREg5XAFZXnemZDqgqInPltCLmxst9z+mMHG/Xti5lO
2z7ySBmgCLYPCaDbkx22S0rrQF6aV0Ms/W+JLDyMiDv5LfhUkvY1U55VPectqladFTVu24xk4g4y
I/ZanxZd+WRhw/kDcXngykvG77vVWK+ak/yIclA9uRMnvpCqnC1m64rf1lNQF234pAK3QQNmxSvP
Y7dGo1KuqYDYh4R1QA5yoNVwSxv26Yn28pIE04IY6YezA0UYkbyx/bw+BMKS9TfBYbSPFeuvLYs8
zg/uoaVtxiBJgv4ugmPPzznlhEEMzev3hqxjMZJ/BvJNzyupMsef28f3dpk/cSgiwAUIB65kCAdv
NURAH1EuSu7ac6nM/KDleCkNRpAhFvS+AfYroVGLWhfAXHq1d9PXFsypubCNhKLZdjjy0h7/FCHK
aZXCynpN+4LFIaf+11aN7WxXqnCjTPsYEWFo75BsRX+CRIPpPVoUzNneR+ribMA25ZR9aetON7gF
Fl62O2KxsW52xdAxJUxN1A/FxcYkmCmBxv74AaQSgOc2Z1KUEFNtRh56rHxeQAlAQfPpFUY3lS3r
2vkNBQl6kzOiBbec/EeBQsIn6t+yChuXQE9z4FioHG5xpeihfwYUFmsx73klxJlhVnBA9YcFzpXN
hF5cf3+KY6ZaUVJe3NqELLg5q53lZT5JfdzSY6QpIdAV9dcx2k/nRhYDBd/apn7Dw7usyzT7FCCZ
8HuvowaRcF9/AwmsmdjXCviK6VJo2ksbNejN/rfVVjsVkF1MaHcd88BbK+VSjIuSMtHesrbzbG5b
ZuITk9lDt/5v34tKb1fvHZ6lDdgz1ArJj52OluLVbyoIUqTzaPfIEtiXPLN+cQUq19GPenKseM+i
zAAn7Al9YVWeVqczU/cd6Z648rN+lvw1PoSrimoeR9Hc/TwVwYIlkBYgYFcpwykjvPv7/01m7XLy
2HWuelynVxCJSRV66hylng7FK4ez7q2pVGQag6/opyFdF93IWAluZHHG5fYcv6leVzoXZylxJOCi
sfmx18/PeFKBmMc1xLvT7LXChVDoIcVT6XrraWwu6otjW+gKB8OUixiehUsU4BpeXuBFp/0lw5Fh
m2Gn/oCvaZJNdS8oq/iDDSqKcxlnizjxjwH5Ems6CiQrU9zmsZyDJzNi/VNcmXvWos4JeB+aXWHI
mQkyJ6/SMr8koJcbaz9ZZPOCKrWKm4Bs/Wb8QxznofoYWqHhE94+JtMAU26WOg0l96yzQmu0thBE
G/oSJb3FCuY7ZLs/oZRzhe/fMUFYWEMuLwGo/0lvFY11+7CYL255LvcDhXRkVdQd45gqYD7AvLwi
pN35Je1GQYtW/rMP7DsY9zrUHYLXoUpm5LD3fFz/6YRYEcwHbFjSpp7SWrEG7onPl+gOktG8lhkg
fIv8NK4CdaMb3IdzOjVkr7/UHm2XxU43v+7O5jQcNmbW2yYpN5t3H+94Iq7LyeAvaAMrep2lydly
JL18l0d8nPwos1hyLW0MiT7VwYeshwlLsfpe+vZtKZQlQjBOQlegbfA+k3nKa++RKFEQB5R9dsU/
HcyVQHR8CVP6kz+PwRhy36UcpOPNrHjQHM3ic4H5HiUfEWkeAKDs8xBUV7flFHKSjr51sVhoDL0e
lUvXQA5GoVZoGKhhU5l7nyVtlkf6057a+2MWesyW+uVkbBqyC4plAHQkRftNcXy1yaxqh2vTwO2c
4LtKOLXV0YOTigO1jJC7DsOYCGBGQfq/cPXWC22oW1P28deb5aEjTy0DuCSoJVmGnKDuOphXxCtF
BVQ9N8vMA6eIr8YwyKHb6UtPjJIeyilQWZm1pO+WMdIgkd7UaiE77ZbDIWyvutvJxpTG9EZEnhtD
Zu2oueJcbwTbXPWIVHKS1wjKZm5OQXku7ppfH1yhCu0F8pkr8fkmpyxvv4DAucpbVeWj04N9ZIdY
bNGhOOMVA4pWu5ys6pYakcVW8+pn7NmtvZ1pVkVe7fmlYvdOk9spqQp66VEgVhBdL1La1ljFKNvK
fCyOPsBclifddf7/I9GjrnI7BNS8bpIGCkQTN8hgwIWR5x3MWYq9ZO8fN4l1lBsIWBeWFGbebjj2
AwKg3E8+LpDb3p7rhR4va2Y/lZQQQ12uJKUhVkfxfJCHopf6YW5Iu9YRXtKzRXlttnM1W2b3Y7Js
YImXOg1YhVoDOHRjusduNikEhim04rMW0At8MODdw4nwEiLDmjMO/Ai/AO3x/WZ4Pskfi22qO3qD
nRjR+MQRFtD/vdTuKG+TCJ48Wrk3VwtLhPql8oEufJtZGHrzmpSWgH9g4XZsLkq9xrlbu9Pr9u0G
HmOAAqqiIHiFUjqjPbzyOGY95KjGuxlxBRMOxeqCG/BU+iRLQgBZZ+Q22lCn9yC1hhrRHS5jCDdH
hbaYnUYEIFHiSHZX7DSdAJk84CmU96vyi+N3eLD/EXrRQcrRth4TVyZbumoImHqF9T5zzY4cgr8m
tU+S3ofNhs92MNSoITxo3CQWx+H8FsZJBL5fcfmR+VxO2nyOSOsd+Ucl0wP6dt5JvJYbWA0Y8/T4
m9VqGHoNMVT2zudS8G5ukBwrJb70JuIvWUgB4GWn149jMaiNjfzVKlYpEJN2nfhXVzr6inwdIBWs
rB4EBI5djIqoPuY+IK42n8goYeWQV044/WzCEA+QpUtgRno8HbdENAfK7KkdULeFC7UbwEDRvLdX
IlXyx6BT1oeIgnFgRAigbInn5K6f1Gyhd8ZFFOx+9k9+xDfcKPhfec+kx6d8AdWmfHpZKlAlL7C5
YAHH9vrf4yH9GBkoi64OrXuETqQv54m6g8ANtETkAIUPHTtf5JKyFiiqeZn0ZkwLJxiuOFz6ynHK
P3y/2Qy38ffmuDPjt1EJ8L2V5tCJF34wnaSSIjmLRrjUGw1OQnrw3YKEUgQGeNXBudP36AQ9Qpcl
6cp69z+abgl/U0a0MirAXw28QFTXjRvQQWjxKtrNV0oagNKGCNNi8kfxJ4bhkqHZ8+Muzr/kO8xM
Ys5UiPjdT1U70Kl2R7f3GywGcpSxkPkffLCNDHEnzg26C1z3QpR0vM9CbVMcMAkjdQvi2n0FiP6/
UFiUY5DLgx5WqUvW+DXB9BBAtenQfzN3lEeevrCPqwsZ/unHTI4u8yBxOllwQ+qJsf5Ok/wxmX0l
rYRwe9wu7PIFmNZB4ab4hsJWWT3BouulQLipY4SJnxrHjOboZFEOyv+wAfKWzbrus2RfPWLFxHtZ
JSIohR3z5jynNgdKjMBeywFiwdRgzwfPKJCzEotORorRvHBqsipPHBj46CINbhFNOKSkUzmoeR8l
ULpMPEJL0MzasbQdcLiz7/3zuqOvKiAr/EzU6SQ+K5DhJY/CFONhNkh41t1vmuQLFsl2F3jBBfte
vy5BNFh6QqvheBPok7vZH32iOHIdJBcxld0Kd3bFDI3+hIRqivPjCeCtbvR5IA6loCUopGCIHyoO
N51n58UXdpPTKV0jVPzJNdhOeL1inTQiiaKUL47FT/v9RsVeUlQoa4J0ZZMeTRHxE67DiLmLMwKj
Ffu6AfEccom66H5Mjqe1LMyd9V/cYk60nKfU9zABi75bvN3b6oIGH84pOXS+FHIJ64njQeH3yVR6
TbBHdlLAbhRt7W2ZWuk1l6m5KtxQzFi72dL1oW1fKhO1uWKRHp7UzQ7KCdAuuqu+i/+VleGcMDxP
gMlAqGF+KRk67qX5N0caEREa/BTWRuc6bC0W9poAkb4PetxbHANjqOPs3/vaiAg/2MSX1xU7zFKq
w2cRsOiRNML7vsQY1kYsjpvzqWLuZmkjsdZmR5DOJXnZUSeUOVveoTszRqksAScYIDLwjAFcFLTX
UE6ixRP932AKgtaGbPwlnvnx/aG71vXAeL5ksg0NO2zCaOJNt6Ill4BIT1MI7SENenkNvxSA8zOV
9hlPZfqsblQZmh+9j9VxfHCoNCh0IuXxZug/5CwZHR7jKqwVzBAVgedYltWpeEXlytsdwVY3Wc5o
tdc/mWlz1wip9U0PBoI7J5YSVFQuuRrT3ScnQqBSoZauY2eGP9zmBbLO444b5fL5h74SNb3rJdW7
+yvhKlE/RfwEjNYO2Q8ztIbyI/QXlT5VlK11S/wxsI6qO+m+TBO9akB20JWWJBrHzgbbEtG7Y+4X
Aq0wA1eS9h3zBYayl5ss8wOukEMmhSQ3F5sU7vdTM+RgmHhPoF5Pui2nir2dgGC1Pu7UEud2wKz7
x2T4BFiFTp1LLgsiy400Dwztds2Lhy/nCp4SfMStYaB5OUay37RDB7ZJj57+JvzS2xfOzfjYzcVB
hrEvDocbB1+qfq9NzpZadXuQfsvwCthjwpkcYYt2CEgluYtJi/qI5va9t5vzsgGEqbHVm9jj4V/D
Kky6vNJ0IbsAQsgeXiurbEPlggQsqjiKIlkVutAizubWTQS2mtxix6GWxwhmT6+nH79Po7iqEz8Q
NTq78wkYEMjxeofIkhu+tPhiYcWH2JQcDBwPpPllrI41Gcr5V8zmuM9T2rhu1NfLMikKlRlyXGb6
+rdUg4OYqa6FDnvN1BfS/p0t4ko2lwmqMuaMKAylZbGxqwsGt8uBbAfK/p8B42LLlxt7WjlsWXK9
oSRQIuZ5aKZ62/Jie0ELJv97FwaiRXSx5tMTjbXcvryZ9+j6Dm6YYYBDuyS0+OYCWaJj2avstbgE
XTcGCX4aZodwuH9cxpKotyzur2MEqqflkMuxelQ3cIbTN5d8BPXUs9KNIQZILQGh/sWXhEvNXuZG
m/XgeoP+WRAEo5dIJd81T+gcr5WowbaYHbz0jHNNCZzuEWYamcLXe1JUrK7wAZ953Z7Q+o9vRghe
0C93/sknqDy6R4/6lcfpDGA7O7djy6s4JAwd56bdsuimi0g6gfvJ+yd3BCHO7QpSZh9DEjNiIjFN
W40lpc4qej/+3LvoGq5F9roai9FbhUWFvoN11u4j0E1cOw9r668nQ8r6BzpS2oyv6z/mSEdWwM+k
lg0xfwQtqbvI87UlC08y4LFTdOFEju4bKmMsk+TGzAFgaF/yBN1KtVuwSWrTNpsLgXh78QqJQoTO
VKS9sE8PJQQIW6ec5bx1n3U29MAyqkD/szuo9NZeuEMcEPjQ6LxTn+Xot2b/mZklkfCaFwGJMgcg
w9rJAy2wQFLWH3b6YD6AIJBdLx9iOfkFMhf99wpES4/I9c5ZQXN4q9VvqZq/GB2edTJHP8jbF+Q2
oLpA1GKmzlIW7zB3OP92ZAfteVWcpoA+f7glb4Xh3GPW71MssVCnLFt3H19j+vc3JHQrC+rJ7sDE
q3OIH3CQtdOUQfDPlRTim9R0wMSWmzk1BnKK6DdOBchMFDgqCvhwcUCK2tSYBjOQEuVtU6aZq1Qk
bKcQQUhqUa5fRwUEX4BebxCh846u2Pkl/cghXcjjWi0oX0Y5GUb4+dlEDUYx86MwWNQrdVVWRivP
WHTaTxrJ7W1TShZyHz881gUm5alXfx2UwWxkReB4bwM6D0u3PTG/t64MB4lbqwSzNumis9w6uURN
FS9KS98uNgB0aBssHtvz2+ns+fR5ztNpxtDURsqwMc7xon/UWgqt6289jkYge116Bvm9Bz29QNhv
y4QCh9m6WJQ/evext4EzGQlkPBZ6WEu+4kcoNZic0a4ZaNWF5z78WcwarIWPBMXJE4AbuL4+5ngN
sAfUWa4Hg1OePL3hWTx6iM7T2nEgJezyBp5+kQ8O8nu8EsipwH5YUBkMLkwiDg+5eB4jKwqpoHQy
Mo5aj0mEpdZ7rkJzRJAP2VbcfoEgWG8C2djpJ9pwlFkoD5CxxyGPTA6JC287QBjM0knkcXG31Jep
PAVcQCJDPjXhbVVWjf9VFJCFmpfjbk1DCp0DjNnCwo6iF5H+i9lnitgnJDiY2+/RsIDn/j7C6LHc
ODV5ninfcxXty9216lRXhi5BzjaPYo+gTyj2l71JufVzWS/efkaOb93uRmZ9dZEb+fu9qjD8V7uN
QpmJatcP/Ht1ymI3bC5vglNp9y9w2FYgb3oh8DohW4zqxwUx5OSvWQ1SR/H5NEoWyFecuHvsvF0W
l62YfiysAnKq2etUraeLnVMoFwNBMsm55Y4Gc1BysvDYizsh6KmLMYmyyr4SfzEkAEvMO80w1C1i
h8BryMO+lz3K4nzXshrWHZslDmDy2etdj/nC0ouX1v3JFsUUxpchnBuMtylp6ZgKQTK3I04jKfSW
O04IfEk+eeqUDXUEM8McyK71hgDz0sSbHoy3euU3Uyk2qT3QC1mhMIo9SxOstKF09rThriLZ6RUo
rr2Cdvby1qamWgqgdo2yxtZMjeCeTJcsCGPVSDNLltzQQUZ9FGFEooX47J1t7J5tzK9MQK3/jxMR
+IbQdWEX4fCAcppSdBILwXQiQtsTTQHVqfJzmMwds8MxbqKkOQI2fDkk3rtJnA7iF63EIgNBCk+4
EXuQpvNU73WEWcI+v3AtPY9AI3/kw+UJpdXXpbzYGFnvU9JS/1Xdzi/PrWyb4UZmKWssE3wxEvqy
Qd32wG1KvVBlG9BgHLuPiQfL3vDMqeGaey6PHJFdjdMwNuHcNujARkNiY3rKohtajK8JtG4iaDZN
jARwWteQwd9GJEvN3oyovRMwYJM97EcncQpTDHccP2NTO3K6JR9IdSfJMqWYQAES1twc9pDvFxld
B2mmZ9waWrlQo3BdxjhYeoyg0NcpxfgTuRqdjKbm7MHJNjGdLVZ5capxNAFOU53LGO3Dby2U20jx
GG/CoE3sI62sYxE036g1TLDbfk7jfUe2hJdmr8X9XqZdAxWC+p1SYAC5iUjhSPvzVWU/rdHCFmet
SlKVbivKvCv8+lfKalJX5/LONmvM2O93mNMYmcgoAeKlC8h99a4+CQ9T2y9z5xyI7x+edOrC5osO
MmDzsmHziz2gNuXCgqMiVFIupdYazCN0W8fLcpSshcxdR48SGjc42b9eFcxNHmRMbUF2GJh9nzxA
p7kPjsqoazxJo4qxRrx9myPUqBIEF8iHfX8TxX04vIHmqIjUUrDPkq1JenJFpdWnaQPfULFiCkjV
4bNldaHTMvoCUMAAiKVn6X2ecpCNAS4ZqWeP0H83KEGjmsggHhcmoV0+wLYpdYG+F72rjUreHe7z
3xYtmIpsQjVO4WKtncqlIHyVsSolQzOQ5QY3UVQhM0vjnEz50AjWtnoMwD5efYWwZuyQIxqlqHup
6o5EiI1dZcXQ7vk3QToHFFqHPlsVzvzelk6k4ZRe1GHdi4feaJA+nAdDML5Rk1mNQ2tjyYD/8Lyn
JfqkEI0Q3L2Rb4wsRSxkkW3A7dGA/8hEx5MGh9Hkibtl/EtL14yb+XpfUuWvZhYKFFOCzo8WhD1y
IFjIBax3+BI9ujqmWGSmTW95CvENrE7+DEeekLLP5dIxOTdlAvvG0fq81Cq8Tqfrl/q9bDLRTxhe
QLKyDTj4nAOnMCshmqpNQsnQTXcp9sXsBu5KiLG1ixcaN02Ns9HbCbvfmT/L3CSuLIhJmSpekMkG
gCicVO+x/JVz6RirUwVCG9KFoqqd+eQ/bCzoPdefIMScdvuToIkdWf2+gSrqQnvx7BHwq1Uts0e+
gs39LUEwTpkOV8mLyPpM7sdQ9IV0UhJDPI5xQ/mPqRRZgsCteqXkSimfd8sx7XaY4f8aTn3MdzZq
4KbrfJ7Zp9a1zZW4kPSJo5GOQA3pAW87ilBocwx0gZ/NtrOA5OPTK7LnqwsdTtfX0276Egh/6pSc
Jb/j0Tgw+I9h2SSkffE3pYZ984jlfafwTx2z/KF0czWekEXwgUzqnYTQFREH2eV841wC3dxN3qFT
NYeyhfb1lyQyUYaTxB8SqcuuMY70+guQ6zzmmqKaRz4rvUq4YuPcS4iBhzTQSw9hJKFcAg7MCHLK
meTPMyenEmOnQI6ExinLWx8G4xNdh+jgad+dm/ffaK595yvhYTJfwDCsmM3IaxPZD6JggIz7ysP0
GMKAgD++4oKmrUoPOADqVdzwQyyJlbpw+NU0oHV3WZkFxXLgWBp69EERjzhteo7XnrmDCq9xqHYf
yYbNtHDLN8RomNVomBHw9pTFzsRgvCF078pYKO04j5xk25vju42aWQbPTHZ6N0CiEDJmujFhnsdm
gdAVQn0XjJLudL/5gfwQ0NW4sfSJYwrhZhbTi/QQU/UZ83GbMWFI+aILoAliEJK7z/AMN99r1gUP
FNHiMD5BKArIk+FaSr8q6rtwtRP6W0HG13mfXavwSsASZuWvDhr+STQfCuRWUv6rFBURgnkXpcSQ
HQUbAlE6pc/qAvkHv8TG92uyBarnB+zKuCDaetHNIowYsBmQXHuk1d+TmXZSYJAOr6xbanDqO4Jx
btY4G36Y+ae/crfFv/md1LPOlKu8VAGY0DOnmgnzeqPsexFTOwElQ9HPelkNqdZ4/icU+MJelUcy
OgfGdcMMgvP4XTlEpJCs1PlkEyzU+Hg1Om+8+V6jFDf2+ECWIuSZMP2cEdln73dSOfKWAEjGC74X
cfRXtso4Vbfi+kLZN1qR7jl4q22yJG4VxLpcj+TFnWv5Td3IugVpT6XfDPLDGzBkYqT+MApJMQkV
noAQA7YGaftHqk06Fv7LiE5BNJSaqpApSELw0mdhT2AIdTymvp1I6Gs5sJvbT7gMJGP5H86AK+BC
dP/++iUEwtBJFgTuMTJ6upbJUrGH/LGlzCCAfaWcZlkC04L6Yd9HQS6QDF82N81AH4ftB8uw6JZ6
ni+Kaaz2WxJ00J65hxqyz8djH+me+GabOQnhv4ppulwb5LVH4TNekKqlq52p/OFDhAHurkm0tjSK
qOEmNAX+0AQ/P0nUAM/hL57fN9O0WLyWfze9ZSth8sa3rlqQNb99lKzOw8gM8/i5vodqn2UwHmKH
oASWry9CT9rkMqt5eaCKQY7vRKEgROWu17u+RjOPLudYTjPtVINClajEmFXFhnZLc6aDi7V6hsWo
Aru6PW9/Kc10PQCeIQdq3ZEow1/P0O5KcUy9QIq1SBvkR+ONeg92vmmbrAr+qWTTUda+ISO/rtmK
JhmT4fiP9WlMwaVd8JkdJwLj6Elm7Ne80Xtg0X4bGhOtTtyxOgByNYDrgXLhbs1HnY+zYt7XI9FQ
9U3yHzXGKMi9Eh3n6ps/1XLobLK2xO0COCQA7+OnQ8r45+/S+9Mtu0CDi28lrasoyUCH32FJTSWV
CCp7kAGzFO66AROGIIzwN/h+pQrOJ6i0cIVeQ0xbwG/MaRf1bfjSTJjcH7XXXPp0SNI+2Hpsx7tV
yzXulZr6Gu5Lw4/BXZ0FM9zKvB9n6bbhNhq9KmW8+L2x6XAy8um7fkMFkvJTrgfJNHwocLSKG3VS
ns5EjqkCRPL6kkj9j7EXpSx4CCkWKJos3GfIklAgD+mySLpqqA2NWubvZhET32v1UeprDnAXSE36
xteOJpS/Itjnto78sEz6n4U3LiilNF1KOlTyWul/pGCvryEfLkSr7qkqv5j2J8F6NBm7aGh4Pn89
qftdJDyRsiMaY7R1JUMm7jXeIa7MmrynzNIkJIgq9V/BE6W+1iWD59qyiDGoejkJIFerA25pgfS3
W9MASZCv9FR0ch9s1lIJd/knP2lYPUADphJw9A0nWECuWI9rS3jXxKM0J721IZjzTEfsc5J+zkaJ
/z+FdV8pzy+PdZY9SFLUq/mjzDgDJy5I+Pbmr/a4d6PUt/G0HjneO8ux9KcaO2CgsTU9KKy0eEh4
B7eSpNNekwQV/gqnqASZahowG3RfyaiPm/Bl5XEs08Iarrjo3OOYjahK6RInW6ou5RMO42AxA7Yw
MW++JFMwO9OF860xqg9BAEiavdyMkmfgupmItt7dQOdR5dkUqMUaBU7Uw83DC2lNZ55Lqklxhzes
KhpF9RvQd2vZSaSB/VCblwIgnJ9DQE+MXoopSum64YPRL04XqbUSam67PBw4NeZRE3WdzEQVbjJX
B6ud1ye9Mga4ykWPcL/nV6TULsQTJJCvMw2wD5lu9AJ8DPBsZoPI4LAMwpFyuXaPlzdbzV3o1Yj4
G3GCc8XLvDctXVFsYD3nucmhSBNp5DDSCxPsLk67/MphzEOCIxThajgOtg1B0lw0huNBdX7wn0Z7
h+WKZH8QmkqPa6/Mf50tVXWhINxsPuTXfcmFKrMdP3Vvnyjxqv4UybIRtz3/Ftkd5TQ5NjadZGjC
osp72urZo11WXPXR9kkb1NsqrpFyehGS5oF//Sx5YDM32uMHLhBG/ZukFQXw/Fp0GlF4wzb32Cxc
rVbRReop0zb4kjDHLvwaZTPrj5b1UUnZUREgKaLQ2iOZ8buPjQle5K/+XwEljvi074cgTU4lqiMo
ykYQUl381Cy0fRZjEZUUbWNA7sGJigPvGw4s2TgJxTw/xCgNNS1qPS+qmc4H4gtRzicC7fy77rny
48sfCOIRKqU4h+Y+gtWrLMh8jihS8ODbjTmzrX+8h9v6Kym1mBsdjz8u8A++gT7gV2S/dzPAstkH
EBYmKzUnItpcnQLK3wwfkp3TJXb+mMlxOhKS8MnJux2mjMCYvku7YwEDTNa2C1vi2TtnD81VDrpg
/E8DUK+D0pC0C67AD6DSCov2oq/g1G/c/+Xx6Cw+JaYNVfzCcKIGrljOISYSrUgha1VOGvQmcm3T
rvaYcxAnfnKAyVnBoYRu5/auvyBinSM4j1/vl8LqbqMyf4p/iNFB3+tc9Rq5kYa4crxG05LUKQ3s
Z+Hs0LFVk6Y0ONkXYbyYNTghjrDEhXDKA1lMFVvfArcYiz+jNIFWcKozCyKkO4eEb3GK0g3z8jgD
3VGGU7uIjA2vKpxxFbLaXlyQrlz8OKqFKa1JBUC34aPHCixenLJ/oIq4D4bc1yV26Zzlk4XZTqGY
2gcNSin9KabOYrbuTHa/8MTBM8klvnvD/B4VJugnNgTruWJX/Ehw6SxwK397I4QCbmbLgDXCDAVK
QQB6vFGVG29DBxxpaWh5pbUPDluJZtaSftpu8/Tka6fg7eK5lM9l/tmGGmGR8w1JYmcuCG7IfpWb
1kJIdPzqs3C6XLdefi6k9m7SqtX6ds1yGW5Gh2GepOAwd00yjNqmG+zhXmpgOeZA6zgiwWPs5tcz
6b3CdGNS89WZ0APSOISqQIORotKSeBqhB9++wG035d8kiz0xkvuRpHxGqJq4EzKLHbcbI2aTc30x
LlxlsIBfp/y4X8NVxeWJplYvfYlykJbkcTvMVJU1rPEatL0FNaG3rnuXx/0TjvtAE7FN5ARtxVDU
SnuNI/3H28tYrBKbS5Acw4powkhRqVOvZOHA6vN2AWX4Cyx3TPMx1jUu/MpwZkN/CdLPadVKt9ci
kgL5YRXvPWJTvaWMRgErtiPGu2+IY7Kyy7M41rbgE7OPQRMBZKK73Sk+XQhf6pTDqDV3gtt9DE8f
5VMMTq42e9ea6VlTObocAMqcebROxs5NSt8e/zFyyBx4W3ykIw/CWgvpFAig8Xb+ZbGEF9XpKzD7
aS+5f7f/D6frSfvAgIWqyUR57RDWrp5uxIMfOrsa54wFO7zsY2UNaA7iJznjdBboJhaTuXEmODyn
BXs2SO43K0DcqKWvQHh4l8uMXMeoeXD9iAB84lCx9ldHjnH/YsbtSyNUjojHjDjWulhf+Q9kCaXH
p/nNXioYBqkrM81RMwmnzAlh1L0CG6PHturPZMRsZ1sg0HDSHuwR6bvOx+YXvHhhyiu2Dwtfui3i
rcXYW9o+uWk6m4CpO26aR0jdOV0ZhXeDHXgr2rPXsR8w+qpi2/Iurw+YtFkIQezMxpC1ADOFZ+X6
tSJaqo1en6QhHPpFajkaqDj1aTMN6cATvnV3QNYLpgLugTPVBAn147n9SKCGoGHHh+LYnJE0CWkg
IlntpNRhtZj483/aVS0sJoO2JxuKtM2Nd1N9qBzmkyRfABk57rHZ/9xWsIh8FdgvYGwwdam0ltwR
+t9Vrqma6hGjtiIx2kh7h/6bQE0jlVxDERb1YhuYrjrNbz61Q+JdLlGoaoJ+G/mqxfrdIL33KcyI
RC6Fx0TLwVb1YBgV1oqKMrIOQmtIAD/fWsJMcExEAHg2MbPDUXeDYvbqgY7KWhnXp3Tec8e826Dj
UvKnLKoe+esmppofouhVzRXUYAN9Rg5k2PIEJsPBI9xQwDGrl6m7AJ6BEwdoU6GkueK9wG24Prri
QhI+hD3QqV/9INzHoFvvkU6bhbW9kDJdBt0k2sOEBGt/byAQXxG/gfUxZyXdChKdbj35DUqudldI
Gvc7www4/a28EHtHIr2gpM/T0K66Vnqe4F3YaqqeWnMHcM9BrPPINxc2Z+Y1r5OliiGCmtgg8ohP
z0etaoS+s4hLD4kUlF+7ab85tMXV6yPa1KMIoqAIo6xGnFzqlVCjYvY2zjTv6FxOGzH/PHAeV3hg
ShtYJG4ObXa3A+vBA3jXfBcrTMKDXJLtgFoHfwd19s1Nxn6OMvZWx8dENneTsHNkK8vKVitt+Vco
Xaw01oKqBA435BJyp/yRY+VgVKJ94yP0uO5vwaiOOyCRZLy41LX1iirO55byoLVqQfJH1Nk0mkg8
NqJhvPQZI76jNZNY5NnQrkUeIENm0sZ+S3qihpzXCP2KqHD0t6dHcSATfxHlBfs4yE01kuul1vXM
1UsIs6PkwRkyxh6g8AdzixE1Ea8yg4vc/5IQoOU34AQiFKZsRJCUspUPLkr25Qb0vFe0wrhxIq+k
yf2nQXSFoiUQPBX/kU/lRIkOp/UTPBBGwrTE51zQfg+1y+pcxLI6sBdnEAmUJmhASGJJ0G38Ks2e
pxk9mSCcDiZ/q/iRC3AZ8to8kIAVoSCuqpT3sThEkAIKO+Qi/cdSGMwHxiR4+oC0zb9t2Ys3O7fk
GdMfFuApcJcXDVbm/zEh1Ia3fvf5MMYWuiI7PSkesvvxnyMusddXu00SN1QDmSMIHFPJKWAcvw8V
bzEuPUhM1F4uxKdarpx3rpbaWHDNX6bGHWHYBfI1o/GudDe6R3Q5ZaZYmDSQEsPmR6soUte0FLZA
3rcBsirgAcP7TACtXtPMaW4MAN6uHsAM6AEZ7eNpQysJId97AUsRcqLJcETC2WP2IbOP4ZqGz1jG
81JVeyqOVyfJ1YWFPbKh6MKkgKdOXb08nORwI1jfFkbKVD3ja+LFt6dqCINuT33ubu0sLEcfAQow
/X3o5Nk0d9hA++fSMjl0UZCfQ3e1h8WcTj40Lw69DrIEZSuFnkq8c6iDbzjP1LY59iJ/VfOHU/vw
yTIFwso4HKD1XUrauA4c9xZA3x0Uh9my94VATdAOED7kP1t0RTwLeSlx5rZy99Mm6TEkJxdVWROQ
IJSKcTA1ZSLsujyf7lHeLtx90Cy/iVnMf9DS9Mx+CTr60tfZcL8rDcPSmd3PhhL4SLBdxnoaRdF8
1marU7eghSJ827/RGTwU6BQv7UT7uY/Baz4l2+fMFO0QV+/wI/+AsYPXRESIymBghhoOKcBdgNW0
NpnvVbv+ht6W+qQwx0rHnZpTXhR7T/bb9E5BumG/jr+TecO/X+JhHAZwd/Ash4NT4HRZx4qsjsiR
r5Iv90hwnhpm/DOHEkiD+r9eyV0nm6flxQe8DCaD2IP8IcxHTDwRoWGSczdstLS28GK5MlaTUpG8
B1J7Wm5HGF0l5bbFJQ6GNLNzB6IvKgtUdj5Pc6KK4jAJGOpy59VKRE4ra0puxT8155X1WgXBGY+M
aUmLFxHJDaUB50J2x9Gf0V1su9RUWm62LHR57bynE032Gij1Sw4mo9feWApSJsJ06aKFPIcliMgN
G7vV1sUpzuHeKiEWiHiktUFqBmVjZXQUP33mgqw/YtREk/PA103r2PtYAp2HR794VLSOc5oPXw7E
AuG10o+4sIHcbIMmrRJivXo8W2ZSJrm+ALLYtNdQPWrHhjkxx5tUxXRJp1scBFlhd1zwligXD3OM
INvwBVfLBHFFsBXCa1JzO5uSzm7buQvCWMYzkUC7GvxRcoAJ+YXDj6ph+/pY9HxPoNXnK3Ibg2XW
bI1PRgVFYL8/n6BRKkB8p+b3ki8LhDjkFz2yBvp/MZo3lWbsiAPvsHCsRC3pWm9Z0qM+ncpyXnpF
wocTQvhijl7URT3mdUoFUFmV64roFIzqHnW9VBys/4FJxJUs1pexiTjVVqWXunLms9Bq2k719/W0
Tm0Z4jxX1WeDZNQ7SpqWXRdd794xsHNyHBvEbrzaKWP9srzSZB22BIngLXeC8aVzChmJANf8hmVx
2yUfeiAHaGmmvG8Mrozb2/+Yf1DM1rocwTcIQ316nj/F0PnA+RcByC5mYBGpLyzoCeIzgos4qj62
E0ek50Uz/GqOXwVZLdUrPT57X2OBh3W43F6ESp4+iPe+KNId4cMOdTA5k8ZF8rynPPA3ic3SKOAa
OZTHMqTn/+kdwOnyuO4Stc1DPC4tGlk7NMAxETtbLocFP7NMTrKp+lXCZzXupswwulEZ3KVfaNPV
Vx+3JxkHM9OeyXn7MEal9qhMxHIhxQKgsP1wzsClDaCQITdx5ws8vNGYV5xQcVKCH4txNO1Sv7gp
R8yo2wI8UGk2qNA0wqJjH95B8gMwJmIX2TwW3UJJpr8GshheXaD+w7whOcpJemIa/KDj4IjSTZ6w
2WJFcNWbfJcNhxhD7BQktIb0qVIKTerswiVR5Oa5o623HrhYdVHEZumZ/9zwCY4ikljCl2ropXbo
zQUlTyzJF5HV8DdYDHTYBhoWT9r1EkHIVgTYgrFn8nauZFOmqmF6/rPOTdUaI29vPkuEHfyfv2lp
FRd2e/eA3hJzzLkqwfEv+XCYi+kf+A/kZEGmvi2+CKCHt4prFQnuW6bSFaeRTkRYfWUfgCI/agps
BOypEO+wu+uXaUJw/iVDteOkd4c8FYDiHbz6euaBKe8rwEkUumiX6DBWPPbwCs1Wmely2fLnU7b+
O7cR/RjP273Fvf1/bw7iFpjyBLaRIwGJQ0O4LxTU6X91JbgraqFHdriRW9Qf/t0NnvTKLDRjYu95
1X5Mda5AvSB/JGgUwxxpyHgTL42cBwsWcsoUZ3AJesiBhIvocU32MTx+Zv8ld5o7TOL183GS67M7
OWcnr9/l+20fTTRnIn6VFsGgMc1b5zTXNkK9Z0j5jnwFrzpinf71Os0CBF6rz4ACUE/OoT0Pb/T3
RhfWF5TUCZAgWAKonadXW6SC+bhcJeKFX4DvTeCrUAvMpbwoAYtPli4yC2+mg0WV7ildljrk9myQ
SrOS6EcSh4f1FOpIwh7iMNIVlPylF/1+AjkxEGempcIK9fF9qdujqBT3Yc1wjLsBvaGWBejHpSCe
c9nZkZ0lBRQWjEzkIVZ7E/JrSz9er2HNjb8nYfgmMW/5QSknn/H2sl6ZaeiFlWwpgHvV/d2ppre4
CDBb3b8m6tgE2/8+Ur77mpr10ZCD50ovNj2xC6k4m5/HjAVwz4zHGIyWdguD1Yjy8ONmDyDDZuP0
eh6dWclrEAa3qQoH63O4YFcB7SW2113gb/LcMzuKxeKIlQ596XK7vLDO7IXFwXNSQyDNc/uM2D3p
r/iA4cIOABpsloAYd1rw2h94IKqPwptZEFTE0ajoZ3ik5mq2R7k0MTAhaLtSs7lfLijf9Tw3+3gt
IPkQGgJKNB8v/W6GJb3wuQ6HkM9mKgEu949jAuMxRsOq2EgS8u51D/2toC1K3rDCCd+FAG7msUyC
A99msxu/m//XGBX28XF4OL3WtQ5nI3c11gQBO6dGD62PmvXEyUY+T6DgIr5MovjAGVs+zSenyJFE
0vJ85z11KRapfUwVdF4VjOGwG+yS0PweMRok2BQV/27LU5+oi8tvvO64efIIjHTi1sNxis9Jg5cS
uGOFjTRTCcP/7tFWgNXMLz/2H0kfGcUbM6rUucCGGHy/CQ80F3zorlau/9oaODoAggu9VElq9aRS
CA3OispduLoskM8OdINUyD6jxaV4PiZWg7T6bbbmC4LM5eTunMvVjsMxrG9MbXNbmrTpnWZTu5dn
zIPA1f04cElVZoja4yfOgkQXgDpW6SgXbtYRIfXMLdYA0X4Be8FjmVoxuQYM04zEPlBJOlPfkfQ1
Tp+5O7b4CRD0WipfkQwshr7ObJEWTOZt1THXyw2YjpbHXX9x7Eck4B2k5iQxQluAED8QRMHndB1/
gGpndbjCWoQyWyzOVLXK13C4y/AGog20tdYfcQhW2VYCT+w0B87Ff8PipaLuKujmx9TdmsNM2PKH
BQAON50FI7GPlXaYSE94S4aUb4htXtyTdRVJLAOpaD65+I62m8A4pBYUjMojOOblsbQIusHJXKRX
yo/Kc/eucLHzbzKnNn4TGAdOSEcrJm9Pcs8gfVjXvCVpJrSdfqSlCXhxtjhNe/ZWiY9szS/wfc35
CurQzUdZSq0tdHkVu+7U1fPXflyd9QWq7N7rqpWKYW6pQFw38tg4gE0zUy/HStArNVCVRHtArIqA
xkYN0Zt4DdVU4+3ib8YWLdJ4PPpYFhtlTBbsURviWW6alBJ+/EQCBVCFEKXWo4iCLGtuCumC2OLP
OSh8iww2ErbTxNRiJcSrrCoiwdQtMXdrLQvEhYNw8VtD9w0S89BVwu6yrojbrSCeQqSNGPl+ONCy
4HP56CCJIwcmqLkM5vNSMdzo+VdYododCLvB+mUX8qhZuK93J7RR+CIr5XrDcPlqqnkZTvi7eD62
//RondCVVsgYBLwgJP9gfy1AWfg8uX9Lj2CZRERCVIING/PXSESzD7UyJQ2C7a+9hrtpzSzS12Om
41xTwowFSZJZotlmK/gObWFAiWGfdPocDBoBfRiKJ6Sa/hqoBNVH983jb+/YB2YsH0RO9ScxBNVe
N6BsqLRajfp08vhfNmauaMBqRK1APhijStNrwz8/wRHAXTaCeOe2h0d7Jfs5+YWVmLf/rf+pTg4V
0ON45Cg/T4dupGb0kixPCoEld3WAYSdH3XXMxLOPcdJIsBPSSIkjkh2NWwUrpSzPh2bQTfU/wc7a
wwYievwGd4+muOuAMD/CqYQ4DIJyicd/yGxs7rDXVTCCSTv5vxVKk46ZZcg/cPrnUITYGCaa4GfW
wLKNAQ9r9xm0wsMRho3Mme5J+qwsZmsQDv1zirzyh+QrUSV46K/zqtYF8Et3JAkKYIWCuFcqZ1Yi
idWzbPLjHrfcLvane3GJWYSe+XcTU98hOySlvCNQf1ydV4W7YLxtPLIXBLPir/d3UQybuaDVUVki
6EOn27tEk7bb6WC+LcW+7i2/Bv8pNAGgTaPWLbCHHTAqucS4rMsAV0PwNAYKoCFNjsFCR+lker1I
4j6HHW9UKAqegmN1fM9uyiceun6iGUhmnmA8RdtmQebnGCEVyaT38Ke9rL0uNxzYSrg+KPYTZJbI
ZLtFFOX1fpCuZivoUz0i2HWPWLnQxjFbkjOZoYQjV6/WNoKWsGFqwkXYZ55sk6qxlCMQ2TyywGTS
ecQ375WAnxnzbfIu3eMQz6IkX6ZVSAivOKIu8So70rf+fMJezX6R8oz/NgoWQC5E7ELG38ezVaCo
gGdYsCSQmt0S30txNbzgh7lsrPjwJIOtvIHYd4BPpcqCM6EbQo+6d4POFss/emWUxm+gFnAn+Y39
KyQ9oRTWZip2F/PK/Fg9xy1dEJpE3cWy5fMZJANqPoXX9mr/JT6u01EsQF9om9AuUkbmgYkIkgBy
/N0Xg+lbIVoIdzE3AJH0AhdUplGmp/e9MMrpb6LGQnHAWYbXjKwq3Jh0SGAZ81L4sqODG4lNLKwp
iYQD4eN9Ia7zxNy6VbaCiOhimRhngE3Pmv+r1+vNrAFHASHQoMF+wBqhAfNLI4FOiKN8yQaJKDRJ
/0UgDAmUw48OIZyLdZ5ZbRvZGG4cFuQHh9Chm0sEiZHG90Aep0vnPBJlgZJVA0/HoeLe0pv/aPoU
P9po8ud9XlrB44co5bX/AP2M5x+5DIH/DiGX81bZnGmwVxZJC0MrKrTDEdvwXNZ8QPdHtCIrSlUT
2ZLdxeBkMaEaKVfyjpY0pveoy5WXdElgvIzKRmj0U9nSWKc8/yBJX0Abg7NpaOFH1lmKRudfYmg+
odJpOEAJzeDeCjVfS/i+z3JwKWkQrmpOeASS1unY5rSR37CwM4xUlwoYaixWek/gm1J0912uXVk2
BPVeser649gMtG51oS3DoUZnpZK8QdS7StrxaY7ExZcf5QQvT+441mVkWbBClCBY4fUKpwq7MDpP
9DLkEPZMkUd3xMEf2cUKu9PsRAkZoYa+DC2vi+tOPfl49gJe/1vyNO18+5KLxZoVQlrED9UvDIyG
YO1whrQG7tX+yMWUdUIZI0XtsR6GaM48mGrdOubpN4gYr3r6VmeClxhdrQ7vwXPekSIycaXK5IAx
ojP/yLvJ5Awbs1gNPNDm6de/J5GSvHkzpy0shygHWR8Vz6fXxPd8Or/DFcPcNxQhD3T1xzapXHdz
6PEs7OQ3TKxf2dBZbMFLAldJiRainvVgELM0fBAfKxDo1E/HFTLolRrDk5f4Ru2CwcPsmDiH9Aid
K86syKXSdbpv6jnJITlPVAZkJoER/4n4XEyah+H3zU/XELUvmSBL78HY5d7/IjRUmlHC3UbwNmpJ
3g9UCFh4L5E2DKSWdJ+u361vSxx6dLKQ4qyYsbHdtbCE4QMtrdMrJbyzzcS8vc246Yb7me56osEh
kpgr7S1V22jCWvmurnNh3I+ousOwFG0JPediBju5+4SSkSeTm+P+v7NB05UKdBN22babNuDdaAS1
JVwZEkNmnuRPz6wiyla6sy74LsdfQFs8WZvRkQ+fiWbXzkjS9xKWdKlHO9xJerUiEOB7c0bn8RsO
2tr7XEWnPrh15rB0uLTfuYw+d8R8167QMPRVzOZY27YJzzVZUoUTYBl3ytrgwwQN6t++k2ZS3w2D
ebEkJMK6797NSmzy3K77YHbl5cugy19MduQGvlluCc2W1dqydORNg8etJlJU95d8t4Rdjq9/sLq0
i67MuVrktBxfDjAlWwI+k7xw75lWCSuw985GKVqtuECvpaWymVEUxDjFUT85Uq32I9s8615j7a79
FPlh0BHbEUGRX6pgxyDs5Gh3KhMQy9AqBqGtldeLoCm7B5pi71z9f/aOcmGu1df7RFolBr1ihiFY
olvHsyXS1lOBi/mi+qsudvfkIyscIhkZ37rQ2xIMEu9c9QdZsh/ZV1X68YFJaDWteJeFpJs8pwzd
6w9fWnhF0MNMtCTHRzkQhORQvEe5/CbJFAhJt/7jsvU8X1Oxcjg9iUDyqwKiRaVE9jItr4gQiQ3z
ybz9BnpC5De3bLpYURbcPj53mr0phMGIgMs4D9ncxUqUP+U5KIy2cpFENaKxxSg3GUCHfXMTS9cr
nRdMoV2Ytq3ZaLbzSaou68eHG5D0d4R8fDyKwo+nBVxPx7K67PGPIqXwgKt7iRTb9ClME4tuZyoz
p2HLJDCmnCUA8lD8GC2irZQ19ppA/RjJKA5HQZHlGLQyiqcp+O7p5P9DCWyhyRg38StfBtMf160k
k/a0HG8GK7VmXZJHFEpD8xip2f83p+eGkN0gite2VQlGPYMd+twLyLnotAV9P/7cdyDkySLWQ6Dc
XnJjdAja68lXrT3rGdJfZ6ck0Xb0JnjChFdxeksCBp4EPQZJWC6rvfMO8DD24nrfX0m0kNg+l7lM
k7dgWQtCE9qgJESPunEqNpfc489HICpsap7nHMqmdQci+Anxlp4SKYGu93awjsKNDLPiID7kth6u
KiZuWr4gg2LxB39BAjodWACa39Yrqvq3Zs5L8jKOEk2ebFdJiHX2nB79sQct+Fd2hkxGVR6ahaPi
NqiF9TRlB1sJ1WnxPcyUQll0AnNvkcaCXTlyVRdsVcQLukTIbXF6ICZaGVjfcPUq+kthMGqmNlmz
g+TP+1r+2/Pg+aos05B3EtgxIQGDNVG3EKi51WdGkkOOfuS1oZJfIZXmsSw7PdmKJ9Pn4qbdZzPO
eMvaBB2lymO9bpHtq2BTP7NTWHKxY7pfK1g0BOVuJkNvuzlEVAX6wc3N9KHg8CCZqJTrJhakyq71
b1fn3xNhzJryWyeKDhFp3uNbA74SVY+E7XgbqsAhivQ9dscmIy95p5aoEdhAlT87Zwk1SrCBkMuL
LYHEQYC+lpIvQsIuvdkseVf2oauXgAMAnLqXkwJzcgYyRUHNcm/A0nET6VmQpWnl/VnB3m5ABMZb
5kA+q/r185YdHr3EpZCQGGkQyEmcEvcT/oJBo0cfcBqVbC2AIrWIjlVvQHRSeLZTGeZF4KPdZAM1
kYhUv4cuKzeiETAWMBWeBYQlw4KI1BEuAAGDXmIYKCDvdDQlCQa/FGvWx7Ej0z+xOYV8A4jetbxQ
aQzaxm0YGdYce8STOZLK4x6LwIv7fweaIf9+va3ViN0rfeqTBPr4Ry+KA8xNQJrEhr5GBkKSa93A
RGkH12ijePJHy48+6gxTgjn1gwhJJ1bD45rZGCxhtwPp5je2ltN1h/iTPGibRn1Eb/250agmbfaM
QXr4jZO+YieBt2Vom42SaI8xAGJKDs9bMIsLsE6iNitSm9bVh8fltl1NWT2pkxoGUZuhd38ohaQW
KNrtINzSeLPNNJYOWUnzO/VUgJgR4p8y+NfpiPO2ba15xP4SYaXFERI5ZgVtSVJmFTw36+5KAomi
uyRFuvhufhOIINZh19ncg5AT4ofvfzWaP26HV8I+sJsDgT+wjAWxh/dukH4taK2HzLrTGzqy1h0t
cDQZHuB+/tximd1NirrfBPuLc/VG8fHWmtX9F9yT/u4DXx3kkzug8MueEUYduHZbSRh2WaOW1f8/
qmII/kZwjWLESfqp9swjCSpeYUaGgOgGwrs/9REgNDS3WF9eahG9w3ICngWLvdzOObOTEz/H9W0m
PL1yw+HFekpgXgVE6pgjFHrd145Qgn7su2VDAGxI5fkhuefSyYihIsqbXsN54V+uvkZ/snk3zbBb
aq3R0oy/A2fAbM51IE3M+dPGJLxT2gqhLaND41+sYd4df0Czfmggv4m3zuS+U6VAy76mPJNedXkU
C5eLCvHYV/lN3k9XX49vRdqsMjBM0Ou59/mNFGoi1TlBAJcJyhiPvujAme4mHMWN0Wa4ZhXxfCiL
dmAfLtUigqYUNE9vlR7o2JWLwuL3O8vV3QCNcOio+2znADav3XqPXsbGck2lRYVLtyjEYk0HC1HU
ln2s8Fr8ycmtDgAmrSybAEcfl8BqSqEUf8xcAIhh7iviJw2QbTblLZtWP9M68008Pfrt90b8eKha
daab0MMOPcDNhOtFRxkylDrQcRarsPrTLAUMGQBgUD3ZFjnTu5El+aruJM6vucDtGcnRM/pjkoTD
5MCGM7QhBULGP2S3fmiAdXunz7oHnHUkhM3OHdMb3hmcWaWuXWo+CM8iRvrhiyjlAb7+PA/lIYBU
Njs3InUfBpfmu8xtZVYEvMUEPWUfvb3/+Uz4lu1hQHdNv500jZ8lOk3QkFPbiXBvM6di0I9i2SQP
twf4/8a+4Znp5JlyNy4vZqjnw0b3T6k6Zk8tUw/T0yYgqZ9T2hW4Hhvnfvz/sxYgM7ga4HiBuWkc
TtDlLCxdUaNjVhmVK1HtbfWrNvym+IBJ+nrnTd3NE4dZTA2pBzHkmQ6sOHYdkgyrt21h3jfWcpUm
BdgMXwPFuqFUpau2QqzYiZby5TwvjVqQHJIEqh3MEhYVfoV/USTNdlVl8ndIAUWmhppddAL5+pca
aUbY88Ihlp8tmueJ53LF9CY8AppJLHq3ufWtwr74VA0HG3UM001PAk4pq2jVabfOMcht4IvOGKiG
HLqUr/KdRwwr32ORuwj2Bic7DUROTuQ+dpgIxX5o3L2LfbOpWhiRhr9wA3qN6AAZYtxJY6fGDS1s
FiQTBK6ZrT4hoWEl8IwkcesyuUYvgdai5AeoOBNtCgRsL9dKUkZ6fdlQGhRKSfgDQ21cAv3GRTWH
/aJFaDINybAEwrelRiU6mwHzwSPudXt75QP+wpQ6pVXEL6Qqwr8ksJSmzDX1w+XT74LoIYgh/cBv
dESljZHAHgodTzIvWzRi1QtJuquX5LAm8VQn6ucfUWEfBJKR12QIU5ByHODvUjEb1zIMxv/gMdZe
uMRyqBtTLdXW/Uy+IdeW3Y9uuUwVjk2pPkpgzyDtWInbM6bea0ureplnEBXvpskPOl4KxrFz3iG2
88v76LozNvlHPG1xtsyNV8yhLF/X7+yW9V6Kr0hscTIQi33utAy75zRzu0XsTTWaNgvHRlhRhVeB
xAGbYffX62XYc7F1Rcr86MDLbiISybhBgjl5ZRz+j419sZ/wvzEv4IFaBfOe3hEsXy4ZaDYgxkN7
N3k2nUYtMntXArpxC9ju4ceFdxcpbzAixebRG5/+8FN4lebv0ChKcRzpYCIRmnsIJxomOCA45Q2x
5HxdQedYrejNahIY8QDsmi8DxRNwSnY/hDqsSaMmx89OVg3n/gbhswmNlrBa4u0Y0vFqEu5VV1oV
DvCdGLePzS2uS5PCkVRX+rgxVcZLa9JHRgbcjZFuJIVFcU6kiLSOJLc5zi9DBqjCsuH+bH4GpvcR
j+mDiF9wzHj2DJuCtLPb/I9rh+UiHTo3iU7byItAK4nr9ffkKKe+zHWFlWYE+MJRMUKmZSgBikvi
BhtrxEvaqE3E1if7BpWj0oidbbaQQwfIm95eQKAMislCtsvs/ZHsUxpGRFNBdX2QBU0sThyO64me
Sem1gz4HGnatSq1l0xrHHUcxW2RcbMoIiOO+9vevp/6MrWqsoSjlGP4TdTnxWXGLOqvLK4tCuQBG
0BkRTodGIOMrvnV3QZcT2MGbjIcXmT3O9C3VbSYnw3AobsI0DyPv8AkG7O0LcLDbm1JMuZgzA550
fPRYsqLygSwC0KcNdK0RGB8kNKlxrVQ2cY9w6ZKEHO2tBJ5pyVrjntEk3Ze2xn7uksQuGh4tbw5n
Rwj8ePHXfatG7PQY3QKQ7BSwgwGo/tUKwt+m2G1dm6QadyFh5sW3vSi22K3qP0W0i1UkvjO3FZzx
3uaM1OMEfI/DJSVlC/blnO3POGR927TVnkj1q3lZ3m3VaG5mu1vDUxlp51eDehtbUJusuheNqzRa
givl248kOprSWriRQGM0uVtz1GtUS3hzW2VQ/Z+F0CFX5CmcaRlbqGZHa8zvIytyKoP/xHg3iC1H
e62FxgNQs7qXYV6j60UMyC1XfJq1ViQNpdY8AU/ZOCeWok4+oilPpcQ4VECzbaNy/tafL+cVPcTZ
faY4YAR+iqcm21FNZEjPxHIY+L9kwm5yEzR1JnahABVU4L86AmZffxecEGwNj01+vk0rqm5EdzcE
16I0Mka1+fP7bwGYa9BA+IZw2P8UuPonwyeY9oeO5JnvEaaBlrPM8NAneOv4qLdqJtdbu0uGOrCf
ZuR0Q0fCSNirYfPJhFyQ/NtgxZYibrU9M+AztCINcGshJfpL9yE7rP0fbcSi6mexGOfJf3nOwAt3
EoCuUwpttuLsF680G4PxUoGy/ZFKtdVDvXqtc0uCIRE4yLzWj9YyW1egNu6cGc/+HocM8C6EOO1i
vdhvZJhdXuX30cMSUKpwqrfAlt/eGcYmmb42+C6T9LlghzbVybhuAFz+XLKxMd6ccwyTEUJtJtJM
PvZsHJswByjdWpvfFF3QxzTqJWEVzLiMBNtpFM+6iJknw2mn2GaAjJTz/XnbCl6FDpk+gK3q8Nae
FyY6IWWAaJrr4ufyfSOX0JyJ8EC/3gKelg4DJQGDBeTxlqpQmWOPlEp/2VPhJKcr/o68REsuWQcK
QjSUprbnykYyTWs5Wzr7GKQP+epg0G0dN6PZ+na0OpQ072Xeyl5RdP/kmzcMgLPsq1lx658A3N8I
jZ50rrdsTPI5iKHFh8rO3h7Xe7FIf7j2B45NVi2RwNp0vsG5a4wdj+f+4KpWK0XUxTNJGitQj0nK
eLWX+Q97KqTSdikICvHRFeco1btvVsd/fKp8kXZkw+opWuqu+E8NV8WkEwW5gYX6C0tk8rCJd4CH
SD1r9rs7jVsEG5tDlBUxrFGNyr4h22QwhWwoz398vwUzj1AQ/xDI76m25GkZjaFuQP+xBdO1Irjx
zSeZ0QY02IvdoWQ5on8SGQokqR64K+U2sUp4aGCFR5lQ9qjqUEQr8O5fHeY7mHBWDi4zvQLDxlpm
VOyOSA1Kr5MG0OxHIHmsNRPWxNdyl1pK18006ifCWF+UHnsOUJHiB6Fc83rHSV6aVoaJMYfFI6Aa
fFLlM8Mzsw2WoaIdziBWRjFjhMkBpY8PFPRqzmCMLbiRT+yT8yRd1xSD3UyPRb2NbL+dQCZQQMvR
0X1sNs2iK5JMHIPZ4cKpQ/4lJsUXDwCdb2VcfjwwfEBUjemMVwgBeLNrQ7mRmv2teBTU8JLp50da
u2ctU6HcOlnED+MN4ARGTE84ahUAVcM3tivbJOn5WS9QpTnpdptrMR4i8VvCciOdUaPjAYlOXclN
TnE62LjVoy9IGCdMbbvJlm3NONEne/yRdVE+zypGs8q+VlsMI2MAfsOFrXdS1JYuyivm24OKy7HF
K4ZCUqD/HGVKgyD3oZTC4+RJ3j/qL1ssjnkHeP1o6a96P41RiK+885LvgmNKEyHqZS4HHbxSTJf8
gSlBzOgPONRq3OihMEKLjj7TKC5eAc079J+siCJhAUezF4HF2wTuupnRJaIvMqZhT8RhOr/dS0ab
VCkpMlBgLvhg4b2Q0RFrMHMZ63a3m5v+bcuwWr9H/Fx9K80+zjW5rOUBsY4H21YqtQpEizKH1+bS
eNZPu1X/hWCneNbxdMcI6RFpB3P9t2rAWLQZwUJRGFI7rKJBNl18dc6T4iBidmkbQt8j/jBQZTSN
uNaAUOTYiz1G2DzxN8S+kCp/flN14Felu2stQFOq0BIcLb3eB8j6WZljk9015yE2WPv+5qVwET9J
zzcg2q/LlqXyz4llQZfxzZvG5uIzypxEiAqfXxRcfb/VqG+EgREjXSkp7vSyk7n7m+qGCtiO4RQN
hhjUJx0zRrrG1ijrTJe5/aOJsfNivkC63mmRC8tZzSwFvqX9Pkso2eWwkv7fqpzwfOHP9nt8DJyu
qmpweKUB0p7PLwSVD3lVdQlHBQMRauT23M89Q+nJIizXej3nThuhDAnAnbgR2Jcam0PkV6xb9/dW
UpZOhN0lA2Mb/2JV6XsbwHMxY0Oxbwg49nLlp9STrPpSXgurW/EaUH5ev3QlOZwgN7glXyxF+D0T
bTAVlMXqA6iB24WpkpV+0RwfmVYL1i64VKaMbdB3YmBYCQPP1m7hau3xFzKRMLjOESIc6fiF6hQE
PCSSvMXwGat1bCmhDfpYO7Uq549pbGUI9o6l+6X9GKqrD8Ris1vw0/GBm6YO+NlcJ0Cpkpt01E1C
aNm+FMcWx3kPa6myihCwB59Cnhdu9nCFgv4HBxAs8bJr/iM9x4Z3wrPwn5iV0yJeON+adDUOaL5U
N6vneT3OwnD7Vb/3+HnAFrdMgM01XQ09XxP4y6M8ynezNMO/RrSER3MAoUT6KreMHVM5pTf53Eln
pNafTBlyomGU+g3HtG4zPciK4NOSCl6Q7asgSh14HovloAnkT8PTR5wbHTmOogOodl0LuD6Q6o/z
vqsxrcx7DJ9A8HIamQF0OcPOIKFf6GsuAu29HHRl5qQjVGYyJypSVIFywwGxJjObFbwtGUTB6c78
oBT94l3kd9XWvO0z3giJKeIEEHOvIwD7gP9wdHzJLOpTSGlCt41dpl++W9uU3RWX1F5P4POPi+bf
PNTwItJSAZDcs2UaWRGrmc+36qk/1vzmV93Jm2Rvf3Luwmo5rdH8ov7tfAhzUQsO8ToC2yHTdlQv
44DVGd9xC6D9x7pVAIq//chsqYV11gm/AypeaqWg40pAs8x5Gcykc8jWzHXY6Y34DLRamZyskPER
yI82W2fR4o3bf2VY+XaT5lmftbMOIM6ExluBCF2yb9/qw5bdMib9nhm1E3PU1MrZoyvvGW2EJu6z
CqWBPsNCgaW8JduBsyWQvgKTNJr2w1DLoWZRnrQB52BSW0Z79keZrxp5Jjw4P2rNy1vhSRjdlmkP
XWagrokvJV+2P4xFByaBNsNc7sP8r5ecgEvtGMLsrNZ8VCPqgp6V6ME3G2p1CRzyImG8IPPzuqi5
e/RUHNwqy1OWBbhec+KG9slTXnf0OTFf8DoRPMjw/PEA8KXI5KYXPtOV9AIFinA8hk0iMxB7djyI
EUfwY8nTSevnLgjBb+RZGJq+HfqeICCLBOvx1GybwqmtJGqY1Wb8uyqOz3Urzm+RTk2LmXRKUXR1
ioYCxyaPiQGYk/JaIdJoJejdzyuzAXjaWZePqD8cW0Tt4PkSKU3d4ocJ1gy+h28bfxSmDUXliK4O
Ds9aZ605p7JaSRDns3Xfnoot5R0+tZBuqVGCNKsAziwLF7bfZRy6qAQBj3esihq4bN4BXO+rEQO5
9v0rjR1WU3KvnSFxlzSQR4FQvIfVhNAs/mjXi9F9f73SEijJ5j2jgQT0/wsAuznq5golRsy4+2aJ
tZA5VhgcvXysZUUFvHr85XICKczTBl+z++9hnXPJ7wclAPMMTbdLLtoJMGunlF1jQJuZ2LmBYcSw
g/hPgHhZHjxvDySQtsL/MTpHyisaHrWSukd+hbZTuZXVKnp6UPNeRIehkH8rCutk+LeresgzUpla
8ItLs/IktSHTJKKd57P9B/Lc9OwDcwewyAVKfyMkrrb6cMG7VrPKbWaiiJztG+bGAKJ3fcsTGxrk
tLux45nsYNvUVejbttIQf2XktRROvefN7VJg30mzMpXdkLewa38S+D2mHRnrYBL28NEKi/a5ii6D
lNI9eS5/HtGVnFlVTPoWGay8rZePJ8Q9vTMrYbGpQJ7wW3fxbBiN4Si0VTu3W8hIOoQ8zFmiV9MI
gXSyPCw7f63mWknsPdF9OupcJbFBNcbiZjFoFzNiP98b8OZv+IVcHVO2dqUh7+ttLkj+imv3jCq/
ui9/4KbavoNesyu4/32SIOafXV0qkHR5M/KMKSnNkrblvR0+U0HQsH5HhvYOgTSFg1pZ7ZWQbJL4
9CL8SvHawG/PZmQt+OX6mV5v414cwmlTmtwMEe0lic03Yr2n7cH+wp25uGil7wwkkLESNYyamozH
+OOvPfxNmNlR5hdMqLSMa38P6EBc80WSoguaNQClOWkvehYpt0sl8aOebxN3WbEa2BrcBt6nD83Q
xl17hhcULqwNt1EgvteAOsOiXSka0PdIFKIAQSOiKkqU8ZlZmvTzRYyxk231EaVjyIxoLS3pQULF
vU8kn5fp9f8GBJ11SrqMiLJyXWD6NnwTzZaOzozugw0Ol0lD8X6pTAoE0bZ7cjJt6Q+NmS+G8nwm
cdkN9MwIAlvHdQlQ36RQtNwhEhWYeqJAs377AaWTNMt2yjbiG8Gs+VBvms87R6cUyhZuzA6bTsuT
YumKpnc8pemgCTUZ4ds6fLsn/+r2onUhX+uJUHwNMcR3IMU8REDCJGhEMow6UzorXYWyw6gNHJYm
H0RKiuz9Qsj7n3nd74SU5ZOiv5dFGc6unWa1KR8gMzEpIfub7PwGX9RAp7AqTzuLXn5ztuOCvd7t
YacsiuuCh38UjMeXfvMJHq/gd6LPd0SJJvnfOd6rjFzJ9PwOrFUgKrI0WY8V6zEkilWgPXKZCt4R
J+8OHNayFf6B7f0LwN8nGg7JS1n7hQsBZn6bbtiLhXyJy4G96sQcU06x7w9npfqWr7HnBN4dn3kZ
Z9/VDT22iDqCEDk/3IHkdtwumrVvGJHbIcyBBgSba3UzrXq1THIyZz3c4O7B/mk+RQRpXbRalpOy
Xy1WpbY2Kgvvjpy5Y4H+5KW9c+V+5htmu2xqCvSiCnKPuElgg4vaxLDQKFb5y2DnasMkX2uRSbX+
YnhA3WKVDxPSv41lt1GcmdSVtyo+juLf6fxHs9hMBsaPQTHDDiZmc0QofJrMNc6Ccfg9S+WHQIDl
DrXoVHt2eDg0aV79ZL4dA0lYZWTLkOqHMu76WcBNB4FI4gAu7nti6UXO5cY2GDJdZtXp3uWZIgB8
is1rigHe0BnBC9bL81bSb7Cw3n9j/hAMo3x7ghOpu1Cp92YjxcH8lMFFopq2riR7plEJ0MZz0Mc3
Snlz+UtcRUzLl0b4Zr6RpUVbwurwAne+FBfwaemGN+oDhzOAXOTxlrL7Q4+Q1EBEIKt5TrBiWe1n
phI+lQoO97Pk0/5EorfZcHI3GW70H4d5gSIfhjhKLQyxFCbnkhxoJakaIH/GLJoWvJR3wcKRuzsI
P3mD6TvMI1GBBmo4ZcaH0Yr2GE/8ZKWsmOb1OQ4stteN4g7Qi/BdvQ8vhMrxwM9vWQ3Vu994mzhz
xPUot9JwwHuN9yiwSOissCaSIPf4QEdVQSOUGfrM9sPynqyUjGdOHZ0ZfI+WsWxDmDK/ACRVpTw7
QKUK1wgQLgvHbhoKjM6yTSPqDlkH6ele156ghXEsJXNhvt7JmzSmbzZyVdFJf1K2M0ITgzMb6UZN
eFm83Y95vN1xJRHBQirjZde1RhOzq8HBAwKjxr8vQEXbgvWQuHkUf3Teo2NefHF75roquRUcwSgR
wu9zuKWiqQP/BoScjHeWJK+DI+F1aemC0jygOSM9MPlSFUGp+CWQ39woW6sjaAsWJFg+61b0IS7b
SHTpYTRmaqm7YqB2qQ1JwxihHNx/VAfoqdlfS6lDLgIRmQJ5JQiGAWISCvr+cAaY95XBOi+znuON
/+jPHPJYwOWhREYL+7S791CQ5KviXes1gWs5EjK22YCi8tvzEoYpmSePrd8adM44nBjLaYPYFWm7
saGjAnaFFPZUg6j2w4zvVIeoubXEKjBfilXWElEUL9If6LIDcHIOIYhjBvwMS3hypAix27M6W2FZ
5DYH1kS3PZ1u5ysflxFeiqpWSt5O6Fzw4WWaRKQL4r8ES0T9Py0/YmxivcNNsVVCVjEogRdYX88/
Y8kyscsALnTojmYBK3hRk5YN94DZ31NyTlRQEg+ckVtYGtWGhmlmO7wgix3Qe+7EAZtv8Tman7t9
v5S4Atp+keZ3F9tDzOd7tOOzZFn9S8pPOf9r/D5XNXh6GsJzwSCq8D5HilBCmIxPO7rrL/mLfsK7
K+KdJkSwl9o7IwKuBjtOTV1GAIs8rqGqA7jth7oecPGIhG8hQzlg6rzXaATO1iCsyF4Ht4EbSCem
5L8H4ZztRvyZItio+VcVjX/CsErFGJUP5ZuJ7Jb04hScNk8NIa3TjStZe+bK7aOJ+hmf01cG78oV
6YLSGZZwgIR5sKMGC92K53UN7xuSha52LN1W52Fu6a3uLMvogmEKWxbl2WtRNGqCLGK2AE88ZPC6
loXD8bMrNZeIH0jL+wafgV3cTAuQPpWDSLp2t/GvZkudxPNY4HjfPgptHYvw4VjhgY4PfY9gAhGS
yxzjJeanKiKIphHLOVq1TI/2IBTSaqIoPnbtz2uYKUF6fz7gGfqsz7FBO6HFfTICxxXphBy2kuMq
bNsJl5829DYeJeg1iQAPP8x1PVh3NtdhEpa/Ye/kQ4P6/fqQMUHxm8d0TqEgozHgoRTIrjNLO5Wj
IPlC1eRzAczixoL/jxImjXfumef8viDHjRWjJvVh7lIWijngE+CuET8pEiUJGfmmDz8P/DfEbNr0
/s9DMH6SB6oi/rbxAnZqHa5vhyt2/HPv1PFsWs7qpqIZyhjq7gDXpkNwiSZZV5FKUajOM/7LZIsG
XXbooImAkQkEFfmzy/3LvMZ5j26aMTUg/bB1m+jKQxBBE9AeoE+L/xTWudElXSSEWiLwnPhsUt4V
RmGzTWHkMuvGj80gpraGZ6YUxvwOCP7xJVTKmWtIabF2D5wUtlZ+30xnCI0MR+mU5JE2/sBasUPG
SwzLZ/2nmhRRdzOEzK7VqNkrWiFqwfqW62hNu6n+C1uOIJnI8lL3Ui7Y9v7a/ipO2zl503v9vttp
M85i9wAHWvJNEWVClKuAELfDAs0J6EXa/5tC3YdB2M8ryME3I0kI0BXIAP2mpyMiRGdvNDYKEvTm
gJO6siW48UU+C2f6MW2nx2X167kaVLNcDCICn9I+YYFf2d0COeaktDAAdscZVi5j16Sj3WHFicII
nZwvxu1NEeL/uoRYgDfcP9qA4rqfD3E8yjeB4UGSjgzV8x/5p2XA9uzOzYfMkkSPDrGBUFi9ABcq
/aADqE5FFmrUx1wFCXytOqnSQsaYAvwKo8cecof2TTNFM727Xudr/XtpUfk2RH4bMZWNmV9Tzdjs
qKOdAEwwLp4ATbu8ij+8WyEMpGGsUiUVce+n+ZeeixJ1dGNEQyocnK98gRFy/UqFbrI2xYehXOoY
mfsPHA2+Tths40LYssJsHYI0KB/X8SQFrRw2UCntLexxPbkEkcSypeZ7R6TeAch+m+BNzRhMCYT2
nSetzTJp2GVFXn0RMt7HzArdM88Ff9W59Ff15no7LiYAc8DSMgSUn/EjWi/wcICKgvOx4K2gIH+N
hRxwf0V9O6Ne4MkJNSWiR/Bn22B1KaDPjYUKeplaNcPQxJjxjyDZSPXA5G0zBEBlZauvLMZNQR3B
qa0G4yf4PSW4lhEe/aQhOLUtf0q5ZMTpjtiRgJ06g8sA9SZylkxN22Nj2BqpltIbUCXPPvu9QzAG
n8GVvLhgqoTBKfeL2sjVKR8hSw32y5WInXMv3LarICw5kJr5/1TCcr8UMT85JxdhZsyR/609ynuZ
F8KAk4hsPPIpcuJ396HoKpiSfiXLj/XjBIHqS9k3mujWs2CoeNo2U2WJGPID2TV6XXu9zDTj5ziN
D0xFW4JYGwwJJPO5xo386Lo4I5NSUjdoizGP2j3QAML0+a1cYv8YRREAR5elcBc8SQbBctTgQTqd
YJlkpm3YOoDiT3Z06ow7/wECCatDrYOQ+TY5BbJQpZYxqVUnjCd9QVFbUtw7N2aBHVJb0KUOXJI0
BavdYvuCMvjARGPDnqeJw5sHbibWv/47aEvpa+6TRZvDq5Rj0jFq5qfbYZYO4SNIvfEZPkrcouzm
WYQiqxpR91D4ao7+We3N5B1O+F0itE5/PM2C5+TNFN7N9xPgz4PX+wUiO/8Cs/T+N64HoqWE3/Qa
+e2890YmGpFxT9xqU8f0ER1/xBM7ZdqfQt2WWLdLrp7YCj+mXYUDNpITBrfFSXj0wBJ+a93O4vKz
NRjE3oNJmDqJevFTPaP6dgNYBRKCy759G3RN4Yl5dNg7m/VMjU1ha7AE5bBIK2x+PhuwpmLgc2zX
HhrBN+izkpB5iBFfKTx1nTKvDuso0aaPrpq7wVJFp3JwAlEKK+G5RjmtTjfWRaWAp5sbEaDlvf+R
eZhAIMiEnbDLYkgJ7BXtMMn4hV78jqr7hljpIQtP7petN66p9nN7xw/R+NlXMqyLSwyERGPN0Gkl
RQ+r9M5j0v9tW/IQiT2M9f+tbOiv52wYndlOLr6ssGpJNKXWWHAYcg/oPUi66TCf04G/PU0npTgS
Rd5Dro/YAgSeu6kcaVzZqwtxq4X0s/5Z+b1VCtWSjr/LT3f/S1UcPMOVSGlHLTHhTWkjSP+1Sv0V
GRQ6ZZqAjW2Fo/8QSYtQ3SoTZkVZSqDTR2tCz9Q7ptCPo7YMPhFY47SnfxprYe2ngfjroB68b4PC
ZvEqqO81UCz0tdU2qtG6mSYiiuSMEfSDZPTYmL8ophzbprbdO71tTT4gq25Hd4LG4YPL0ASo3R2S
TwzEuN8OgdD1oYjyJ8lHR58C8Cmex8qY9defNbK5zSbJRfSRQJZx80tfWVsj+Ml3pCXkwWgUeMhK
AXg+lh/w/je00MgeiWFaOyTr7oIH1rIwOuU1ewcvq91I7JIrwxROhAv7X0Pmr4yLacwkflksLXuR
tGtau8arOFhOclBEeDnS80s1etaPdDkqUAM4NpKr9RruusYfUeNn8CWKf6cUyk/BW4hpeKhrp5rs
h2J7eou2m39MKkqxLk0JWZNAEPjuYCW52hllaFaMm4TaPkJqulEvre1tPhvxLI1qMLpyYl67LG30
Ou7Z0q0SKFbAiJ3a/19UeJn8Wl0iN3LAC5qu3UeqLpKMFUGh+oyK/QlPfOjbFVH/DW5jD1C1U17w
SlNbjLCRW+B1WqqiPniE918K6xU+33L0TfgH3tJwjkh63INO7yxE4MsnjPi2syne2hs1p0zaqzOx
YJfNRrVsgAIYh4I/m5J96CSdM7qnKE9GlUnSf9uEgynGVVqj4NNST1Tia+ONCiOXP1CmyekmFMBi
Gn2NEguNX4MDRUGGuG0T/FgKpXhdoLbtcTzR57FGmpmoWOJx1JZlyU054XlFYQZoa/+l46hKNTej
Y02ysxFsKMdZC3f4nGZjChVmIPx5z5JtCiuaVFrSyT7St2Q+1q3fosPt0I8EVC95hdxl1r6YFkYg
Eoon5rfDvvWekdPpVsM5G5gTRT+xtviysYPEHySEQzJZ7FB/YdEuQ/Yxk5dtct0N/+oibvd61CKB
33zWhXjy9HyhyAvPmw9Hn0vC/AVFhJIjp6JLqIudHASYwGvvqUjHp7aYFlCMRbTs4HsMol9WhdmA
9ZdtAXcmM62aINHMkaFmExplfCENNVZJqoZaWAYYFAMIU453JP+SbxxrmTjAK3DnYMhOjgT3NkxQ
r4zGWwkuAv5O8qRhHyQJRlnHRKPoy/4NvnELRiauzUDvHIKsqkJMnd5K+f24QaXk08wETK/Xdkl2
1UGcHwRwOCoT/JlEqMINEqNDvz+TnfHuwFr2+fTJYrYtLeFyQPKdAWll9pnTaLrwqTXRaJ9Dblzw
R0TN9Qu2o+xU6JLpk5s4QO623qrhH1SpwpcmIBSMqMeBZrh18K5buIeEV5E1PvXz2Vyrnn1yzd36
JMK3+BlgiL/cq6GAMIrAUWFHi6ZmhG7XJDO0UpOV/R3ks5+xFRU7waS/kf0uohB7NL/0gd7B/uOF
GYVt3uFttSJ2m+BglTPtr0OpkSnh2uXKFi+uHM3S8jLjMYTQcZPfb3o3UhSSBO3PifXyJiL70OdJ
zV1eKZjB7x9icQsSRs2tuvntwZykr/TL2uBqD0D9Tqn57GEIjUlTUSJBUIOijFMNEmiYBxv+S5Sb
XCaFoucouYc5Kr6mx17Ll/vMHSkSWqoe7Z7LPqMjVCQyiG8FoUEc9qRMUe2kQx7gbD8I/c+EC7vk
oKVhTviWQ0GjhFf4UaDmGMETMguW4trz+1i33Kq2uhzP08H7BmpL3G4LJRE16Qrfe7cNDdFV0j5l
N1luDBWDNCvurImlQYCnN/hb4gAS5AoqoOvw6v5WQwR7XB9YsZ0yKcllBPgCdHqS0bzHk5PMcm0Y
Vv1lUFqf5EUVEluttkEgK5szYXpEXR2+H4FTz8GfVgCkXnqiDJy0jCFXVuowY3j68lckf2TkaC76
tLJaQyXWCKo9mWX8o9oEzFJxUDjQ0+myXFoQ+u1HVtBgKY658+s/HFdx5zb0ixepVTBSjvdnIt4n
lke/I5NFNmi/j0+TXYyUhGtdSQQWP9kzhyajukoQ1Ybm5BTGPUpgL/4YeyAx7UYysQrfeHbgjei8
EfuNhljtlxWLTjPG7Xt3YyZXqgPW38S+XAO1zYu7knlMcs4hE4JdXM+wzG46e8srfF1OH1OZunoM
f0Oc/IFAIo2Gg0FxP93486Ev9Qj8y3gmbHe+wDdtRH7RuNCmlsNUer9p/n67ta6Dt1n+UKXqnBVr
TX5ANeZ1M72vHdf/AdWBPPL0OEStTeYKQtdsT2LVgj6dPpUJ0+Bf83rCzBvDbL66P4sN9QRPq6eH
xdSts9xR2u+L4bL36oBXIRHj5zL2cUOCuMMHPtfzk49ktn3yGcFV5QzDHPyGkbbeyISf3To9Obgb
O2Qou6+Gwlw8I/k6f4KcTw77r4MZkUaU7Wra2EDoVE6IJI9hmVtybinONL+st0QSHwUJCcaFK5BL
srhJnh+oLnRFFVva2wnqjKm3pPjcsvON0/I+RkYJXtWAtvgRuIgVJ3fQKJlPZlErgOtMr0vBoTAS
pHZXDLN/8+T7ZLT8k7G3TGmz84PXU1iaY9hIKZMoTWVP7AbMJq9FgiO76hBv8piLZPV2xIy+6cEW
fpGySg/D9q0v1+qY/zd1bCsRGGDXEay9hxpwB+pbdKE0EqePbqCyjqGKFTc5pEN/jkqAstfMga0s
3sciMHnk0nXMcgRt3uvxczDz+ZGy1HdRrWP5W2mIpLLCu81S39jB976ky6U0xOQVcwodpB3OlTux
d+/KSo7yLapgBmqe4robLTjyXxpaOqrUek3sx0LfkM8IQuMt+HlJWE8JMgNS1/vMl+HY0n4uds+6
I1069KMniSM9GTQ68wQm3QtbPAwXU43DcfLs4bwXxtZn+vXec/6YG4irkRpNRMDSap8cSyouvpBT
CDLaXKT2+S5lgORfsKTrQqkSagkWrDcbymRYa+pKhfdUOB5BS0BxKhmoRNo9nMyycdMtuvxdJwOb
7aKDjeLCwfzeX8vFFKSR3f+XiySobPVKFdfUIIsP5gTvpYk3j6scsuU3HpidZYYoDc5NJfWPRyBm
quqY2WkFBimkQ1omf5hCKB2D+G28RGCiJTv+TDdy/8GeRZCmSdjWqyIKKOtvWezZQnpYLcrpxwIg
MgrOa9smlJw6DkQ6dgDpMMkWwdxb+gPdZzgtFulpwmFPCAzOkyEdkjv2cQbqZg1BDZhLYehojsn4
XbZm6ybLtRBPSdSWv4vIaP9hd2hFPLXPh102cVFk+FpwqBqsahUg+GZp0ePySdeCC1FTSDB+5Kxk
V3zQnQ54pwzxLNuOlPkxQvwxrYLSYJuJpAcwZwrwcw4HeGrsNiVbaiuHS3XE24HKbE/KZ297+PZB
aP+8VaiMXI7YGChqFYYBaC/F/4LsdyJKZRoiJ3lV/fzgkBJC0lsGBM5qyagvcE9tTt1hUKQ8/0Ii
LsRXe4/cM40cTjBw9VP6Lq5LY9YZsV7iIKMwcdAcYRqzTU27gM+SNCNCREMM6l17xn26Ro1f3rxV
XHY7S2hHyxBQJHnqvWDNwHSZuxuqO4HWNG+OhtHT3W7GIKWXQzh0wyeqxfALnnGY4x8aXp261c5M
9Fzor+R3uw9SRYFFSLXzPqxOl/hf8mCXBfNAAma1DXiXL5Cx2in6rejKYMQ+EIdXZRknBRKUZnPW
mfE5mSyFozvjWcXaAoxYqhV5hGqSwt8pZoWL9bNOakd/wOBj/tBN4ERv3+njyiVlGS2D8MkZKmMy
fS0PorYZeGUFKLln0IsGy85PIgfvp6Vnr8cCZ6ixonr0B9vXwvXlrS159oHBefAtaLdOft+OBkyO
Ya2GSItXLNjy5GQ9xcefFsdMf1As7EHO2vkvECY1A9V/3k+6wg6bfI338U3W2VBnNz4rY/uzApaY
AqvhcTu3Q519Zdv7NICFPkg5D8wKmBeuyGGLLIMH7M3hHx8EWBKfcFo8T0l7ZC9xFoSWofUmLDjp
ipMh4x1tUIFRx/2QAZhuzXJ3mraWxL5KYBVDAHqXknCruOpZqnG2KFGSclM7PaQHFmhdr2t8JSKg
1BEzf8sDCH6gWkEtgqgp7QSdg4HjTPB3neN5ThbqOlDLdVnG1ZKekiAwLkEpEIZXEehJULnVdHqW
r78Nb1LMX1FKGmBm0HW1CMSHCcB/V61kdIWB7kBiGh3k/mdgpJraeVUmtfBdPvVxklx/RPz7vAf5
fs6gSPuzBgksCnlpWe4BxU+n1BOM/Iwy9k0buMlrnIOO3hL1H7/7O3Q8i1pmzPevzTzf2aGvEbhq
gyb2CWRUL4CWswvuE4Luwrb6RxFg3hknzQK8WnC9YiouQWYd6BeOPeb2KOufamgFFR+NhNMVvyEm
iu80JP//6D3HBcWQ77RQZiyY+42lwJuSLm7oVmRtuSBINfxfkq/i80TlFktwDb666spXIMRL4Ss1
CcOV4QsA97MgGgphXnVyOH55g2rNkXS6sIbgLL0HkuF41ZIdeYBPTrjZJjolREYOHtKfmf9Xpstp
e74exkKwoH7+jZnEMfHI135GXp15opzJ1LW7CddNphYQpbWiIbwFofo9NFt75p4VuIM+xvEdVezn
tQf4S7wH4UiWkmvrOlEjxIGzhQbgq8xD6GZm+zHMQ7GqJLItsWBBWFdRkpl0C8YzROaDshiE0i9R
9OKCWhq1q5vTLdiMOj5cql4hYI0q5Nz5AoDCmDnW+fuglCeqw6s1+Asmx0yiBqFEHleD1Wlsx3MN
UQNb+3zcTaRqj+nTXNMXjw4uKFlmaIEUeTTOpTWGLX6MVHUHx1YEb+ZMt4uut5FJYvGn//84RGDx
sneXI08P+8gJLp0xQ48/xP7JeunZ2+/d5N60GJfL4YT0THrEpHCRVsJHhDfbFcKRqmtvjPS1Bv0L
RbLEz408XoBSwWiiPfbapweS9R8IuX1Ws0p7emVmEKklLBn3+W9qqrii2nUQIDoS8xdZSRO92lAL
xwXUzmr6xUFQjsNAsStFpJe0UlYMNBcyOfyAm4TvGQtng53QBowdWpWW88i3SfoJDdmI5xnurf/+
zwz23FOmv4cEDN+wGQ8ssfpaMWJOQLuq7n42KZatw6sXn2Njfeffcg8ihxtMnPxCSJMh+elFEvS9
vmHkHuZYXbh6Sa6/2fFmlV+7cB9Mnzg4le4JtiH+fWvRRGzMQo+73fyc3CemwW8ljco9w7itW9Z9
3M8T3sE0T6TvYYZk8C0b86NirNEH+9TGN7ZKoCC4HzLz9aJhAqkLznMLDEkT357XMBu+yZT4Xu2e
pyBC4BJ2sBSfp0RPcTPWFPMDLmAksPdwoHLHUWhxtvonY93vWmmCEfi2grnlwm/JOUOkpd3T5H4E
bsz9Bd91kGH4PXE1eR6E+RGiIBZ+WkvQx0HSMR14hBHurKw5R12apfeHzdoAjtuhbvcGQWuPWIP+
95k6vOEfRD6yS6tCnsAhYiNkdlGGVBi2s6ntDc97FB46uRPYvf1+JOFMmSQGgSCw/xPyRXbjNVK+
yb4SjQ8mk/AkdQWJXr9LfTKfmz1VhgzP5WUzg5lyLwSFpdwVM3Ayy3hTbInZpYn0E4UqYXePyNxM
fgaNhIXN/Slcaf8W0RLOT/P1/K/nIGHOqaT2Em8/ya22zEfnmJBSXb3Thq9NOcz1fuqpjTKcJmPV
ayjUwJE2j7aeRGpfhc44bwCnF3/apNPQPq0b+x5nWvuja9M6JFIh7C81RW01cwzg1vTpDNFQTt6R
LoUQHgTxtp2rW60qOkovNokPQkMZt1J9a1dPDr5TT8mSUkGGzoFHMnayzGXtbrv5BzOtYUXbGxKG
CyVfj0Smsk4ceDuOz3ypIKOakf4iKRfBU+QDOCXi8wCjbNiECfS90LZRZ9trf36wcVGbYwWtEVW1
KLBfZDgS12mOxdAG6ZLOkKU2MFQUZNEWALCbigvDD+vReXqdvRmHFzPLL41CXUeYjMrg/76gf3hi
k9ldh58kSVCbH/iytsJopfBZ+LO0uz3sS0QS8Zzv76zxKICH223+71V38+aAQv00lPpw56oEvZZK
KcgeIZEEWgBwRBzdkDDy/XL3zsl8KJ4TErc0eo1jdFuDxjaG1BngO+wN2sJ4qgbzB84ITY9Hxz3r
Az742hnAr8loUNkk6lfCGR60HuwK8Y92MCvR7scu7xoin5OGo+KoetA1bC3tqq9Z/yj6sUFE2Jqc
iPvAzKAH2zLongnbrvxh9BSoBTI8c/VA4iF8rBiySjztaWH0jgo7YaXDXRoHq3CfSM2BMuZfBBlj
aJBo9dRT6+LaxvBS97N2H14BF7FmnkPRFjsfQLlf+ZvHU7GbmBYuqlx37GGyuok1FmfzUbPZcpst
Guqs5QZsc1YdoxZjVXnjXZVLpKml9yUIb5VexGntIh10oZk6NE5nKfGZyl5CoWzDxbt41X5TRyI9
glYE4bqz4K/6eXB0P2miRPpoZNW/PSgyrP3tBl3PIv2vMiav0Z+HIxz9xRiNO2mT3zFwBJHgjjh+
eoyyBYY4SKAiHqG10arTJcD5Z0+7qB0mdh1LBoyVmjcFZX2YvsKAN/VY1JRFC+jK5PywuV6sovlz
sdZy4iLCkf5Ja0WZYK5vDlHpyz8prq7O6CARob8p1zHQGXj0fpyZMGl4vYcKqwnX0zfNFY5bIDzQ
q9Mx3YgjoIK8WSazIS5GR1iRZDFU1vIxXSuxlVxi0Z+3Zwgin97YXkU8Z0Ri5cNmjsT5PGN3e5TK
79OvKzJVOzL34WGl9Ev1cmE1zrQd87nLZZC5Z2MKkOKvdo8AsDVLK0ayxrjUlaU9ayOd67n5bwK6
KwKXzMpYqDw/8m1Je6BFnzPSjfJo+lS9FE6Nmqx8Ld2TfZ0UizCfJPQmiuYPR6SPGhz2M86KuWEu
lQ/U1Du6rROuH6ZFBwwM0w6uGwpDkxuCb8SAKRLto1Jv8KkmEp1SVQPzb6ke53dFxQ9ujcoJs12v
ngM4RVjG9V5b9KLJX02miVp7rFQ64LmCTFFut7KbJiBtpQKWhbFIdl9wXMdPGbStXcmb+Uewiac5
lmgKVkg4kjsQEd0WO6JvsEizedFTGnwT/w0Mq4lt5i0YYSxWLNFQQPPfQcCibwWdVkeoXIRQL1PZ
gOI0xGadIAcX7hPJaj/P8d+SW3F0XPfHD972GYnduBmLbsl8MVL/GrLoFRV/cqRVBhB7NDj0++Rm
TJ/r2LYmkCs/wEnyZZmnE8Zy8C9vWnEdA3AGmiIiR4HJEh0xR3p8z0Nl5/McsRZLxYbjAkUP1gtW
lUO74WGYdnOSXPOY0vvlNTawuCeAs+gQEAH/WK+75n6dXy26HJCIw90hRP0yqzVepqq44GiwKWD1
EafLpOCJdCbmZx5xSOkSk6SUMCbu/sH6SpeyY4b2D7th1MLql/XDd2xs/8oeNAiCWPjF0K7C1EeY
GQvfJc/qnKSNwSTRfmQOWoGedy5m2u1oLZOJzta+d6EtXiNj/c7qhAGgEHZQVjs6QP79fyJ9knDc
p4Lxcy6UOiixDpwcJOY5jPjispNxyOy5dRATrY95guhKJA0OFNEtcgiYWBZZAbIMIMX/t5B19fdy
5ofq+hXoxAaVJcDNLDrH6Xu6LqP1wjXA1ov3QcFwURivdQy6p2HJmsdTCprwcYZo6XrJIoUZv52l
Sqpgaq9uhqM95LGb/q3tjRMzV4/RruNFzWY0rleAfFUOpPUiAU8I7IJX/iWraOGVvZ+7m3G5j/OK
kODesZyKXZWyH+UCqGGvrcPR/IzkxyykfF27Z09fHekzCsZXwX3WjZQH7LDcN7fKa/LYMU2tMT8Y
rqosfo86VTSShRklYJPKM8AjbAHolRwFlUK9J63dIrD1hUp+zepEP0DUlp7e7xkfji/uWDRDKwb/
gCBcOIY/VN+2DpOx1JzgmcwwTwtkvMFzgK+2ikZT3QMc42CAhwwochYSL4dqaD3W7KWSTYqJs4c2
yQmyA49kuyuk0fcKf4J/k5vXwRMqxGBq6ktfDKdcqsJblgfa+XbdBSFb8qXR3MBF1tOKnAtqcGQ9
yjdvyzvdCow/jgrplgKrYQ7Fmx6OFor3jny9pDVbLJKl93ogoAHqzp4W719COvv0Il9fL6g2oAje
R34ruyEpxwIQwHalo0yGeepT4Zw1XARYWzTa6wxhyuq0DxdwHeZNm5pMYVIh3iQd/zkgdNjHC0FY
hpGU/3k0XGvgnXPjClP0mJMU6lsvCBwo6tBTAscwm9tDKlFA/im2JZWUyLjncfH8dOYJJFTF5KsG
6Rv6valErUBtAF0B+qqSIxYTxK4wDM0GA4omGhPff3tgmatnaTMr+p6qjMEuYzbzc4waBT1uq1/2
aZ7uy5m0FwQrBKv/pE/ua9bdDVIyMIiXY5Tu+P3HtPk+YRiqlGUHW9YDwxiLRdQiYML3FHcT7TC8
fT4faMUTMXAc4NFq3PGHYWAhSVDf5nYpDekTxLHz+qKCVPszU/Oqpe97T0LVXDbeIrUtcZsklJNY
bS/N+ME3o+Q7UpUFZVJnaE+e+lZmrM0AAhj86chb0wi7fnL2EWpBvRocuH0g8TikDWHzm28XRji3
9Ea2n30Vkx3NyQAINtdkeXfc4323oEPHQCODGRsc8izui65ai8C6lA2CVgF5wl1KFRgTf2yOQG7T
Fl2JwhRpfXDa1QZxQH8lMSR1yP/REyr04bfl7X+YF0mxKfCF2VmADByV51g5WQTT2VfAmTv7uwY/
oXRvMsW+JUpWhnI3g//I3d9s5hmhAvx/FMAlF6mdlHB2UTV3tsvnzyzAxPLJfqf8AzjqrAPDIvfJ
n8Znpc9vB2GiU22Z0LaHgGBIfvRt7qs/eHUQcrgGcNwj1xIb8Pg8wFY1diN68q/ZViEl7thNk1W1
kdyZERxoBJgMhTueFYw5nSnNtmQUNjxXGyyUMGkidNa/2602KL8hBLR7Ywx1RvmujAv9VbNAalib
ENl9MlzCs12tqPIvXRsRLzlzMz7WwwqRvDYH2qv1wPUE1Mrb9C6/XHc+e4NiY866okt0QKsD8Xhr
SipvsFKBMUWhE5aTM891YWSKWp4qyWxDBfYBNk4I8DeRuqa+w7hiL6Veu+hnQDBLGo+bVO/fsX6Y
1BXzIJenyNW7KVK9dLOmIVkWpKmtDPENj+tvJzezmgVM+2piVDPPEIJSSE7u1sZvhbLNxgB9Fd1f
C3GXDMAqM/gyHjdaHYkr1USLX6l9WCLvalGBdGX4B2ty/1qWsNl+X2Rk8bUoiUahQST01/+9X1/i
nAJbfOlP+OT8dpdv4ctxQCKeWMsCzT3q20Jdmv6h0LGPLfg4vQEbkHbn3VcobbedOaEVsPsx7Jlk
pVWaBXCU8jVYYGAuG8FMfW0MsKDXQ+RgnB+TLRYd9tlaaKhgFaIVxSxddsgqltkC8IfXvxtC5Bpn
/GRzmv4O6BtYKZNrHmOe0+69ptqIR/k98zPvFbW0LfCMoXT2j9cS/x+b0oOMPuAJUkw5QxIQGTAY
P6VBKOBvS859+tyAB10WRHjifq61Ebh0YcgRgP2NEkGKevVjz9PmIzhTqj3OkInhZOA366DYaAzA
/senU4P47HTGjVskzzEXgjNRHXGP+z9hrwB8ykBog+o0nCEDVIR8u7RtH9C5QP2vtXO91LT+3fr2
AsqO411CbCDnd+gCwaNP0SDNq2JSZO9pFTMXqEO0WPUowfUBEFxyhFtEOKmY6bNJTC09TEEVUHC7
2twm45ekW/ggbdDg7KmqyLmWSXFfmh3ZEIqqsKUf+mk31WcsF6KD/oZxJoGo/Mil7brPmgv770Q8
4hNyGlGAvbr1OvFZWDoSntmEc8t1/pcWNnhCSL/NjJAYk9OXQgFhMYJbYye9HznEiCRYzVD8fIPH
Se5j0QBezMnFBDg8D4syQKBYVgUt9wUxWbTZrH3bX8y4/TwK3SwgpED6aCgCR6odxuk56FJ+j4vP
vcqb0wISOhY43vBGKU1uMscxvPRqQIuEmidCTukBEqxKXjSfIYikXYCMZbIylripeZnJIUL6JOA3
oqNx3GsXv5uVs5gADuqDU03i1S4qXjrG82snFsOvfZHr7gnQVUOJ2Y+nTVokOc9zOSoQJPoO9ll0
Q0TNfaCausZWzJeu0/4KBNJbtghPIfazICNsQiKnxoX1d3i/lf8BYmYbq1nMPWGkw7nf+auKidzc
USWtvIBH7b1O7ZU7Vaa6iEnaJCJB+Xa5Uq8H1bglf1OFqe2pDLIIVKG2TKij69W8XC/A7z33xIe3
XEqnteMSoAMdSVBn+YE8POQQNoo9ag0ce9/Ci10iJmiSRPTUhed6oH8xJqhKsankiusIhcR4zEA4
Xl4PPle7lbW87scWUrptHjv+aLlTsTO/7kWFfIOD/4nYifG3MWXbdtygBd9l0gmB2x4zqTqTbifM
yAVN71DlPCVJ0AFpUEOGHisXZTdf2lE+HPH1yThIQCK+Z1ss0YCFdl5XBsN6fbBlTnDgbjMzW3oM
m3rPWTJw1tgJBvtyYobsd+NnmmB9ITrcserxVHdD1UT3CPVClWAoeuiIwsQBDSt3ru3oFn8XYsVi
9xgs/5PDVX1wudg6qghjhlatRr+XvSalJYRuqAAaZHD7efuwLV2/zNaeF1JfF/uZ//Iw+wEQ5c39
giFRYGv1Mu2QzJs06tk5EuDMYrnR1Is5ckEIcYgszXZlT98DChQxCXKK8yklaBqcnFlHklfsq51B
tnisC2hU/zwHkSskfPmIQBQrFOeUkhXeEBqjYFSV6PIVAqxAf9X/p4ivx/ZVuFLxi3KSMtu+lVsQ
t9ZqkfROipZhX4/wkHjofCR9htRtTNo1GX7zAtZlTfP0VPwhVOWO9PLzLh+ZzW8FJ756ccNrBlkC
55rCDxD0MPoeXRjGFv2U/qfhtjhxxGhIRlml54J+QGfPyAnMGg+0ALLhV9vTYFt8ZVCUO/O6vhfo
7pM/hIixUV0pjMMJri7wJWgn23q/sC6wGt22Sc5iIZox81yZ+ZpaAW6Vw/KN77ZmuMHmPHZmXXm+
6OxeL+ivIomaouyhmWW8195CKUkTH39jb7ctGoQW/PT+Jv+dMCbCjivJvP93u2N/9IhG00LNoGPQ
Hgiwsb2cw4XVJpJhB+4UFoDarjg4+/ggpdLc2s8HJtYO9eXgQS7KNVKBbhGiEzJvqUD/nr9QclsQ
1GVZs7yoQmPFk4Q3oym5ebfZjTPISN3xS0s0iIIf6WC0YvS7+uM52EpauayZn5su1sYxzxAW21Bl
QFFmaRpFzrzQ76YjVLej9Y91q5QpwduVUNj8/KADYFO6GNBw+ZeDRjzn0/77am4WLATbZWIdb+tx
n3mP8J7/54W7N1xL0QNPwyazczI7PqoxO8iX064Lj2B7ZMP9tn7TE+Ex4pcyQHkUqLYg/ALWe/3b
0IfP27tIuxjxuJ1T7rUzIyzmgbDq2gErN+V/lrio7j8Lqj9TlZ5OkUvsybSKHQf321tpTDy12YEq
eweO78dESostOwyQyIy5WUYOTKn2wysJfYSrQXfzIvW4Cz4FcXFdmkKOklljFlnmpaS4OeNfxjak
9EO3Z27Trs+yRYJSSl1eypWztLgg/1Dzzp7/KqeOKI4OPKA8C3hA3hvQ02Gwqpn2gEqUG8QBPevV
fuxOUeBj8NjNfugA6AxarJqmvOiCzUtrOunAgHDcPJOBdyD7eF2MKoGL1s+p6d3D98Qr2CuXdCza
eD0DrUqdUSU9OWF/oiQfXzMQWU9IA9fLvWY6jMqnXfzi7DEkvaMPZOXDqOI4xdKsSS63PicGEX91
x8csp+VYhz8smV+s319ylVdu5AiKTUmjyzrsJLlG5Oy3NePRO31mWmGET/WYA62KA6yoMGEsSv9M
VSxfSWeABT2DS6quRWrgtQJoiE0kqBIc+1oaW8lRi6YnNXgBLiioIutC3BzW5tD2gWSt1np8mUlb
QhOQ8C6gvLm+IaBoKs1gLKNdIjSl/VRdbI2lXxuzbjfJVjDtKMMoNjf44ROr5LyseODQWgLy3z6A
aPFulaEvA5QUOuqRJfpBbd0BebHk44uQkNc52+XC1oP6dM5hLQeAsgJgrmj3qRJOFoO1Q7wWBYVN
GjWQRCMHxxr9VctXcbIcu7GJwFlgRgMwv8OH7uSCeVs5JA2bYtqEV8paWM46dhxF3WUltsIBfCDN
fGgZuo55n/Nf9oExI4rMjlb8ZFZFgSIC8ja8nn9WLHgEiouHkwOUgAC5tM5wCDMMre9Ppnw+cy5i
3nWiKmO3oezNTpesxYXzE00he580PY1NmHNmMz3QRqTnPfk700dHhDfrVwfAJJNDrUwpbfP4Lhxe
odSWvEu+TJtmbjcPmLIJjl46qXsT9faYPL8Ve6ErpCVLcPr9Dh04HOAKKFOF6+Rif1xbjBLE1DSn
Fn3vkLM47jxPP+IhHQFeeWS69TqNdQ+JexJWRrGTQs941jhvX3ClWdu1igrN/M4PNd1f6JHotWsA
qoEOx5DTvvMPrMziTTzPiFXSslUAYZcF+7SZkKA4IecaqJOXwVfCPbv4VRsbUByDVJwUHFgI0GGh
Xi2XvQirZA7NZdLJ9S4vIEt9q9Tgz1KzV7RrJVVxSJUnz5aGxpDmKs5S/J/ojhmT+aZuBINWdgEx
BQ2ey26ZTUqxgs0NPx416wDgp8T+wkZd4SHN31qtq/kDxONkq+ebt7Zm8L/Wv8Bxf0cW6rU9+5NU
cyIL5JezSf4cqTNM8w20LuZ01j1Dy4det0GVus5NG5/jqYvcWAIANSk1PmvHSKUqp6gZMasiCYp8
p8p+3cGvbHSobszgcJX6lBRrWbNG1kMNN/+vvNhd+rLY9vsa2SJgIzu6LI8sG1qMsG+FljYWNTuN
b0UpRoIhLRpjEp2xqX6Lh+dHjgnl/0xTgZkmPKMmomrTY3PCeutKMV9yN8ibT6P4RGFICmkw3ZLo
41Mf8gdTECy4sL094X9M5+oG1xl90vREyWNjyw+tscLax0gwFNUsTMTqCbY5S4LYB9X4yCv0m2nj
dBzOB/2Gcakd7Oj8ummCyLBXhamyll0S4DZCWx815qt+OITFa/HCXjNGBz1wrcAgrEGDVE3EwYK7
8nw8O9VNmYBLKhTnIOyrJsj8GiHONlE4brE8SD9b96U8Uqme6AfnBeDks6BRMCauohBGLtvwokMk
bO9RpkLwaXmQtWGBRSC9brWGWiz6//hZ+mT66r4pTlWVhW8FS/wrSXnsi9D2Uzp+Jak2/6VoT0qc
rPwihtgiI5Q8yEQgUsdg/oYY3gwysoaIkNtyGiHBNVNLUg/W0hRr/Fxc0DY16Z3ctwGOm9ZTS+QT
0UwRFj8eDpdbUn67MV2oUbux6HDvwhZHPM9fAFprKwmA/VUcUg39FJtiGSImLfyQ6oJvLynqoMo9
ZRSh00qOPvkgL/+4Tqf2O3fy7fZvOwRca8G+FOKPDUCB2BJ6K8fDW6VAXLzyiGUhSaqm0tgQAssw
WHaEgWH+Ds6wch2xVnhB7b9Fe1FBAZqmg6BZXqWQTnOUS8vDxB32YZt5SHEEW4CCg7vUCeBgFzX0
Hls6zcuXEvJmN38GuDIp1P6yVxcrnLYrAxLfoHqwuUKNg2D0ki6cWQC1Wi673ryqcphPRdFXUI92
xDc8gn+A19YoxNFuqJ+l+7h+njjmEATa6Y6/52Bz93G1UTVL2m0Ho2mrM+PO6Zzdf1C1SfSMZkpX
vK7S4dT8mn7BokchzEbQTule/BhO95FUkYz7M0C0IRjOpxaKgkmic1TIR/blp9xPp5MGPenbwjB/
L6CL2o+AM/eqS00AE/DYbrn3dqQqyIJDdf9O11BGYZMar65x9T7OP99ItCQf2SS7qC1omNCeJ06E
jM+pmvF0ULLmfspmmgMDEd80Dnyw0/fixwYue9V7a9HVVeFZo21LOBLfXuM0U7bpWqU3W8ztLf7+
qlkAEspNDHAmnH3/KvHOfhbLgIjMo/RK1aeCCJhoff/xf/ZlLzzcUeiKqkv6gefwuks39ZbaDPCQ
NZ2aLImgRcHoN7yXtdvzusOJq/HKAcbjrtrm1LCazEHeAYvJ6XB+5uaZc//AWTAiGTmtea8ototv
m4SgQhhWR3WsOW6Z6hiSy9Pm+4gXByyQZe+EgkQNalb12q1kPbGhMWPTGvjFzdwVOo+TXVn3CIsw
roGGOj4b0m0t4MGxF5jAFSVcUpeczyU1LRFYUT6fbCtVSFx9fSam8yr60I2F9+xN3l8pKRQWZA9i
0lOQrtCJl9Zt06DghGnbOq0MV6M36NM+IpZb7NJBlvevL9BZlYe0VF0a5wx0nfMgI1VgqZwNAt5M
9eQvGNCNMDnj1SJlyFym9KmSo/U/ffcGxNqzBYEyuGgloo4McuRfgdraaR/kL6/nAPF/Y7YMG+k/
N0M5gtPEz4E4VPHl+kCrAgAPzXxIeSMvKhRc4w+W+xER4lox8v31WYgMryFqJ3Rf8SVq5hCkelQb
f9jx85a7SaP5vynDK9otwECWwpF8LrP1bhDaKsd5h3G9ux893qdRrigFnCdpqxdQz4u1O/1gAH3h
LrbPe4YoYx6zPatt3CKEbC0InPMvywQfJEyTvok2gKyIX/REwB5nA8AYfEzE2DVNP00yuOa1hEYC
zD7n6c+9MtlQqttFl5ACAbF9ELLKceXBZ/oa7eBdTHTpQWhjI0eqx+a6oth8uJE2xdocHLzg0mNc
lhnra7W1KVeEQi0YR4QXO8OwGT6jKNRZ1RHk25tWjwOQyuMz8Qu6BegFmU46WjmV8/qnfeDdamNz
S5L8lbFN2I4y/e3Mtg0wluolBR+4okyjbFsJMRuE6QreGszx+x6uyFzlE2dj3oglFzH/FukE4K7E
gtC76p9xl7Kk75B//l+mmjFA0X/OMr805m3qgoW64pGqVLp9hOXy6Uia0WowkM+1aj9QM871JIAO
MtB6xYVYJGRuTPsfFyZMki6vf6W/2PVj7L+TdBhTAai+MLgnnRGUQlWXbphrWZZ5SoQSbnh+JRyA
bUxgbW7cz2KhloUVa6MC9WK4W0CjHfEgZxvGogVhDWhfvHdmaA1b/p2/a6k1oeBAp5t9XUiuk/J4
zj7hL95ZU63OG1UNWLwuqBW4UbBBH3IcUnm+jFMWd001UTMHzNvCNuRWSrkCRMuJtgwzGbFXy0Nc
/cPVXawoB0bslaRD4rJKD/5bFuL0j6gKiZtIZtIgFurUE/s/p/NI0ypaLgZyiJNJzOI7JE75mxul
pMGSSC9yi5x0mcvsiFLAVHpbDc2KpxtGqx28CZziTUX1HVoZnKu5CULXBZJK31s7oFbH33y2nVLe
Hy9NWhI9mE1iAQlNVVcoMXLqaRwjPQOYBms6kdkyncZL/m9TiIsQoYo1p4XVCl6j3WmCJs00txB2
TtFM7YTdWmh+e6IR6Qs5Or9AjSOiABUZP4EREJ/yz8v3Ue5yGIRW/kf992VuG7TdeHI8Ist4IXtL
F9uiz1f5F3hhEARHJhaNfwdvgNc4lWJD+nKn4tUO9u3Vm8GlZ5v0dvBOS6xasTNszEK31Y7KH7CG
4gICUxIJq57A2hkhWVQ5jCl2fFzfowM/ZE1zvl+54GDmCV/RTaOC6K9YcBv+lNY7HuuwtRJxEuXs
wlS2VnKAGzOWx218qNjvOyioP3Asqjd0t67Gy7zTtUYyFH7TgqKD9l+k24O0OqU7nXuKvQKUDcH9
wPWrWRw2MlXZDaF57J+vgXCLsHDVmYaAL/8TkHWd6qUR0K2D2PLfUwoCBSI5q33bsf9u8hLsN0JY
4LQZUNMtBOQgDUFgjFzYfZN5QqpyiLEUGO62XAJJ4MXqg8uHvqOgZw7TsK2oA+jJ9S2Y1ycQs+ZZ
DOFULMBXu1rpCAmVK4Ow2nwI0wvBt2w6LJcBJZaxqP1oFw68xRx5icNKzH4Whd8SeFjPw8xa6d3f
qNS9jSVTS6QD/oBqWVN7V7GRGP5XQsDOM0bWXljE49B+l24AyDPdjNEpdeHpnlDSa+Bt00+WAlqb
ennrtit/PgwRvmaaqlUCkn/IuAGFuXvpCZ/j4hhqMlygvTsPbKNDXv8p8QjKPt8VDUwCasD+qMep
t3AvItx6Yki2ggWNIMvCdBvVXhlG1HoGtEqtKnG+Q8m+ZNGHZehIg0s5fBZpyTIgDXudi0lYZbGp
51453oNq6rPluQtGvuoCxze+7W++X4XpmxBbtqM/UJHGXMcoTXMxtFFo1gjNt9HJchN9trnsE6Qw
X6exclp32Hy8Fok8waDk0PQw3AuMUcb5vrch7m1hRY3E1Bui4j5Ylb1bqlb6xwf+SwGkSU3itAkk
ivgo86qHlQoWXUclvXjkFd2Mw0SHc2nIPwr8qFzPJlyDcnEfLEwM7VAy7xAIX5kMw8HxT0FSa3gx
li9YfVhiOTXeNoOzKyLxH74z/6AIKHlfk/xYa9u+n0mwqWwjsrIy2CxKN5rwyUizITdS6cEY6lM0
a1LM+4Sr+n2XtCbvRgz/3fo6+60j+c1kvBeDvk3yCUICRnE40L4lWc29MLzk0lR5PxNzKc7rM/h5
7Oh+tAH4UsI1xzTnz4gIxkOyvSt90wMY5q0jlJhfhHYGZ2kIsOo6wMovyP7NWejONeSfTUKqd8CG
LfzDf+MnTkvJgbj7bcSX+1MJDyZQ3z/EnAqe3UeK7tdjLuL5+tYTMC1E87zDVI2/vrgI5LTLwJIW
GuDfjfRJWBF2uxnNaMtrWJ93osnupN6MMhK5+1hXaHh0Boxf41lelTfjAQXXpLNj4xcqExpVJ5+A
MFkS0UnqOeWOG2yHehwpTl0Vpv4SWWvMARPV7GHwIbYPfMlJDly7x85TnlGJuQe9BBaldeX+HWFG
27KjHd65Vk41FYUWxno3nDe0xWrOIGuaFfH7U32SlnuHH6kFRm4xtCyisPdplrZt+hOXyMKzkWD8
veHqgWM1pr5h09nSHDTyrMwD9KRG47+f1kDQv5XLQrtCYc71c6wIpr6V2R8CLYZ1yyoQXlfLB9NA
CkLM04aoRSuJwcbee35U5l/CXHI9JmntidkhUNkOFJN8NdKpDpSZxE4nOReGaiY2UwK88WPhLTOY
gTMTYbhkqYTX6UVPQBcw3WR4YmgbZReDGgeR1q24JdosN4CrEGEC7Z771QfH6n2kt8eBSF9f5IXX
njWrc3c8Jq8CydofYZ53Fw7ZKiOmH/X5epTYWcCAtmhT/FtEdkmGatG/9c214PXHVqua6EpQRweD
mDX+bMgre48ZCFIMxNqVTv+xpgSuKdmPJy2STSvze8Lvnf1z6hHNoVRiRmgDq1+4EdfTB1mtKZz2
PpU2jMTuJkeoA8aQDnRY3EGkmhHmeD4DLcWZkE7+eTI7mPrGgOeSkjDFfZFE5BWiVImNSvp8ZpkF
7o7HhTFns6NUX6eO4Unr1vFybqnkiY45NekFtyIShu0VhQaZ8XAhVOavABbstSLdKKsMnZWJlekE
gIWSLjNYRm95orYI0xoAsSOyIHLut7Bnpu90wiKKaGPk62hFm5sGhUuKXRMrPJ7H4nQ6Pejyj2lc
crD5jxyOcT++FPL0iUujaAOLBV4dxfT4ay6kp06mRqlpvo0bGHjtRHk46P5EbyvNlUuenzP8SWs5
VJgY50kipQ4WolnytqnrpRd9b3Qz2GwJzHpa70TU/wbzcXhtX+BZjY0swiyCywCM1Z0JDsWHuX27
6rKWH67GO/R5exIwhJKimCfcckl+5Or1SbY532JprKjfH5UWgPgaDlW3MK2u6kKKkeWt3iDOZgR6
Zo08fuaXlAT5SxPjv1q2nyoHY79KNwKGKCERJATnVvLFdaQKTEbhGVwKm3T+82NUzypG0uvzra07
Lh734h9oNZTn62fMrjpIGoXd1cFsn/xgNtzLCzl5wptCbYTnaj+O6ib0P3PAEJ/Be4bhRsMHtnof
nEyySIekdYC3VIPhhI8NuL77wpBApCiEqcW1ZZ8EoHOIkaeYqjETmpJbf/29QECMcfj2H2ZXhjLG
G4I6gF/pmNEcwmidVfRFn+gvv/Gj9RS6eBXGgskeEMtwZ+8YS+CaclUGkGqtNPkH0NbnwCvky6Lx
wnvbWdZhQFyUvN2oJMS3zRmGHrZdeUO1SrbwFHuvi7gryKQKF4Adcpi6oKuft5sTfX5/I1ONnIUt
T7HCFvIbXxdpqp/ubcKm4PvrE/jaXLDobKlKJyZrQ5v4jMULWC6nSVS+G2RLHFxCqYXYviOEVSRA
X25PPePiwqmntV9tDZAo1KWanypuRkQi0DXwPBS7Qwpj8Urtr4kWxLoxmSxNPa6QrQkjIOectLf8
gPS5/zFl7OeXQg4Bo4Iz2woJiv6pNF+ux/PPJARSkcjNVasVsgN+vf4rz73wT5eS3wKByjf5halo
R/ZKf1oFuWOJOnJI/a9D97V9nLRVHfkawyHBjMVRzI1vVVlIP2jJIOMnmFZCj6ZZqa5FTy/KT2JE
Pl4P0MUys4j46/HD18ADRGR/3HzEZCvsSNq1FRDGIpS0VfHg6yMbJvJ6tlWhl0DZ1nXuyTjNQamk
dyAk6Vlu4g5wy9lLEVm/IpmgmT/b38AoKltebILBVuWHM150Wp9B+s6y/c2IWMru2GTwFCZIx6R6
nf6A+BvdfrcOJASvGg3izaiB77W+GICk26Cj9dMdkwGX5i7viakXHJSwKnsCi22jlBCF3X1tInIh
/obRU+td70zex72HKcXdFahi2OHzBg+WUfLJAn8QDQ68eGkXJmBYTREAJICwlzVx3oY/woyHY5Is
wl4cFQbsYL4q8MRNOrMn0Pfpcmiyk9jE7eddW8DClwG1SBSmV6R/q6HACZUiPNUKHavmtX5/nsdc
zzXcQSEmzHIk2CPZ23+38edUmdZYA8Ax4x1R2l714Ve/sLYNDUAda8XYwrYnA3CXcF7x7KEgf1c7
LdU0ts09hg8ZfZ954hgjVdif+icX6fWbucAcID+jT+LbdusRfAjyQ0Xp0Zq4JhmvI3AAzuU5X+I3
yD6i8QBAVi097b2evf7X7NVkmhpH/aD8iaIjpl8ztGZpEvF4rYvnMsRZhtWQ6l8SXGyvrtXp1zX5
T1mgVM/XQztu8kh4ikBEOJEP8nt+hnq5Nvts1Qxz6XnJQjp+GfsFVBb+Nv+M+tp4/ia+r4Rsb/e7
/4K8dFcxNo7z16uHOEdEakPt7yup9m9Qr9EJ+qc3B7SxL3V/OqpgJcrUcaikrOExQ+g2G4bcNEps
aVhyZSZlUEJicnK8HwhfUrAoy3TtdO6FJOmQVx7FUt2TEGVL8h7ch/oqUhFAPY9DG8fFBGHoayqt
h4FHP1Rn/lFgMLlqAZdH7q4EHFglMvbgzk2ITsjkaJjWU80iqPj0VqmCgihszzt3dlSgCJuJY500
z9izxvkC2ef7fbBM2p5/r0Bmc4bmBUow7baDxrKHFKwqlgdCXBuLenkF1JsqeVH+jBCdRRx3SMlD
XreHDgCr51Vj7vgItxBnVsEjY7uNyAFEYJDVeulUKxmTXX6rImd2s9Aw2AIP3HH1Ld64uIl8s/qU
aJwvytvgMe14l+BdCj9l1PYhHGNiAkwIzkWSud8SRJdMLx4U1jIel1t8+Uo0xlbYtaLdKrAwUsQ4
PPCJ31MRyuY4AS8NmsMt3x6uXOz9FgdKxjRC9tvT3bRGqpMDGT8VvjZTV1hJEoF3P2cd40jG99gy
dTwdxP8VlkcQl2k2svrdLkpgLYhcnLSq1U8g9Q9J+9ZWJyTGf0id+1yWn/Ak7HjsvS5CtFUDPjdT
skT1z3MgwIUvr68z/M8Kez6FRVwHpdl9c1X97LYUZ/7QMS1xzTJKPOys14d5RhyE/10sHSZE9c1N
YLIZ5r3W7kc1wLTahRBclJpN3i0RjyEhAjVyR3ZDb1+ysFIWKQYssKZ2pvkcaQIml15U4VmIMaME
9M8Bn8SV3diQx9j7N8Y5Mg2hVDV9EHuNC3ktLGeFVSgNWoT9Yb6HCh0QyDGnYIXD4g59Jgbby+Z3
WDRXuyy6y7ICxkjQ+2kAGwF6gMRP02Pgeib0J8A7EzLAmdj8ua3r8nlnkM+F2veAxoTkJKRlwrFa
ftHUtVvuoFvMpuvRt+TdKnHRw0Tx7m1Kuvq2dCG6/VlgLhEl8QYsTPaEjDNo+IJ59DZRIovxZjPD
uQ6THaF8VoEK9bDPA3z5q+XLSeGzrxW7vNj24z47tAPkkoIKrxRgbroCzWjJiIbZyQzaHDrAN/C9
CVU6bl9uwMpJ13J5QJk4HJlK+RjfshSLX+h1aZ1PyaHaSOjSpoLWN2N312M+vd6rG3wz8eYnroYa
d3Z2j9kcCXP/SReyF5O4E5X5nGs0DvUTQsw0SnGl2Lo17RuwOjKJz9M99lTRe5A0kXltMVl9VwzV
x4zm5jgkcvbs5ZT7M8IACOSL3/Lb9Ij06wwHDp20MEg5yHbfxtY7uYBsphDxmBOeU7Dhkx9JcmZl
B1PhptNjvX/n+2DxzTJ/MYG+tGG0wpUpGGujhd1eQl5KzSLUkGG8lxlhltbJis4hUuduTkK41Ylt
X2KD9LQJz4J+PG8oITJRGCm8Fo1uXOnj+jzmrt1GsnrLj0rE2xcPbeZLWM7Mhk/QtY9NKkTxKg8K
JvCYJb2eHCjTToqPc2qzXQpeGS+yLUOUy8/1Xw3jgIw2oTba9wj1p9v+iLVLOgHVQ2aT0QgxhDSj
Rzwaz1F69Xp9TC3+hW7ulL4UZnZj+bUMPpf6fvOz2n0OvtGJT8xZ+fIhBn9OfSTgtpPhjA+JqJn4
GizBSy/EI70vaLbMlT3xmUifYe4wlOS476FAsPOy2R6AcYWROH3HN/XPG3wG7dQucxdWTfwO5BaT
yP/iqzXB5RLpDsCiAR78Ome7pkD0cLQwEIbuVfPoLTDVE515WAUOIoV3c57DQoFzcnsBvRWhvowV
3bhn8Mc1ZmrQaWKQSOuJbcHyOhmIhqT3VuWBNU/3Kx0T2cjElvwhvQOJhIiAtewKpq1WcKtOUTPU
2p/s7bISt46Db71++9vPTxrci/jXNhmUdEvwMgvEVaB5Ap33B9p318oCrOLgGnfXKyhPQSC5o4ct
kfhitWPBnPoTdai9WdQdFJuqb8YfUBiIgjsA8V7E8nHleM1lI7bLq4PGm1pIUYS9+UlXmAr4mAm9
6Q6IgC/zOrm1Ai0Yq+ZB3r6G/lkWKVMPWbEZXZkNz9bbb25AthzSODczfMfg+aw40H4HDiZqANYK
zrMAD5HoiLYJbJs7EK+BhVTChpZ+bZe/L5XpYMeICNUy4CyfRy8bflFp0VJPTDXim+6R6wNZhz7U
SfgGYzhoD6VlhteWrIty02r059d1fLdyNwWaV1GFwMMwu+0396KDBhcKzYjIUPWPuXtbelYaAnX3
KarK5F0UWI/6VdUktTtDcHnSOTxjjdyyaxf4q2VqyIYOMRD+cqA5ncFZx1w8Sm5RA9RbGin2ZVCV
s8RBXkRaq7q+/USMVVVun8fxFCSxPvHaoeLsBCShi6Pn603Y2nS1U67UcyB0idlP46JD5OTyfyYA
vlyyN08R4K+06yyAV7xfE6sPId2F9lU3q2+qUx0PJxOeFSaJ43hPTgFcEblA01R5gglyEwCdlAg5
2Zl6jaOYOwwqnm49OS7K7xc2ZLvz4Plam9prD6JYfhIVTtem9QF3FWqvgWajlueo+XVzo9RxYtam
7P9k3bBlPBQWinaryA4EOUCUalr06oKQotPaAvL0LKoHEL+h1Iribd48i98pIhGYBMtTZRBlHU62
7mabXrrw8XdhvY+j1cgp5kXVHLicHdOYqdBKceUI/RWxryYjLITLsuXpxFUrJL1aqs4M12yxlARt
QIQIIcOrQ+yx7ouovfgL7lkSrOTG8+ioE6HF+E/7gHOOMgrawUIG9PYfJrLu5PLd1dxNTAxxpCrE
HjLopFH0kezsBpX6X799DMdfWnahnvZ0Z9ggGXrVqioDbxiiTbghC9rKpngi0xPJNa2tL9kxWx+y
KsBeRA747n8bL8WnaBqNy8woY8e8pWHAOd9NldZxQRehj0E7hhXCOM3T4aaO2Xsl7UBSHLWYFi+5
EsEoE9ZH1cL5DfSWKGNV5TqQd3xc9cmbC6JgqWr6s2ap55UlJjtTu8cIgQ4Bl3hMXlxXbnKz+DWL
DilVVo79ANilJEnL5TlyBzfvjxwiRauhS5pnAGuXXapVMYqv95KscVUwmAU69UrtpvK9/YcoGFaL
8PFNmE5OXoX9ERGcaSBqFWHdF0YKZSJeZn5gi+ryc9fiorqC09b1h9R+Ene81fJyEI3mEphNbd/x
/EnEJWTrzxeiJg6C4ZchuY63iSkcoo7sLzW7ugY/6+2jNzDKFvQqy35XYbsgSuBtlev5ulNe0d8l
9MrYyO5wXR1L0S3uqtG6dO1r5j/9hz8QN9/4pxR9sK6WoPL97OeWXP8OrzyhQsTpBu2SsBVtzZs+
YiwcKdyYFr3PJoiyQo3NvCrFOGY00bozmpr9rcK5UgN7GkPkhvdgkFVztA7pindyr4OvpLnb4fPW
1CqhtccIU0jCwjEQsvw3JpT+MdhPQDTXGAeRxcHqoqQTE5moFasUTYCPCFuZhaZUlSmQqkOtxmoj
E2xmBEqPuIiXUEgq3yU8eOixXhpNhKFuG3cllj3iZZGdsrJq8Do7fXb9akVrPiuCCzQzJH5GWnH6
4633ngg3f7q82fVB0OBGEYGMaRe4nuD57HYutkfv+MJpL5jUbqzaGNr1ILIDDf30sdO/CMZt+Lq8
+vObzUp/fA+3Jh1LDnZeWmjjttfj1Needgg9y6SNtphA/EjkD64nGRP31NRozdbOfvuoyvV9uzyj
Te/M9seMCxdmnDMV6ZFYS+qg+/o9wQ+n/vr7vl0BwVgMzC56hlrN0/Hj4UQ51K01T4wVYTgyaGJv
6EvtSk89CaEPQZgKW8ZW/g2QGQP7RXtgxyhFiNOPVyaFtD2buwoSkH179107DFEaqhS0qaDQMm2d
pfmKpOUZNqpIGOwRx3UMiOJdeLiIXLEcaJddP8eDrza739jOB8RNnTW5JQ8P07maf1STsMdzRlxD
qtCMRHrWnSdWOWwYVLKzHEVVFzgfDZSljx4zfBlcs6aBLFVr76kXGVeYFdHXDSREoJjV2VEVXXcb
7g5h57Z2SPlS2RiewOtPLISGJ+AgBhI1p3J59rC0Y5rbZrc1WYjFx4zgFbwO1ZDWItrZM1pM3W4y
50KavAHtqRXQvLSSxGLy93r5hP+IqmF4P8dRrdCsCrP+Q9E4vf6hRO89YQxMH5otfo771W4heETu
xdAyvR49XDkfs698bOKZzbc6nG6auMDAdTxe3ecaaNGng79D15N45IlURUmhIl+rVxdD5l+6OuTY
LEgrhpyYH7kjzEVBl5vLGjieIJ/XtbzADipAVGgmQ3hogl6m9YRZgQMIEBREDYcytHnvM/bCV/BQ
K1LoVEbxw+JlKouU5EIzXqoy3ZSBLNlKxL+dvcyNMC0KF3qAFQSyQhn6j+H4HE45FJu2ZT+RDoL+
0p40O9YqNBgVMUvy/VRaYT4PBr0MNMiO1QCXEji1WHjevS4blDqA0l0+rwYjsofD3c+4R9IxzCrf
ip0ZdeANYgio/TAPOXr4+Yj2B6UxtIQCpG3BFpLfgaMd02N5cgzP7AVhF+KoDSQRUvf5sYcLpBi/
SdUT2KiD4Jd0JWCwM3lGLKFrObSjZCS4bz+zrc0pYXbh0fFd8xIHva8RY7LB52cD1VyJOZnsbwIY
69auYPwZjI4ah75UN+sheD2XPlW+PTrBHUQN33L0FpIQsYj10FrYx8CPfN22v/Wv5DmY2PZLHqbT
6pW1M9YzFKUNoWkkPCteTyjYK+8OOoTR6SWccnE2LPO8IAG1hmit3oI/oVuEoTVcF3u8zXnTn7Xr
IsEZVq8lG29kGl3enbngmtj0o0WqT8WI0VnXhAi1jyilrMz1j67xyAvczOoolFY5V86prv/MNFFc
DLaxAEFuIltd8jOzgWbNCI7BTTZMmaZpBbaxEt9MpqBsbICc0Cse6Kyv6LD5XWjqx5r1qKti28ik
Xj967WnKU9fPXlSSl/2k3pQg//QNZld/n2KwYIaB6fWFAE4lDTXhRi7OIL5hAW6NeRv6cQjmLtH9
KKdb2A0XmSfQrObbOGBsPIgCsfr+aJhRpoXCkB3VG9OKGy11NwhBuRE1zN3VWYV4B/t/LglfD4nS
aHCA3GUYBM7QsGlTAA8RzeEk1kaokqlS4AqFEMriVFjK9KELPR+PmwpdgyhLvWKyLXAYy6n9DlrN
uAubVT3iACOIPaetEhc4hu451+5FGNMkw1te+kXfXdZfJOBXgaNnPa936jp+m1G1Z5dQ1IBRdCSM
3kZJNLyHuCTBEgy7PgP4JPqKYptqjAZe2Pc5gv7Yh3aUXW8cESht7wWKe0eXeD4GwWBqBZXnVJPr
84oUeyG1MxS99XXu4ct1KmIR0tvL4VQseTpPAylEgCM2t7aSnAXU4KKZFq7wbFOaJ7J3Cr9x6E5+
kxPMs7tzu+CwPy3KifhGwv1gnOXezbWQ3+P24Uv5AaW4ykbtiJFAvWx9aIb5zHDQVnHr58oQwysc
a1qA+8BLawgCBLmR3JerFTKcJsDZ164u3PANIne5pwpsXY/O8oba/ZDVQgUebpTb0ppc2qwAiCfz
Oy/ynX81FX8xveW/lSQ7fK1gBXk0qxaHsKsz3PpqXDZDFhvwolX7FbKBuHXq0I6R0vUrxBXFLTxI
qe97R0NNRtTkERdQSIU/FsWdN+gF5abJI/Dv+qax3/SiM0xCdgdQzfDGzgL3GrRL2nqrB5cYL++J
M/vKaPlHrlHHDus/EmUFizzIeVdGkEja6dDL7F67dJMcoGFpDnB2IjRZJU0mLo4gq9iJXqFcZRha
XBIFI3gKQAaRntVuujvxJUDfNC++hNxlecyrzjfPc6GhWJYK5bMKiOOzBBlBVN3/YuZkkiw6TsbF
6u9+txEggXo2YCH2t3Iv2W5pGq3sdS/2+UPBAboTBhoCff42O52XeQzUtJ56zYtBHomlkT0b8Cw5
ZDoCDhQsWLf5t7VWwDlxDfaqF2p52o+8HJ0OfLgvgL2uJDloC71nxk4cbExfqJ0+lF7TVI8/B/7S
E0FdEF2ZnX2LRgh92LvM9d1/PMZ7+AwRncYo87/7wFvUyvCEZoiT99kChNcM8wtnlabUvrnsjQHQ
jdRQjLNvnGSJCGofQK2uaVQSW4FcI0BCTVRbOSDLuNaosfj3hopCgKBHGhixyiL1AHeGbuSP5EeE
+6YvyaWOTPpYfajjOJ2O+6L1TJbn6tuhG/B0zMlAXckJZ/Jn8c6yUYtdToImS7IlkrMRACeGIP+Y
a7IyWCtwjCPfEr1e8ZVd2+tSvyAqGDwZgVAAYqM9K1wTMt6Lv9NayKqzRMzh4os8yHiOCBOORYZY
yZb9PvB9qJtpaoir6l5fFYijwoofOs8t7vH6MeibXE/Hcg6h//Rk5gBSV0FXW86H/Bl559WXFjp8
nwR1WZ6nNGSRrVX2GKH7w7z4L5ZsYnL3pHmC1THxAI9SPP4Ljqja8OPn/sFy4AScEwlqnyJkNW5B
6rDeXE0N3PBk+a8VR7lroXjnoHiSOaugUXm0q6l5TMRQzDusQa1esBP1IssxIAt7KODxG0uATaOw
Q4v/9vfelfz3r1ynqFs7qlAx+95f+9ZCUiZH9UIQNZUgJ8cZuBBJWZmwTQFKHF5+GJrp+csqaXeQ
KTvqkQ9+AYJRZn1Z8tTAykiISZuLuRGQchg02FZniGYCr3gV3/rXQCO3TNJvK9OF4EPS5sAq1EQb
Aii169aRRo235HLUcyvMrSbMbcc1XfsC+3s+nAYUH5NBp2dy9m6t/BKF+nBikurYSUNNbuepQN6W
V+E4xhBOeLcjmO4GhQf/ox5uzrukZiZii5ENMCLFaThOVcOjZasJsfnXO1kJi+yadtKcmQUosXUX
Eejf9JQiTizeaEnW83TcS7sJZuCiARU3ldty9B2ZBuLgZbEen1tbEMSDuL3CMWHgnEmIppQPr5GY
rDunAilMY7+GBlw4HCmG2MxovqanWdoe7sciHlE91VA3SvYvTooFhzeM607cQ2yti/fNSjGK/JWU
Qq960pIoOmcja8jwtPwpTN7QeF+4JcZt1liR23LRE9Rg4yQHjS31lUd4x6g1HJkKmdazrZfhOc4D
kduqACAkLSV2GCoUDBanZUQ+tR30WHTT7KKrFJJM3ioNT4wjdK3vgFismscr06JvZDSOGcHhZd9l
NiwkY1suUU3zwIeSuzVJKTytmvw+HvA36baCa1tz+/WE0vQ0mLZ0Al3D8vuQLAvukR4Yp84pNker
H8aryIDVFC6YFgz7piDPh57w0TE/ZA6OuZ8uD1NV7zUas5LcASVzkb/oirsFAT8ACDm8HjE9kss7
QhGx8UPcQTLjbAAEuIbvf1QXKai6QBybGKFS/rPY83LT0u8jLe6cQFtwPcaX/AriXf6DjSOIs5iR
GMedTTjhrW8QkVTuystgrIl3qk1T3S2nRLX4fIHAely/4uyMqfOKikRTo8Gcq0H976U3HS7Fg4z7
vYjByFN7oZsAq0zLvDlFZ4XESfNT2Q6CYntXcvQMn6pk8d4nQmV+8TXy8NTswn2FmusrXat9xbKf
vNjAxw4/vgFPRadnUzBfVcDJEl8NoSLQLg83DlLGMf9byLpk4YGO0+I4qzkgDuZIxDsYjNq1V0f8
nULPi/QijXkGIr6S44mMTevBxcR7Y0SE/4RhK0LJ0P53X4/EWXX8JdMIJ2j9RWyR6w+vg3ZqCzGR
TxGyI7Zj5Y7/0HrW6R8Kzzn2UoH3IpTCmgnaRb3QoHvKmZe0Ntt/nSxatzXrQ0pDy+GTFReIN8EJ
USpc1EWGUS1kyeV/RVRsbBztCQlC4caP1lXXQfHtrgIcnOOj6/B+SlavcilO43TmFOv5ILbwoank
no41OP7VWFda8u2haRC5ySbGsiTh8rs8R7xQHVHOy/lE+1FfL9CYqbHTgpOpT8uLGpF1CCaSwG3X
hr1ZBrVbb56CCFegiZ8pOssMq4NYB8jfpHjVsYuvJSu2e31LHLeW2/tayQ9VWWuWgQoA6oDjks49
x/EXWwhWkrrAVghNCpDH/dlRD4KvrarqNocLg6eENa1+cjBI6NcXMrrX/m0A2xIIoZ9vwjSFt07G
55RSM1iOUrhycQMg4K1ICUCBPN7MYC3wGZ4O+ZiPwRYhNLv0KgzNsciksqnSFsNQBBfXjMGj5dXK
4um10N/DSVvVtX7dxLXpl4iC04vaOVoPUD2OinNsM1CrF/qoNKKynq824K3T6I9Al/M4lvDxOQke
n9gpqWltCvVgeN5QNFYl6QYlSAlMMCBeAlvZ+iZejcrbzEHAz/A1cGWsysTsJTcs6xUOIaN+Gxbs
ICo7HcP2LTTA21j+For+zfhtLsOHVLaQKdP2Bzp4pj4Zcz9pe2qMY0T84kEnxw7mv/+Qa0Qub/GH
s29BXY307ZkZdC1Nsc425gwYdFxLzTlfU/D45Qru+S4KSow5bmMef3lZv+XXFrBUqbjOMpHm2R5t
ovdMjbf69b744GltEi5BodlmgPCWSGOoefJbnAtdomraN6seMuwDWwzeXGic5rPP/h3BE7XO9pK0
vz1aJxZOs5WAR4ZdDxgxwZiZTkjXhS2DJGUNKAfzdBN0y/pWnRVAXzKjEnk2l2LYSOjjKyz/XdMg
X+VMCPcOO+w4fPjaERZWT3XdKK7O9yPRiiDi+PO8hMh4XYijxnKApBFo1BcUNcOJrLE3im1kLDQm
XBPp3BJUplO69NTZ6dngH+mclLUA/qJS+NuX20vOUyQHrEkIkeMBTqRzdUOB3zrJZ2Ue8EQSlMP2
217+eixhCwqZ1dxY4j5N6ntZ3Ik2yPZwGNjNpkN0iRr2iReftXxdXbrRSkpgUKK+tzNmVx/C9dEm
Mn/PyarE7gXX6sCEhsC+lIitj84zUo84uYSsfSPaMkZoVgN++I71fynKQWH8cfRHI0BOmexUIegn
b+bKn53B29Y1YkgDe5ZCx/9ZDInxpQfKtb5AK5oSljDDtWkjXAJDNCtEebCKnWmSaw8Elror2vW8
Hn44gcn62Rz0CSZZu3YEe+DwcWYZxm7vGo8q2yfG+ImWUMGrHRmp2GxrwJSUmPeODPHjNxFzw62/
UyTxtMBC+6ley28lKPZAdOjPPOs9J5Bcf39fVlIjwtd2SIz4QE/iwwsLVk3uvBZx1FEBq9dQnH+Z
s+RRCwP9YTm332FaQouoqPnpl6xTOqsSEB7zaRCaRNkxKzwtmnNrR/PWsvZC1pjDYz5Mt5qClqeX
PLcVXN8vOcmjJ0c3Xc7QuRJRIZZTDgttK6YfugKlZv2tCwdJSUZL6asns+TJfPggjvxJ8fshI0P9
CuHAhSb06SRI1X03tpJVweuEG7qMmM14ZzX3LsiRm7hFjihoKGZsF2F44Am1aWKTYZ9x0KUUOl19
rib/l/kS+j/M8Q5PFGRjbSmTYKDZs38+epZ/ntNaJa+cLEaA3tpx05q36+s7yVVnrY75dyVxl5bO
Nr7Vf2rKZBIgCMZ8V2AXhF8WtnNEFYov9wZ7mv4T1MHHA76B1wnpKNM7BRJuLq1pom3KSUHuWq4A
T3XtaN9e/x4qfYv4av050yhFQ9vFktbRxL7/pqWnTvc7JgZyCSzqJQMdrTi6BDCt9W0yTZjQUmza
+EVz+fCZ5NmyPbu9WsY/C34n5uQ70GTVwTrxR30Sx16fIZ0HqoKKusAp6S7x7MyJbXic8CJ//Rlw
oPD557E8L5ffFEHAqkLlxPhqfoUXZERFv3EGv3zcT2TdCQdolHq/goqkgZ3J5fLYnZtrQ1idj23f
8SkyrqJH7ygNcNzMeoaC2jMZLUxAuR8jBAgh/IYvlz30B8v/b+xP0omExfrUaoC8P4xk6Q9hPf5X
wYNITQZNxXJmgKvM1GQFLLKbtO04fagKDRQgT+2yN/ZhKY7dXZAz/nLWvrQqdHlUjAqeFbhIj6WT
EK+4Y3WWjQAMo2UyLGV1m9r77514xqC3fp/8BTs0iF8dezD+GCRBb7bVDC+OOgIrNTB3Y22HZcu1
9U1oM/Jy95qqA6rebi/dClQJEbYX/DgzZS/rWW5+fvM+HgFHRQQRmu7crc875MO0zCLlG++sIYUo
lYbGnhO4FQnW4ixZZ/2JNBhrRO9GxN4hkVmEvYICcVqwhWVIh/XJI/IO+UIzlFjPjhVP0tsCRSB6
inkYZ4Ef2JRdlxQU6JwS3RQXcIRyePYbxLaXJZaMFij0j0NoDfuZ8O5aZsE4Vyqu3UnVsCDQPC7o
gM1KafL0EZKi90UG+ohbfzgpLAFf7IRWAzYXqlU/fdPQuODe1FwSoLAmrrOkbpMoUyFgp3hk46zZ
iZmHsrXoejDNX+Viq0aytPHdYkh+cXq5nDTTK2w4pUqPStk6m66JXtU9huM2h96dV8a9j+cT4C9H
lcMJ2a54FuvLxJ0TGj0tWVdBDzOrvOLy6oeq9NBVbyHzVRKLQmvLJCS0RTgTX7fGlR3y/C2OQMDf
7O0/fbhDiYxCUsQrB0AMEGyJOAblNiEZEoYGYu1Pkoaw/5jhmPm241q55t5206IOB/w5TT5q6i4f
qnoqR2WQMbbyA3DTE47VheeBCBu+2fW/VJZn2iTr4oFMg86j+/U2APzIgdSpdYc3xlJBeViEfvGe
kIfoW+qnaFkefzP2Djo6Zazst74z3p9/4OxVHkszU44wnrU7DxijoozzNLpKurtO0I8LrMGgT2eS
f1dFssyC3yul0y0fc3YibPvHREY6qEQb36NzY5KPH/5/p63/1wihOodkFA+3pq/vjjIQB7oKSzzU
j1zZ35Yg5ZvX0CzmJQLXqmASoJ5EbZvfHtFOP6ma1/z47AdacobKJNv/jAEOdL/Ar+ByTGdgHNIQ
gJHWMTQHp15LL0RUMxsYVc8poP39elJNeisjLZ/+JL4SZAl8VD16SBUp0O9CROQZFpGIJaeego70
yn7MYQMSXYZiXyNlaNW1SDrPn7XBlJShxCU6QED1FBMhLKhtOKC10STEXAMI70smLBE11sSyZiBz
a5Yq+KItqqBM3XvbjmSUfzFgwBGp2InJGz4mZqZGUinnT8EZHckLa5U3GKYoCcGiBNhBVG+cyIB7
+68h/B44IPnIYmIdqQQRh+Pc49tCLLlNsc08E99X0Fz+fBJ2ijlalrTgIlAhBEYMLuOy2geWM1Te
AcsXJ7TiJ7erP9b1HVDJcR1ZQksZES5Z9aNxlsIfn3FvNWtsfAQYAdnkuMfNWDi1dwcgF3C2D/Ti
uh00v0MYI250HTiwLIzoHQcashwXQx4jkftyWPad8bZKrCluuArlS1evAn2HDxU4RZ+AQjYF8JV5
70T0mzt0EmBPNxye01z6OKAwydQ217RBjm0D1LR66jmnTGT1jTToDYq0yYKoioBPAV/4kUuixoe3
NqbaGJT1FztwmAgQXdcHXPrLaTD5RScczNu/ifa7Rq9P0I1PaJSMrNPrqHZcCqc8yXN9cTj8GKAy
v47JdadtmxzR0g89gWNLbNYKWOrC4j0YkD3J1aRJvP642/RL9yvMB74tDbbHSER3tP31KdQgCIa+
pau73f99QvQXDvmh7SUeV/dXbQVNGmA8zbQS0ZCpwLrMxNHNFj23sC1tKTv7LIdy8WNzHvAAp8qY
U3RZ6vY+tk7XxEl3cVtaR86n4vyOMN+NCDvinsGNEuIHa8gPCTjj8FrjaUL0xxyxtnrOMmYih1/a
CU3JL+0fJDs7jBwAjNHuc4oILScLwEoHBk992SJ4yhtNrPBs99slmMAlGKDCstizfen1a/QFcHL+
jfzF5cV66u80iNKjJ66oeR1n+wxsNblpkER2FqWd85FIMJq75xx9wwNQXIOGrq1fahlstgYUKqHY
Y14vA/zaU9ZSADO657p7WRRX0I9C2XjvLucEe/eXuH1swl1A/Z8foeOfWA/IHWeLPiujSfShaWPJ
KH52Mz3uSw2KEvYZ2hz+Aqjw4Gu1bT+ubMPqd3PoJ9Y63j5EF0exi+Z3YlB6gHqb8vwn4nGENUJ1
Qte02LS9ifSuT2ycFyrKoCqVuwcUTWbnFnBBH7mKbO0pJ78SyiU2Oh0pcZW7/H/q7YpNcjgR/Zp2
MH4Nf6/OOt/BsZEP5VgOEnrIpepUjVKRlutDAv0Pvw1WWsvY07qFpz+Jb5UFBGzITVufn+r8tfA7
zYmqARUubzl/ROzee/Ep9zfcBA16lzDk9mrMiXibwW1nDed7d8eXOP2Zx1orAtI7qJHr+zBmmBa3
FELeFbOaMBtZJJavulBtocLIJYloNQyYTQmJSwObkiPK7rgf/RieuFvuIkpR1+qRl16/W9lgFc+p
yEG6MfFE7uVuKRpkyGn0LeE0cc5azPzIjxEKKlW3K71Cko12DkzNYaZtf8k6x9z1gERm3aE2ybKG
7PYcOtLGo5reuGsr8nztYPSSbqLtVwgX+Wf4YIjWRYTYqBvn9z/o2iAEyVz6R33yCQdj9Q3oGSJ9
GcbyqCHj6Sg6+gus6MqiUzteAT3NYhQ6lfsvkW4nj0Gp9FGpKG4LIkbOYoJhib4oPa+HMLrVMUbn
Xt7XAiANvQSXFzrCE/p8WXmrQYIPLkqNf473ly0q1eklJry05yOPjuB3Rj/xyQYtd3MAighuOalM
LrvhmDvHayPpTlVoDsolSIFpKeNVZ7ecw/HFBYCbBsz0zFl7TQRfa7f6n51QClrfhVsJO2w601FS
mWlUoXTQtNbqHx7Yr/igOqCCV34fIFWYHkUV0QTuMUgJxFO4vth0Pfxb9fMGMQ5U4EbeGHH1VoxX
lkVOkblZyj5u0/ECgnoRqezmQ5NBee90sc/zyaCNRRjlhqnbWAQNTtLoRNVilk+n3+8BxQMUDQIo
lZpI/sfUADTimNRI+qgHpwUxunhk6kAKTw/l4nKQDUrEFYaGlqEvNfSBKzZxFosVk8SHukWdOyIH
gJbWsOtK4cKxNVjvI8jkeja10DAi+Do1CrrADA2oeM6qhJbLVKA4hCFOybYdhOfZfd+0RjpdW9lB
gTHJpQqNsX65AiIHgWQ+sQ87qqq7WP5LlXczV4hrD4gsbzxscZTS7ScLeb4hZmD1WC6NMdV0Elj2
1WrZIl6p3I4sB7Gm+tbZFrz3/E3IbkfmNRspFghRki1d0dl2dkFLZAMdNeeJP3sqDkJRtT8oCUBw
A6imIbiU3xCiG7dSYVF3kxCqBHM/3LdgiVUmaaG9WW47hwnCRyaWwYr5ai3vne4Y7K0j0sAlVNYt
GNHUH78SbW9TpJjAIIgOA+uROEg62SsvAwLMPzz0TuW/cNJBxpmjCwtV/aQRbYNvk9tbDPPut/jT
V7KmuxIhm3Jci6eX3uPJp9p/DkCXAVtgxPcjC5lGml/dwLLEPIwHuXa06OWc6qn8dGbHonkpxy2P
HMNHFk9QJaY6diLu021gXTlz8czWcv8veaaYaGf/FyA+UMo4h/T83PahTAPA6+j2wCX8b/uwbf+r
lxxdKTUqaCbhTkbjXMrU+xO7SAKNDL9ctHiioVvTYvClxVjmpdfEBKpjvjJXlime459QnZ1QYTad
qiLRXeN2Sr2OqWRwPbhcsmMv9R0y9wMp47cxV1KOfd5r/eDHp+leTiIbsSMT1O+SsnHU9h2zAsBW
sWE+PpsHY/e9ZROy4oWH0jEYvcpf8NMdbL7BayO3nFByx57RDzldbhsf4ghSQYuPbHj7bK5cKpE0
bmMNo9YZ7ZuI1c1X5aWSyvf7/E9tyoA0jHLOE2ztsbzrZyts3sIurVFu0P7nDuCT5oK8HaWRd06O
YtA8nrHldyxTYzDmE4zsQIrFjyKZApEDRqdEnad5ynQQAYIJPpeJN9aEvu/O/X3VPtZR/tCphtgA
A/w1b3vRzHdpCaDD4nlBYVqgsWo/u2bTEcm0QZxZPAjD+hQbCDlKRLjvKylu0XcTMgfN9f067jHZ
BFzZxcAjHJuI8HPBzh+GYY5zuobfvif6Soki+0Wv+0Gz34C6i3+FQBtH6ThybbzZWRRclOVmCHuP
biGBhiIeat1ZnBttc/6/WE3sCacEYuqsi/JmZBcO07PFuDZmx0Bxn3y86b1Zr5gLLHnDLZhGxg9O
XDIdxEA4pnS8dzXJi4k4gDIbPB1x1ginqLUSQ7ptlmSrQjiACb4ITnxe36Yt1/D8VIbCsY43V+TQ
TvCZcXrJRK+wmbRLCJ/ThMo9yR9rou863DjCihVCq4sZC2T6pXQq88KCe09xOyalqcHCttjIEECa
kSBIEZZLOQA15EP3bW5RzawgH0epln921PF+7iIPcbA4JAv8PW0oYCn53A8grhsd7gRMA53C2RF0
/NW/i0Dq/CDCYC8LSpaCNC5+mSkO7iWsREJ4xiyjq41JdseNrxcffQSkj1SYaOS0NKftA2HoT0VN
YafkBD+8J91Yj4UhnusjFn7h2jZhBhvTbAy8VsBu+VsTHUy1mYD1AyHf/pvBsd3vQIgzMGSlwFXx
SQM06M4xBVxlDbPgSayKcG0PH5J9wP9zZ7AsuUuahoCBo3ZNAYD9SHu82EVDdo+c1IizKY48rDu3
yaXznwq+jd4ykCd7pcpoVB2SVAFKBX7kCN0AGCpp2d27knZVM4N7T9p+EH6hD+9EbcnmrExVsl6c
b2xOG+l4gsOqLSmoTgafZ2/MhAOtq3sjowWCSSjwByc7bdWnkWgLuMkeZOw+m6MzDzpL9T3YuNFW
Tf1Ia0yb5IG13A34vTpkdjVjkk7iCKbsI0VugV11FfvR4SVvHUxH1ahVrC+7UQ2woA1w0cdQPsKI
TONdnkCKT0xGHRTt3iSFwxhMG5Ul9MTzM6Hk++ZGYmtA6R/9HX4LHXWNs0t98r4QiQus8pT3Y/Nb
NHWrxlTknYPKY9XBnHREuoIH/IIitzO/t3LCxeJY+pZKPAyYegXjcjStpTsbVyqRak29uHy1lKwU
FAoEE2U3FQgVmsI3wNCxZx4VyZBETL00bIvn/YoWrnaj3mzISWcIqAGKyXF3Dy3KL83J8V+J3hrH
DBAayuHkRh1ZAicgZoSF4vYVzdGn+AacAEwTqjEyre/kt/tTJ90AHHLoW5kAKlBfB7E0TukQzifa
0MTLQNfmHCuXveR/p/vgT47jY42YXDuvNadEITFJ+uDYqK2HA7r8sA4sRdhNyMohKhlD6Lkw/T14
AMid9Gt16AGSdHhNsRNs04DqJ1Oz1OO1UwS31bG6fSS9RFDkB88u4QrDVJsQay8QmqO0vs29f6Jk
d9IkjM/jdhkfcr/Lk8V6dDTso2+lDULBuO6021hwEbX+dFq5/sv4wwjCl1MimSFgLyfoKzUIUt/P
6md/fuotVxiFuUdawUy8wTuqCzenloX/52uxx6qoHptccda7S6SgudWkgTyRpeJ/2NE2p3pa8ycY
VHVAEy0YEKg8p8brC7KySSaHLGSGPqT714D7QzFz4VDLKCcw5s37q2DFeN00mx7DvbCvwGnRwZEZ
etuKfh+2rcGeSmweXj2xi8jPmy5It3SYjWZDJCoeiwiIDwjF04RBJsdshU+VGfIYg3t/tndXsq2u
JR0N05cbFJRuYDR3XI+JiGFSPaWF7SOcFWcJrl1z11gn4egtulVupg/6fbgtCfQu91oPdxOxPW0V
9GyLo5R5RkaLUl1kXzyFZJxvYwYkUJ6rkBqrB3ukhffzFmXpgbma5gNWCxhY/ir9tpDDEuKl5+tH
rZnZomD055ftYrDIlP9VPsUEwPuRFktUMTptV02sZohBTWDRJU53TwFdJ/9UakFe1MJzdwt3EcIM
hDymZmt+y9/WeaSRsI1IWpIz5dRQan7Mmh135CSSEzt2+qHX2s8+HHZG4btrdzon6kfDoBu/qNpN
Q+bPU3VLfKs8l7XuJsEaq6Hlmh59cCDLcwV8fS1uLSbGt6wHNL26Usa1w6tOaEbbFydWyoaAVRT6
rtpJBJW8jYaP0i6Y/zwHjfJvia5PUoaVzIa1YhGEYjKmmQYVGcnH9tRAYI+vahO0UJMZXq5+gA30
Q2dJKDhvNS/4gb/dzzr10Lhem+0C0AdmYEaZz4RvSCuvwZ1J2N9gYTJ+7VNx7HEmaAoemo8GDBh4
NrZXo4rZFbOB3HvQuLlwnnxl/MDmQ59zard3/TJsLYdOxJ7RTRkmLoHFQzfFQVX3eaFpJwQhG27V
y9zDihrOwjj8HJreTbYAd1+EyfN8TUZIT49mfA7i27bpqmYEz6kqldUmlaxAjMcBjKn5zeOja40U
PnRieC/PLNh63G/2RWLnFFPUtJYl7KaIvluwlCBQ90LuVjD2NT87SA+9x1aTsPLkeYXsJdCvULK5
I/EVnysXzE71n76+2BgsaZKTq20x3LjaK/LC0QREOG76vEWKCCxIUX0kg7MIpKr7wAaVVmHzu9PD
oVYdCvE6RhUZoR9P2Szk/vMlmPAOb3SFj93osS6OXC3G/sgXMivaTeX24GuboQwufrTuZ6BQ4Lny
Y+oFGSpR9AyWNkL8jga2bolo82pH0C8sbLnc9uNS1s3k1SiUy4224dPtuhC03ea5upa1HNRMtkCL
u8rQa/7PuSSfrmqlYgbFp9FQPzMxeY8YNPOcsHIDDQl4quUns7HQdnrXfHxxs+rkORU12s7Aa9PD
byGnAvhGPxriFQVEuID52ic6N+q0Os2jfYQnX6XYwBLpe1wbiNcEfdAHt3mtIRinPw7oQ9F3l134
4nTdok04TAy/qkuX16KoQ54+PDAuTB8buFb7JIthtNfdPAg/jWlNTCRsfmu8k/gHe5HHhDyugnCC
4lfakKmafPoU0VBNt8G78J98GFzJLXWeHkApVKtKqfs2PINX/+7s+HH+Lvxii9P9taTbbWaeVuuP
KbsDsZzJ2mvkhoBdhqJcxLy/v3zJzbKlBBYFoAl31LdhmOuTkjB6kmDgP4Nk+4g4T5FqgMaaoaNV
5zfWCkWTsndgSJrY3NfQXQeu5SRF5Xz/kMqkUACUCqomJrIx/pCSRdvifMha0ElultdMPqRXLyCe
ZZffRahCT9Tt/gQ4/2bjqHzdIdK/xO3lXQMAYX00oe0aYnJ5Wr3bMCm+b5g9bae1dlooiI9Mqhrh
hVWp98ykaknfXnhxsyGduCFah75LU0IGVjQjWo32vB07OxqS5yn9zn4iXM+jfmbe+cw2+NvTr95U
kekjN6jCeJVLSgbBAalexfYI7xcJFA3qEMOVnkSa+UdzNPJrcG1Gixvy3Dra7Q6PtIJCArtBYuKj
ZMkL31O6aHmdgnozcY7US7Rx/swwPtlmoJi21a2ys1+wHMgwEvaqdBhXS+6xZnS3tX6unWiNN82g
7I8gY7HtAaWN8NU/hgcxKDtg6NU5kh0wxOfMH3aj+mq6DIiEY9W9GbwjNU+UviVBWTbrltRF/WXY
3FGfmi7S8oVuisTGAwgo+U8q9YuGvMK18abbDC1UH4EiK+7qDWHmU7XQ0bL6P354fU/Eh6bLNbtC
md0I4Nj9MtWHhQP88ikdaFYcKLNv85S+f5P/PQgZ6vZfdYudsq+oYt3vQlZl3wa7mdSr0wniJ9Ps
UcbNuk6bEs89GQve81yZbvngZrg2Ics2c+rbn31E3Ad9TVQ8WQU8QEA3uL+O9vBGJgZ7bF4jb8cT
4Dfh4veYE0GZVBCyBYKvllXSxPf/zC5LKPUcAZIqxS0izr00Qx5xLWPCak4/LPhwCxILmuf8isTo
la33xG/+cuhMHMCTz7B0hTuj2DSBdZeSuR2t7bE21RHQcGMPH4lUHy8jkAX429DaT895/j3d3wRj
mC8ctzrJTQcfbFEZZYqti81wviRJ+yeWfKYQw+ZUACK7et+cbyT6zFsKziVcU8mZqWYhM3krQPjX
ifa07uQmDMqX6OxLa3g/P2IqqdRURDYvsk7YSYuTcqtl4mv4hNuziLBvKp1MgxRGFbTrB4gU9w+V
SLbRE2HAvLtANiuxmkCsZ1Pi5T6saLoFzaMwRVHupBw5HGDvy72IiP7s3roqElBwWujDuzg8+VKt
RKEpuPQlc9CDoYohb2GY2q1GHvGfcwCh2M2B7d3tsmjgWiYtbyk5YSGyIQeXxMjNqCFgImcBN4F9
YCgxxmZAMBG8Eb1XCQPxuj1ZIxI07kRfOM94BX3sVELVao6VlJ2dqp+vBCpuI+LU+axW8xfTNQgI
4ADxNBcxOm/My4FrquejxPJbD6+EMt8Vlm1A/BvnYQqyGF09KM39Nwb+0LFC+8vdJkwUakB89Xdt
7e4VrFXowyqGMtjx6D7PY7RjQ1vkZ9i0+WuukJm9eFeX7Y14HOGrp3He5+BeY97f2JJHYCtBK6OZ
wunFHPmFf6WuuBPVG1YhL3wv/cISdW4VK41lVldSY1sDDma9jGS/Rn4etPZYcksCVOvRXToUApqf
5dfGByh7r7M+nZb3NcbwDBbizRdEjcDyOMLFp4SX84MMrE3BeD49Oj+yb650kt5PItAonsv/9dtr
1ykuz7Oc5m2sdWe01fOo9mmsK6vYrqbTbTH39eJlEIoBSWx/uIy13Xtt6thkP4b/QX6ka2kbEmJ8
3nzkQbJmAAx6jbgdb32UuowymHqly8y4eFa2BMtaw+SSpXmuzXDsd71eFiBYvhVyJdOTnFdtWEbU
JqRwv0+CEY9gdfbFrEFPVACl1lwQUhcnbeAsQHnOd0fL1EwLaOJk5sZ/ODIkWyRQhVYDkKxIbXJb
pnmOQr9FleVaZ+YvE7x8h4Z3XDQe9k2Tk/1wcaBfw0Qf4XWsU8u5VJb8Yfk0W9K9ZG6es4AFUkzt
pT0FcAU+tHv4J8Tz/unpfM2hOerNUsfoCXzXHRoHgnAx+bhp/peGNjpxCuaE3iufqIp1T/GI+81X
1Anyb8+GxHKup9cOONw40pY4PDhm8DH3g5+YqB5VBDg2rNeZ2oYg+mv14bi/3tXC17sryfOWXCpY
WUuzJijBjSzwkoVebJQxOm57fCi7DG0QGTDFjgXJRwjKbvKdzB5DOnI4zcVYhO9pd45rcXjEvJlz
Q7HBMfee7cNUWS82c6FlVqWcWcC5I8Se9AAmHBRY6RXR88Vc856RkyYYY+hoYmxYI7QonuSJgJQa
xKb6x5VCD8r7FvSgFPVDJgMeWNPg23FZi98xOtcFAuV7uRCVx8kajg7U5H07IjBc93cP9qY2LknS
5zuj/kNcLpSmZxujS/AWFR0CYqsYoxuqla0qg/QRJBjZ8spfOfUkoNH4dF3H31GgTy5jf0p+xjb3
CgP3eKtsi7ajas9021VRXe7x5yvHjdf898aTb/lR53B6Zh2BquacXDAJeKSWUbSEwzqvBVHY7Fkt
e96nqyqsiqzxKR/TO4pdN33eBJEfVD39vphDmjrvJ97vR+zRrMfAqjPiSN7DGOHG/v0Txdqn99Ow
hIphJocLZkP+u0xcgPdZVG5dRnR5NRZ4UexhqQkyCaZfrF5Q+Q6TyVR77Fxdfj3aVNgXMGvu//Vq
xVe4ZCvEnjCKw2Kx3wYAA8XurA1AjAi0hMIlyNfFswmeTseoj1YZMIb93KZoDB0v2780w+uKrKgj
J6p+1/68U/nSzSzIVddiY3iHOOJty/XZZvWPXv15fFMa+uEr69cBaGyAJpwntk1b8U8DVbIrQb+G
Jy+7MgjspjiBz4K2ZoBsShOS1SO/TjXlgsuG9px+JIGtj3M6Hg6IX2S3TTChqKDsKOn3kX/LalGe
FDhfWlU0ouiB7PiC1Uue50aIuMtFV8f6sf3b0MPViM5EU94TVCWdrWTQB8ujAdVzY/DlH/NTJM3i
r2F8BF/DAcQIA9GJGNenc/AjYaxxLBh01zQgOSiqjaWJoNI/cLtFKr17TTw+52EQ6R4j4xHG6+MY
tZaTN4FGeMm4XK43WucUtEYF5kBCsn/lJw8LJbPDf97cfU6JTAefWwMBMtbEkEfi5EphFdtNtjmJ
nJA1ng6AuzdLySq2tYsQRGxDAl7wihZPiyYQ6udysH9mNp3X+4Yp1ETlWjfGoJpYL7KZEIxKgWHq
xVs9wb/4BBI4sl0iD3apsaJ6/Umpel+novt3I3jCXqofa9PszcZ1Jd166pEGhyhE0HqRTaNELY78
UWFQUHjsUqq6ow2Z+/zVePXeG5nCY32a6N3BkNC3ThQFhJ2MK/BIIGO31bNUW2FO3+Ue8zLsb0ml
m08xqnmt1+zkS2kkUNJWpLhJ+jxQKNWDpPP82Uyxw01XNMviN5/DW6l2OSAW/xWKWr1B/V85Nig0
P67yFYd863gBf276tWdM4LVqU0CV4Dca/rrv0hUrMhglS5poe0BTqQ4SHlKDp91JxS++F67N+g0a
RQu9axbRovbBM/IFZs3Em2+rBeJl+5DC4w4RVzjt+o+MkZUfS92zVYAVdz3pXH9ZRgUiYoUERzz7
ILgUtGyfJncnZ1Whg4gfb0NaJw1gkAmP1UZE78eLpFeDzGwj16s49iBl2LK+63QjtGOzYTKPL7uy
WQ8qKGGFfMGz9CEwfBcnWAeQzHHNe4x3rrvQmwGZHI0/RS5Fw6wpDakuubOHlpcPfRSYOuJrr3LE
QpL0Jl+OXNRsMcjYkWFGdIV5vAeWMAV7VLFzEivV/KJHlBYz/8JnXhhmaTodD7JcrLuoKD7FHcKs
JtAgkimQTc/4ftt8RfRmx5IhfwuoYZQXKjm9/qkIyAt6LjzFI997dFKSlVS00fLHlrtltrV7is7+
UKly3H1bF+Spmm9jROa537A/gVNnzuNoJRXGDRQksva5Yn2wL//VLDNlB6XdmX3/Q3+1nuBmMuhk
LtYO1Rf7iNfdjsRZOhaNSaYPwCsO7/zEqJKGHb5ZoF5dEcjJoojXNTm1tw9sogrQYDHSHFcsM3iu
i8UD+GVeej0fa7qIBdBzmiZvvKLeKXRl/+UZhp1ISZzwvgl33IA7fMTA5FmE+KpLUS5KJhp/cSBw
VDyid1GPomdxV7xVk6KIe9IPsjyJWlp39Xd+Ix1xenESQrssPVhHOuuoTS7+zmHgT7mnsSXDtil7
MECqTwlHM5LZHJNg2fQ1rYp3NbphgjTYtI3094me8qCTrf3cDnkiI+kt+PTf6NfOOY3FtalsOa9D
OXAXqfs6KcxHaBH110TfRYxlCB6O07yg74gkxdgctgq5Sbtd7r+O76nN+kxCRxayq0ObPn3mjhfV
LvZe1nJsCjIc2kExahgIbiTLxnANpDvYpgJ14Ot/jg8lPY4mYk3ZoM/buyGxDAbNnaOXIx6OW3IO
v6TfCrwGunr0GxwfbgzwjZNQi0XmjNdw6eiOvHE1XL7Jz8hoo5gHyuBP0cN14le/73W9+w2FPXZS
SnyBl79q21IAAPIhHUEkwVjaFsDU3WgiqNjbUuaIITckB1BWdg0aWt41HM99Hjo/lHXdz9J6s2WC
A5M0qQ+XMdojK43/cq1puwXMGgqNu5AoggTW0jS5fkyAM9BrpRbikqEI0rZXs32WmdkMLNAkW+mN
l+L90RAsd2FE9rhyQJAds4TxIyF4rB+fxW3jQhOIpUAAyomOiICd+qZSZgeBLY9qIECNEGR1+c+N
uT1B0LvaEJWavQRAZye4YGfK7et4nmsZ/cWEcTVtDK/l91CoxQbL963SN2RdRYbVEOjyZfjnXeBx
+Uk/IXhhjKc7g7ZKRzQqiMsJxj5E0+CQhff582SwpL25ZYZdKudKC3jRBZMfeCEZ2w7XPkYyqqpq
rvOhJKSj0W/Wtg9FSOAYhcVoiSjdEPdJKSWiFNud1Qt10oCGW9QZvyovPDU0Pg3+NaYKUyhexg70
Dkp9TLzra6x2BD2ewrB06PezQ6FsgZOOTlUoPrQynoVpJtRWDyntjjP2C9VBt21RF3bKyJsOmqAI
nwY1FpyAuq/rfm9C3dsWE8X5ZLHBPPw1dXZWwfr+K5FgY9Uq0vui1ZgWKbeZa8lC/euzpVKVXGee
jIaTBjTzBQQDEK1uEmTMnki/A6sdLZDXF+S7WSDNvn3IyckNIdGvPoX12jpDZCxqC6OCAfGwpUr8
N/uLVwLDIMMDlm+zHD2U99drgGuIPtoAjbAPfkdc/q31T8GHdOsFvCE30NHSVXzWRQD11XgrcCUr
y848CiGy/42AlIm+wuI8CxPwz4Dkp+xOj7z29tLZBvcvOJr3oeYvUvxEj9JICWkhmDFwoyQY2xoM
qkz8gKYRgAy3xSCOLzqIaQL/glH0TZA6V0sJbSyfOfyuNNyms+1fa3ZrdR8wydP1Vk5rV8Sq9lS1
+UxeHD7tmWVWv9TU0D1n58f+WiZ0FMf3+LbFwQHLuBTnATCGu8mM4wyeIuVMmwvAh3ctDydBd8Qa
GNDSvqJHJtDTu4jILHktQXv/1w+fkSFkSWXwHvJ7nCThAg+nxA+R94nzw/3+2xhJqgRZWWEPmk5l
eZWEjHBYrAZqKQ4wuWNLRzS/+pNHRk3nE1ICCXTMPpCnkx2IaGpUZsfknFxYrr1ySrqZIlzi4v46
0XI0uGsWrWJoOtZvXXSw11xlN8EOqnNpHwImX2CuQdFyBItHuy4ZczzoZePaQfuLTNfWQoYWifZs
o8oDHAc8XYBfx0VDU3lUmWjgKYSrvOPKzxl/Wov4/o4PZwJxgPPQOJNBjwSKeJk8Smw2GagDld1e
wgvwq6ZHT9Fc9UoUqDrnIBe5sD2jLygBKTHjPKF3fkg7mOUeI0N3paZd1kCc+42wVqiB2kWGVddw
LfcVCtcTC/EwKxYjAV2qkRVJqfJMMDy+1U2J0w+DEw4Jje/FbMSc795CDirV+3vzrC+vgQZ/ctCO
3jrP4shBcnHxKjp5I8sChuwq7EdIBTXvyHxv9+avL3VGwR1Y2lmS2xCpN5T9cooANDPkAfYPfKMY
fIQmHQQF9bp4jWH7vMCyY7b/J7hbQ2dkIaZvtUQ0eeE4J2olu9O766HHJC0oYf0R8tKS0pAPlkPo
PnTpkNvPLdoLYOqMXqHMTGDBFK1mtX7MmbIfnZ8WoPZ80yvKviiYpbs3pwCLEzzGvOC3RznrI3Xu
A/srtObv6CMQJZua46A4Mzw9bQ4GT02HGk4kFgNeXP6DwDuDNk7+kR4dlOgt/2RBvDP8iAFPRS6J
w/5FQ+8O0JRKfm5JtXtNOXdb+j/PkGvIgX22t0PLmYahW+4vYkwYLVdw/v5Zqki7bB4Y5raWf8m5
IwllKP132zEaDABA48NS4iaaC4SksLPJIb+NDJkP6afcrAfM+8zGoPFgEGruuiANtUcvTDbkyoex
aFN8TkIHkS3hV1gE+HDG5jCFr9AT2bqQUqe5AdIx+N8M/ntOb8bbOUSb/vHm2h0ZGQWf9+jezOPP
NQyLEHqyorWpKADNuho9XJLmX6IzK7A75m8UADNO6f6B2jw2gKUZYtpxqxb4VWmZogHId+QsHNLJ
cqitUuPtG8+d72nSWhvgQoNdgRadDFK6VKMb423dGzsbqz9CpUywjDDtiACsbYu8mODjLW7LSSch
A212RLAzIEv0ktKLXLnix/PRwU2t4slOUaQA9nt3DWg3b2AR8N/SBE7DE7nYJ8UcZpcqtB6H2ms3
zm24dM6Ad/qDF18m01BKuDZxlsXiDT+VFfwGyPPnBRIODi6/zFloYqJ/2k++MsQs+gDdVyJQwDhD
lDYfX8uY/et4eY+9v3GEWdOpm0jZJGjLNhGEYNGfRE4yUBDEo4bBRJpE4jRobQGY+f25K0Imwvxt
nv4ZCKQb+QpzRKR6lrDfrdRXb8H7aD7OF5edvpYHhJ4l50xeJXJvePHSrFXNl78exADkr6FB4+S/
TBIc6UaEhbGvUYN0bVLUQLNEmgPGqzek+JSwsRhEwA3xtTQ+qWL3J3NU/cXYVUDE1K9L6t/iLLKQ
yVRHnPmTbg9+oZaR+gmpKhox0NI6jsl86y+zWmaxW5RNOGiYt0p6bHT9dUo1B0a1zdJvF6KcRzFO
zHhvO9CzlDrdTE0N5LzfBixIbgY5Qyp3F0xfYru2WlimNQOewKgUqdqXVBQMpF6b6oHdiEQ1cjrG
dbb/7EhLhgl7CJwZL4XflcLPpujYsRGWb9Co1+ZVtFL8I/AAuXrrzP7gLLTU+yx1OpplpfT2SNC+
c+G89db44BF5o04zk6LqVGVijJUfuOHAFvzGX0ldQgCwA2ZfBTCP0mFzUpEsBVTZToiSML4P9GBk
CCRA5cZsqk+Nm48G8dMec01qyyorFVJ1WpGrAbZp5wFDWO8TuR56SEBJWWeX5+W7gE3eWTKkDsvw
C0Oke7ucjeMCy5D00IhRiZt36aReTkIjKJY4347DYfB2ojgsqTziK57+ATpw34/2LuKS76f+Gf9t
Y/mHLE1LkK2A/oKolG5XtyMoaKMpSz7Gg6bGsmveQJm2KS9TOAuie7DuAdYINbkASvr4/G+FIVrc
o+XpFEiYrYTgiEIE4OC4hGfcSpKfGWtamDaXVz6hC7PD6lKt4NnUudxae4sdbbJ82xCfsXxrVze1
3tbvRyEgRssHIc66DzqBT2OL9k/AvH5GFQvaMo3zD2bYrkwmtyGh4SpWgHj72aEknOILfHx3O7+I
geuZwhogMbezHC/P07L0EjiUjIBlTp2kKasvZNmb9MZqnCET+FXPqHaaLBXFsAr12Uwf5OKNrygx
rwUMUptNXYvhyYp8ip8vTuz+wKpVifdwHN26lQfwD01q/CxewuZ4sUe5WrXLHZDRcuWgXnb0PZuS
OiRIdlk1fB1sdxDfNIAxhJC/9xT5OloUQvZA7fnjQFwTUa5roIIGeSA+ggrbv5xjCfunMOUqSShb
Y9HOb63awHPM7S6xJ37LKPVqPShY4UiMng8A06VO5Iq6Eg+jjV8qhGJhti/54noPzyHNcVLhe3M5
Htnh5CIJDFcHfgcO/dKtJfWLEIpf+3xUJxtbaWdxRjvA33Rwf0Ep3TVUU3Z0E7J19jp42Ay6CH0J
5e8mAZ2b45YKgb4BtqfHCTHxQ+QscYGMOxgPk6rTAlurEGP9tkb6J677DOBnvIV+eIctL4FTVkOw
/JIDzsI5AIhjlfeteV1aD71JyqigtRptXYJM6GzoM8NTtl+WZnMcmPk7dXWe2uoiG2HUQLeeVOSv
J4KcB39iGVwigPjOI96nwdMCR5OQ/kPsrmRE8UYyKqPvbktJUTuasYlJtUP28RES1mnQX1Z7kqkL
1Upbuste6GRNValzx95/JMrCl31tSQRoXM9YAYwhMYDXVN7JhsL3wLtJWQaJLZ5XrCRqW0NliLT6
Kwkd6owZLGDFUk+9wXNXteqzIz5LLOL/MN7G7YivYf/xkB/zoypIpGiSl9dNWPfmZIRGFiLY6BtU
tvAudGZBYZLg0qxWG5WUlrXQJcGUUoJllKPvYBJvXyFiD58hcgfJD5X6tTX1sMcK4fkeDh3p/j9W
t8G+EYvo+z9hdWuFoAl3i2jJoOTap2BvEbBr7hcG4TeLUopZQWZjBKx/4yBfQKGr/AaEGpr9P5/6
pw0oB/o1OOHJc5Ihv3xFkFAZRMuv61wOHGREoPPI8LPdLYn3URX7f6NROFSU9uB/jpmZJjcsWopd
MUfEFd3mouhCufQipM3Rc4QnImiaQc4U+Ysx7OogXgXraVgUoCLdwDkpRGMLI6lsNHU2kDYjExwV
rX2r8QXpBwmffFn5f0JedkqfSWT9ql/TG/HVrP3S0RgmB94KXQJ4GMz2ZvDai4ifOU8AJx5QJgCQ
b0QdKr8OxL9AQFL6UfG7azna06jFa8rCOtT5DYj9DmDzLfW6D/9vRETeoXLKRWfi+KEFEc/l354i
eTM+dZH9BPavZyx/cXzQA7vT+xox547jjRY0S7+dAAeJ5eSgwskxCem9X3Hmw7nYr4H1JeqdU3ie
cRdsEA4myxVXHOzOTJ5S4KsmdW9HSFbj6nnsmQf1alFYgOwMO6PHxrStcGTX9MtrHX9xB6THVTaT
Z1mG7LgnsNHvoYHieRW8ymLAPl6mLdytP1Ehe5CQXCbIfeo2n+ANvuoUVJUMRvmCBU0mOlQ2gEy4
5BemyN+l5MHj6xFdQL9WZBGKreYLYePx2a+pQJYT5LBpTfXk2I7fBsV4I159Dsah1eWZ/2oZ4NBV
PmVYgmdoH25nMB2yBqXDUQvxWrtl3/AD3ChLnfjhzMTpRbWUKiPSwnPaOzfOd9z4VvVVgxvEgiPu
+nBEyZaggGaWd+9d8n6aTJaZN67x3lrdcQdowvEHMUB9hvoeO13/jB5sTmmJy5pJocntOW75XgCO
uGWYdsbb4VHP4QVCCrVbjGF39lQniAZ5N3juQ+K3Tx2+uZ00y0V0FnKRyfkcdrSBj5/HUq6HhkB9
gC62Fg4ynX77I25zkKTdBL2KDyK00Pjvpr5EmlRZcCItTp2HOFqLB9NrDNbvlQpkzgtmV12sbYRV
v0WRobbn3NE68SNAFLzt2j8ll6W0bXd0cR95cmop3nFjLD0+4naufAIm9m9yVSAZEBI6aPO2ysi2
46dn4Pzw0bXiO4isgVLjyBVSxybaAELHFpZkBolM9qmcS7jGflr3H5j16gBlo2NgtowFXPUPyoQY
pNLRglCurwxs1cn+Hr8BrVF4tXFycIj/rtqwhYmTLZNjUIyOn5j6ezMAxrq36pUE8Np2VBaoo3x0
yFx6C3i5NxcKQp/jsU95wcmn3dfbIYhJIi+4quPVgi7DM/DsY77TQwgFIPWxuRKX5SbxhL6KTVAZ
8n5EBTNiiI0hqSaByJJU1h18MyOmbKDe7wJqy/ThwspFhdIO+5t1fJwYNvWUvmHIDNhVdCD++tUy
Gkc+2ILWimizkdw/lTWCVp31wPn0dbvHZ9wopHf6vIMNHHueLrDVY2xcQDFdkh8dDO4JaJGhl4Nh
vJuLh3zG2GcQ1gRx4HLpFSopFySMe0BX7NsiN36t+Hskj9l3e4IV2ieYPQFReCmoSgTSbVQqxdvC
Q4e6XUYdJgW+CPTuHRG3z5ZL7/O+VKoYMQVHzpkJ0+lEgvD5VQrPEc2xffgpU080MPdQyvyCfyLA
UwqDFCtdpPf4Bsho8ZpKyiKrPl6Oxv7YsMqKNIvPZgTOF6vzstJGe/FPviNrxdCW3tewxajaRwoH
bUbjKZRr6xramkUXg0OMGShnfWjomV7c4rN8Y+vdPf8BNnOK7Be8urIfGjOapIE8N2OslFc+fI77
YJbd1qXWaWR4dxNAcIb3lkwHTjGIvs+owEahfBRTvz3T13ys9SqmdfXOjK+0F5izk8xv7Jt6RGmT
+aPdn2FSggjOEStUzbAlvDOYh0evwA9nVzqy4pz5wEZOz+2VzSHOVyptEdqlx7BiM6DsBfLS6Jf5
FYt6AnfMCuKPlXRJvkmofCiaBOxpw3ipAF1io48eAVDKA4wZkk5FY53CJENIn+BSiAlYtszehOCy
sWJLt7PalSf0t1lBVhq+cdjhIXCwpFRVil8g96zw4HP11J+CanRiamgErJp4URnqVB1cMvYu/na6
PakVQtRWMD46kByBWWfBucIhBLbP/5mGlFsLpRg/1r8WSDACLfawbQLjf9hTlGJA2KcZlxbgo1sV
uu65XaA7R6rRaP2jJWUD4BHpNRhsSm46KuP393lY2qM/CVlpU2we/ZGQfnALtLvbDs/P854q+NfJ
ZCl4I3vgHTuYTQlo27sy/UzPfZ6cqjMxKMcnNsRmHtE/8ZotSKMI93HgV82s4JpQy/K01xW1URiR
nEq+9s1SEnkOy+1X2BexlTz7FBsTsUtp1qPZ1seHTwcxrirKzPUgWCCKD0KK1xb69J1yYM6bdqT7
LDS3zvJN/VPsKIuNn6oOhaCSZo3wI0jdMDcaS0k2BeIWAV9vWJViBYZIq6xBuJm4vhAtMbpR88pU
hEdwBz46z2r7CLWND2mLiTHhpKqk421qQ5/hDMr0d9PjkvkXt3TQssMpuqgMvGNaaYmEt5A1D5VH
zHh7K1uAMW9+F5ieoFX0znJ/fOaicYAmrSb9T3cSuFWKs7w3vo4QRFqswufLKMhWJmAqVHock6fW
jRp07JHmeTZJuoru65/px4lOAbl0Hb2B3HO7wJOBllRhs+OQqIgLE+dZX7/gk/fVlfppxxLM1CWf
30otzurJ2NaWKFMxalcW1Ltpqa/MGhenR3tsGxes+Fsao1IuOkgucqznKkNOT0cksc8B5XWR7X7a
Koro04FpCP8qut4r+6fHcBw2EknpFGtoI0DvZt9xTgeeRDr10T9y1n7mhjxUDtwFujMHXzqM+/He
8KZ6Mo90aWsW6cLNKmTeJdHgMQi5uyCHV79LcdAUlSzeocURGBsb7/6Ow1nrtpyqag90IYytaWMN
HH/lSlsNz++8p58P5aTKDYr1l0Bmh3nTOOptOgtK1yXVZsH3Obg55iWlOh6vSS6KEfnlZfNqrcR4
iEgFh+u4fkmZBAnJ8sYOr1nfmD1TmKv8GYG/owV+Qe9kj16fioYUKyu8z+mYjKScHKN33PO5oyJC
9OEbjZqkIoH8/omn1FqdCVyQKdWbfo943nfXScDsK4b5nugvoHYc9Fw4KOnmSuE/2RGHmugBLAcI
uT4nWnHREskXdRuTNUUPac3n4dtpM35jh4Q3mZ6nKTNtU785vC9N5yNTufF9osEhr6RXgTh+nM0O
w7c5ss6Fb4wAzXXXErVlDqG5XDO7NbhVGeH5odJExZnZ9IC/8ae14amwZULSfpH4xg5P4W3PiI+b
7SFIWPYzwMlW6/kD73bu7xN2A14eL5pfNUWrmo4wSTSvWU7hiV/PcD3W32gRGlAAaiEh2yAmEHDe
iOHXUZMsg6CDtUhk2RwNFg4ZhHoNruxStoO5jpcRaWtE6YXj4Vr8mUfhaJjAjDKEvpVoqohyiksi
YHRJUJzuHGxqme+bIi5FKMPaqGxGafGyRc6xgHg1bvipepnfQBSmvuNJKHnXnJN3xkHpvZHEuMFM
z7kRNY7N4I0x37rs042+56vFy656lVwsGYTVkEe2XVzsGb92YoZtP/bEs1hDf53X3t91azuF9HTv
TVUdU3KsIbRTtYaYH1O9rPqGYDV1Ze4JpdTgB4ymNxUGfHI+gEKaxJmJSM0WA3ehwooJzRwk+qA7
wvGJQxaR4X7Tp1hJCBz6Klkftp/hHPzRaM2TzxkNB9aMEaekeAip9BbCAkLIPC/boymgOpBFvsOu
k8aniIx6LjTl5fubM41MGMzieQx+Baxsr876Qj5hdx+Sqwmb15NbM/AN1L1eQ3YlRVFHDzz9tpd+
gs6E/WfHi64YAKXWyxyAWfO77afJYTa1KIV/RjQl1+F9ZUHfIDwSbn/VJhHdmthhgiHn6B3MVmLo
6rUNdDAKCDTBV7F4+PgzJUPFP/TQ1FyChhZa40KsVFw67yeIumJkvesHfwWylN5Oek80HC3RFohp
MPxeqJ7rE8pCIuhOEQ4k+ZxsAHMVxV/PDofkN0T0R2Kgis8FSOGvDyDebLDFu2IiSbj+MfnMyeKr
wtIA5Nk1Mpvb2rYsqqDXEBd/wijFpaKdaXknWc2kzLV3Plr2LRN8IAGuBG589xovkvSbSZ8Scwol
J+JYkrYiTGORSveWF6uyQsSa2qCbQBZcufHpyZ2tkbjgGYuWcwnWOthVDGTlKYGfwJQfYT97yADR
EsavuZ0H1dOQaaMvCs+7fw7JWOvGIwwnu+k77zZvkDOiROd1Jo7oHjkxu7Tsth27nXRAUzOe0VIE
dO8hdMgYqESzCQAgLPvBuYZKwsfDMbGXTubY3DeIQPAltVtWJXshD3qm1mYkKE3//Ig4X4JB1aI+
pNzJ7r7EH/v5++50aJjE7StLJgMH+KBgH7YM9pyGJWEVTSyW4D6EindmhnM99OMOv/zEKU4pQFAc
GLq2oxTo+HB+R0tFsBHqdISslad5F1zIOdUlIytXVz428WGQoXks4WZcFPoLvwVtiMVrYuoggH1M
mdLlgdHo22J7dzn+sWBElQ97ebDuC7mjdPYkEuHimfg9cA2Dyg62DxoUXbkbgcwtBFp6SYpGdriB
BIEfjtvfjK1zZOg7vxTx10fUnrdotaPavboy7Uty8mpY37UqLpSXldqxOs1GbnBHKKvFGKVeW6Cw
5DB5gpaG9nmuK6RuiEYRfIsiy+pnsV9DnnGdr5+5LzZokLaNsNEtbyr9FzVwvwCDL/tXXZRO46/b
XzEleFBHJzCk9wBbRDexHLSOdMqaWqcd8aU+st7T9q/oB+wUtrpyzXkKcK+fyCPDSCRtnczfcg6X
CJGrVPGA7rXhP0xz2mGtadDsHfLEFo+75SItfKcElv8dgs/jk94RkIpEzoJt2jsZMyhLKY+Grl+z
6I6rDKQHOBMVstz0nCIERwBzhXktpECTKDi0cvJAkxMMZzmLWrPuNK78J4qDbOZ2/1RKgAcp5nO8
VQ8RcIfB0RJhjWinf20AAYlGsNgd+f/A68Y4njOxPAWSopFORALbgNXS167rgIqV+BKiEW6GOXxK
AoiEQVwbGsBgYfDDZ9FJW2AhxRGrCmzjADqBzpXa1p3gYXf+FlDFKq3jUIZoRvcwwMwGflcCE3pS
/ty8OmjuDUNHyBsZK/l5qhVTAt+fiohz6JujaW4jZOYocPCnyvfPfZ7JBEu6AHvYGFD7GptnURDK
j2U+yGUZdJA4MYRBLd3HMCXv+kjG0htbytKeHX7yDMfFOgV7ktsfyW046Z1JMpnrDgTNuA7+t0jQ
K1YWhT2D0Ffg5At16I+MIlknghltrikq3pKwgo9Mzd2Jt/o2yAE55PbVOWvhn8XcrrBSKa8a8PuD
NAksMwrPmyJmmf4z6X8Y3nazjHsnaAmlFoJK2YJlWlLxnklOatZa+mqXxVKQfedflJFS2wcStaxY
sr3UkzrC+X9sIbvYULb6RbM8dM018HiWDa8hlsLyApn/NOQPg5F4GH8xRSRCk5MkOCPBNpEuwU2S
bY8UThGUzcuwa4Ufk1ANasy1ihVaceikNslzr7zj/OHnJfrth1UQeQIhbcxGK8k//C/hsMgeRCiq
OBoZhWILWcEGqY2iFku9frTbjk7XI5MAIKxzcaEBDjRl211qryTXchPSzyajODTM5ALejRjAgHiO
7CLaiH00hlWhew2VpZ2MrxpF69QfbG29GKYyDPgvAw36XIKBVUOAhIy4bjoD5CCSvZXMQON79Jzo
IZilr2hdHKawBTpZYiwlWYIoDWtwEbSmjpN1ulBqqdYxzeepznahq2Q7Yr7o6+ixkBmOXii7+Flt
hol8Cms3GJ4XENRTVCu3OfDBvdYcogpqU+PbZ2dyFWHh5UKS7/13E+o7gU7zffI8C1EimXlHnyPO
HxhPn8rlJlT0ePWK3yfTcrp0Gd8rlME9GYE+K7mLXoeEzhYc055IIM8Vd+ylpumZ3VnL7qWpEArl
Kcmi9N5czylYnBlG2iqZKXBSBPpmuBVdPDypOJVu4cnNdCG6S+8vabKU5BFiHbSRVCTv3KK5coVU
tKTLSKASkEv1UsbqtxA2SuPORJ1Ng3y+/ViylVWqI0me+Oe678vrr82ugn/xMEg0AN1ACEeAjcnS
EqF6d5MmTCgsotTF7bPsjHNTHUl0fQlwwysBb5tjkVd24bIPRPl3bHHS0agBEg518e4nKcKY8Yzy
EgKXG2aqa6m/52/iCYrD7jIWw1KdndQFKSjdHvCCzYeGwwre6GooEKQU6UoBTY+nbOX7my0+EefN
A4xgVtWJZy+leJi5L0rMfexB9K9QGRClV+q3HxU4Ivthx8Ig261k3c4EauCzZQRpz90ZMdAbhPGZ
TTD9sp/YZh8bymUPKmBXhgztjDYwAWqdSb+m/lhNA97SGuYc2uIsQMnM+x0FYtXntR3FC4uFfayK
NI13R7pAfSfX4FDpJNSTaiWHlNHHTaDOUNnW6qLc5oglupgLeSGt5yCnjgQI0OBkO+mlrzAMH/OK
RtJ9JM3qGcmMIjf2BJH7VpFJiYonX1q9EDWvoBypVjmcM5rvy72B//e1t8H2K+KzEFimRhgLX+5T
FFH3PX/rCaAKRzmvzLfoHva0lIxJgNkHEaJr6bfuzCsCLQDf7gLmoyET4CN4y+8WAb60VZQ9P5NU
52oR5OFlLYakJfowG5nYcPIWJ34wd20gWvF8MT42MvBkyOubOAgDmxRvBZcDttKQohbMt5iZuPNz
0gBLKK6VvLLFK5Lkxp9oeivd/26GjC1uI5l09Mf3ETyLmq6jSMX6Y+2Ahj+kVhzjXXXyqYqAZA/7
R/XXj9M4VMo3hWJbIxkx15ikd9MyYXa1A0xXCXr/0Hja8DSMqAoNitVjiJmeHhp6MdlnZIqOUIrM
gzEPElIfAjK+s4smWinkbcPTuvIpqch82K0aNBhOVo7mk+nT7rzKwtj6tUjd3ARL9zUnP6+cPktP
lmdhWAtOYkn6mKNd8/z/BjP2HkEpQs3ajyYQS7oTcosjGTR4fy874Lkli7TPhs98m4+1BZvfeHkV
zAuZJsZjz+UWc0oXTr7o2bVwYAzXDyCIJd+chx8bKNRlOiMxuZt8wsr8zkVQ7eEWtbcqxFxmcs87
j/O4Tr1yJhuTTF61+tFR3WahnID7u6nbPCi37PG7GPXTjFCRIypegz9qWYvuQxR7CrGucuuJpagG
6sZqJLUlbkzdXFH30zAHMtCSrNc8/l0MVuQKr9irR6Tqe6WBFesHEohV2uOBvGGqx2kvXXsfqjfc
1YSU1WH6O+zQWPR+jwtTFvoXdKkk+w08hrZ3X3ovPZw94DyzH9OjjOppc2zY1Ad1iWi9f9CLdhpk
EGvMmsVEH+ENvTjJaKpdTtaDMfYa0SEv5sIVALAoULP5gpbRfRYp4UT+cNHjTIVlmajHlm50KJ3p
t9Agc/qM9T+h3oVw6QFQXl/lJ8T1dvt+DIWERyejPvmHJopa11qiLNfuM9ITvVFVbxU1apDx5fbI
eXH9w6xUMWPRmJGlGO42bLg3t9cli+RNz7jgJIXfyXXoP0TP57WuHyk1ntFnlZJdPEOQJtGsezfJ
wzgWcGHVc5h44YSZalEv2EGQdTBxje9UDGa5dEE1H4G5Pu7b2TrCtli36n7upxDKNdk/NDDlNE0I
Gig7SXxwU9svb2odEfeMKhIyc2q6kmebyE3fAdH9KhbOknYqkYrdPvqnW42ZM7idyzlMtti8kFsO
n6cW3VW/lTR6I6TCSx41hmuoWLKOycucxXv9r14wYWS8oENE9YAFBXvjRRnRweeYapnLWyYck5eS
S0e2tJdaf/akTajcbbTwzIuLM9u7EhYX4zqWLmzy8QmQtGDKZHQbezkIHbCgB/9fgFpuawtPNig1
zwKaUGXypWlBO32xjw4OL2vFiJJ60rxysjdDlnbUMq2V4yrAUAIFaJJZy4gsxlvPHcPhztpbxyl7
z+Kb+2lgsIUEk7JQObVZ8LFSW74FG4QMpO/DLIOTIcN3lpXxrEFFkOhwaMuwQLD1D20Kdnz7DTnb
F6zNnbFtAlPXsam4GVcY7LdkAmqp/uFIEWv9mLihN4Q6ETKBZNOdycJusbM8vt4paSVUT27T9K7j
wQcNrDxX5isAFofbn23Ih5uijp0ZAv1r74HUCLwotLDLirvRcLHo8+Lk6v4sRGeSPalDTIRCkJFM
saVdghOHZ4SnQ0H8Ao4b1gEhlnXzcUGvOpZc7m7fO40Zh05ZNcryjPNumaTruRPJFxPzlbrNsDSq
6Vzlp8IR2btdtPkC8MGfpYSRjQPf8DlddNzkGTURvCyXuKTInp2BGGBSVeK9nuozeaQ7xlLr02yj
cRKEz7wpHcyXwPOiJV+C4/ELbYCohaHHSbYtTwY2Y22BrQCXZDjKZY1SnNuzSIEkdWpquUaDaUv2
lchmx3xYEbP0M8EuenBGSBzdXUwRdbOHpAYmLDeVcS4de4xNeUee1C3e/PdfmETiBCf8p1SYt/pp
/LIbNuhjt1wcZF8Z+OlJCm+tmYc72HSU2wsyVJQ227tJ9kchCVWSNdvg8hlFiJUCXnnXBQKK4zCw
Ly9DBGKWt5jC76QtegWcJRTKXXgRI2AtKyX+oXjU69TxYjIP4AykbhDdGWaf+rIpOZrxAqVvwJ8n
NgkyT1io7E6tLty0uBq7LBmvMUvj8skSZz1vD/MnwXNnyBWVGWv0HwvU8Dk/mr1mcJ8WzwRhRKOo
ZFXKa86VAK+cDBMHUEYQUfOMxI7Czxy6F2IEU1GmtqZ4i6z9mG1hQcEoTN6En4XCRKdOELq7/SQ5
d5PSDTV1xf2G7F+B3PtQYh0kRZWGTAVwRnRlZRYEANzqght02mEYe0hQenc5xrnUhLuaif2538hZ
lAGApNOXFCySAJwWwYIV6Wb45IxpFTh3i7GnmJ9jSX03y00ceSja9f9kWDdJkqTPS2sY24RcDBMm
2Ie8cG32dCUtbCLzOaFetffvUkrVl/DIHLrcDqJM3DpZIFYVpypCGatfJV5+cAp+iRwcay/qbfO8
RAsCmj0/mLVMcBFH7pnfyWuRpqXgg/QYjcG0Z+pLdo590AsbjIHB2rzyP70QFKKr+1Tz3XYvZ13d
hPArCVe2huKDvN++nZp1b60EVGo/h9fd3bjthbSIidKrUPs0MUek0A17L31EAOF2bsLDYBETB6HS
bgDGOl49h0E8johk1kqm1fTTs3CCfjlvckfP+781czaT+CkWnoHA2JjOfNo07NOZRTr9Ngb/JHb5
PpaDLFP+clQ536Eaxq8Ov0Snt5HcnhVB32k3xlQm1lcxE7UqsN915EzAxDLbDYshPT2LQG06BKw+
3vrQgJD5eXtTaE7Lg11yFfQj4pTfeuImiTYqk4LEBJ+3Q0HAu1h6dSJQ1wb8DiKRk4BPQsOy3Z4E
+wCeKRM4tNUezRA594Ot8Lnvwn8iyI1ugTcBItinMWh9bH3++RKIOjX9gRQOLpsW7Ps5AjZxEnyP
JMavW5n9jY+lfImvHXKhDIjzRwvJuU31Gfi5nLZVlQwH3NXFJ4wJK9SjtPrjVRV+JCQESt2dQmO8
Pzz8fZ8EoPVpUFFJswQCMYCFDd8pyw1wbtRAYf7IkTFYI7ZVqFzOmWhDjzPxKTs98hhmE/vBHp6N
9o5V/6BHG7pKQYWKAKd2iwVa6h+SjS6cUH2+fxETUNOia9fHNGCXSqiBXsIsR7p+8mWWcpR3zLqI
OY3brmDVybD00ULaIOUPXFQBc6AKW9QDjDJdhTaOX8l1qBkCDvkZN5xbsUxVeDz7S+tagsHoJboq
7+FSbGtfgAq1+wMpP4Dp7gGLzDcOkuvQ0jjflGKzWDUxwO7SEXAciiUjjYlZB3avS5QRS/usAWy/
XznrBiJekgPgmkO0zcKfdcxIJJjZqJA/SwuadpjVm1JCxJRvtE6rBfYW9CF4O+X24ieYs1uM/vr7
j7xrGRvB2XA2cBvjVQYzYwo2f1nZnbB1ML95X68TVAkcRKO6BThzr5pgKPBu0qgGDTY7ud/OjfWO
iNUOdpNk1NyfsgGTjH4lKTEcUmwx29VEfViRxnQsCzFtM/HkLgq20q33K/KD4NUxuG4Mqaw90ktM
ONZKZ1B7cWhk4sr+/nO2Yymy3wR7VkbkrZFjJi+MejJg1SITOkPSBw5IdgnHp8n/PlgM1YRGni7o
b8pIyfEHdprprTj32tGc+vOs9SOTkvYnuShUEH/aIvHvrD/v41iB7YflCKeyzg+DBfszwxJwz+/j
L2S+xSUVWMNuQZf/YToFGrFhpLR5rC2Ut/MK5pCcXmj/72gPBgKHGEUYYCy7PrsfhWYn1J6c5FfY
uc4pIpaEZvbTPh+2IIBPknNM2hlTBsktHkyY+YygBCyq0p8hYyKnKbzKnq8xR7fmCyika7tdMFsZ
9uCx4WBgfWYsjiAzgUFBA8MNz9t9CIzacQOMGHffpJEf22Y8lCr5O5OJuK7BUZDdT2UIsgaeq8Ak
zVVJxCOEFoDspY2eqJCg0N/lcQvE79X/X9/Y8DZKwGPG7K9+71IEjr9M6JkZYmqk6i011WRuhb5p
ICl/rN9VHrTTbVTVKN24QSgvTudhxZCIkNV/7unnV/044nRN8t9UD6Cd157eTm8JtIhZzHnZjSwf
p5aLDwhzgJYTO2u4J6ZKYBD2emSxb4FYsJU6Kcz6upPSw///s3yBP4c2i4fStlbSTKvsxtYwIYRF
cBtm93ICEhGFEuVimFgDhB6ZC5YLyjohJhI3OmYOUNhynvqlpATTVE+QQDBB/utS/HTjQHcPPHOe
mTREWSTQPp+an3pFAi/egoeSTpYRnuIz72s1luBUieCxwszX/fhTPc8XAQtEXu0dHmXpwDf1WnzO
kxuw6jVReMcMuLyschuBNiG42/4xg4Yors+yfs7ZL9kfHWwdrVsGFZSp4hheBU8PHg1XF/sZiPxz
+lue8lSeIjNYrXONUT7/n7ZjbWMDM/mRHPUZEwQggVpp3xExm0s+tPXqK2PX0dKu1O2IMFegUeTL
VKF7rLvDae8REXEJMq1+RONQruXxmEV69D+2Uu0fiViaBXs+6e5ONMCmdrw84QFWLsGJ9n/O52x6
pCq2fpXKWl8AofEQ7Vo8MvTSx/3wks2R7Aixd9DdK5qA6YHdEBC5QsLwlI48QhzhaNwdbxsltgUk
dMA6mwHoJvSHOwad2rzn7lScUsFTxzL75K1WIWbA75Z0FK06ozW9x4bOidnAzi8DB60fSxDmk12A
taATzMNVvkQdEON3WphM/nK72WQvbZnFfPWICqTCKg0BK0kAeGP1EmCVEauOl1zWmiFLK+6wXS+9
pMj3xljVZw7//K/9lhiWE/h2nPk0unLsyoyoBWD6PHLUWCmfTAfQwsPk87zQjED0Dydb9RZ21kDd
e3MQhHjF2A4Xs2QfVLP5nlaaRXnDEgHQ2Z4ran07SfJLUoDnz3nTZxzYukv0V8JBfLoC18v4ZWQ6
lDrVu9h65JqtGeWHZySuKzOn91e+im6jJlBgCJxhh+/NFv7Qgsr7ozT7M/AHmudK+vpWPi2c9GWP
WyoejQm1tYzeXpXOVVfvZrgVa+fnVf5e6L6ot7nWAuHCne8cfiinlnfHZu869FEv56lIQCyVRFyZ
K6hxywLCu4VmUY0tib0kKfD/TyJIeQemAjHtkuMw/zABbTisoh5olbxXMZOiw2iJ1C4o5AbixkcN
iTBqPr1bnwLmGm5PuoUmyn7tBVh6v5JwwKB3KwELrVdfZalVgqqBr8nBZ4F35LG+6E4LEmrVVSkN
QYsVOaVrnWpjBxvTdk0zIJMkny43F0K49zn4osxOMVTaNSSiZ4V1sHFcecIXoI/SJfV1yN9ojhMQ
5mVk14L8ASBzZMTGBpLKse7oHHGm4QKWG+XGognzokd3rWZts5kPoJp8o+/IUdyOp/EDBRuixzBN
XFjPuidMeoCeeoF4Px5yHwi0Ti83MyPhPthZ/2HwZkpKL0LvMlWk5EWCvmRf3D4+bvWMmxf7obYv
JN46tCa9jQi5SRiCfvbSP3V/ByhKpI0DvL6HN0EleHE5vJzt9orrfpIVWcs/vzwlHFLlhlMsJgAm
HR6EgfSD/VyWx0oWiMQ07O+RmIv2qccNm3hNgqerdUtne1cokggQ6/5CiE2aiZxyZhfThWQQQHmj
aYzfWZ/YBVXn+Xoa4IhfVn3dPtedbCv0jOcQ/4Oe0D2UtGUcMgeiEw1DLmASNTYmCZtGKBMtW3h1
ZFVOPFk163q13InW84m42Sct4BduBHGYVtgF4+wv2YI2lK/d/NQhKfxK9Dv7KX3Fy/SWtawobY7p
J19pOzi3WpnKhrNWk+3JHj1dD6e2plBffofTCkxSKh+WaE4z1rJQ5zr3T7Z4HSKg6GGwcIjvP2Cr
yacK3/LW+dmKLcKvhp8C1xV4OTBdoE8+VJ5YnANfgbdEKrrQfVWGvTdcdQZdFvucqAkN3jQnL1Oc
JxBX8NWywTAd3DeLFFmiNpw1x67ErRvzc2IA0yjhsdUjqSc2k0whgpN69QahA7Uyy2qVf6+ytSDV
ga+HJqGVhMWmX6N+t3qkvWMD1wF/TypRvYn0v+iN5brjhVxl5t7eixMra1A9M4tO2pmnxbPgUOQ7
HKw2W47mj4uRYOarHcBIIMbuNJvkF4kBM0aIKShsESNaj/WWJXbeHtEbSiSkTl1O8Mw/3IhA0SmZ
n7cB28C+EU4/IehDWeBBbWSRgRN7nW5s/ghspR4bhpUrH3XLURqg0M3SyIwNWgkc6y6qmUBk/HA5
C7lil2QUJke1jxzXanWKQj+2ZnA0A+MwgSXs6QkoLQY+XO/MmhUNc7oWdNoWZslT0mcHX2mWrLIq
qgP/hIKOjeYgj9QZlT82I/0+SgcF97MNqjS50lTDWdm7+nZG7RDK3zYbSgPaVyZosFxjjpYnebD+
OsOiMY394IBViW52yLs5zBOQMRCR7jJHSSnN1yaqMPKvJfUrxj+FzbUfLjeOq3GI5eylrxuRJyXg
bH830SLJAGGKJfoP6j3CKFnqUuZjLB2x2TydKWrONv7vHRt+u3UeSGflEnMRSQsrfDLlAKllfEuq
R9u5pkYf0ydZAR/Z157zTUe/yLR3tJK8DZd2ypRW2qk5QgJkkso1GOsXU7KtIb5PnvDK8KvYoL0R
B4mtUNJbHRsId2eUmi4g5SGiQb9hxbq4qkGIpM+cROpAwZ65/6X+CX7j7CSswC7GTftZZdFdjWgs
rnXRa9FWDwknvCWgnzkpg6NvwWRyuBgnEiGMbALtuFHPkZDxGI/so+EVrylt+E4UhC7fD1PhlNSg
pdtBxWzBQohAqveD7kl5KwD1N4VTWyosrxyt9GzN9kLH90fZ4YVHdt7v9QfsbJMnwz7hTL/Oiu/C
JGOxXop7BDY4lPZUUighTRNZ1aAILwX3qFCSv9g4cg1QGMldg9fhNt+DnH+z7KurY7lecMPf0vnG
7UhyhALuBdKIFeRhap/lzFLfgl21Sf2CZRAmC0807UOVFFeE3cHzKSo9GjJ+Jx55vzOTmZ8fDlmK
M6HWuRFxyWnEng1zGnlX7HGbpbc8Esd5a4bUUFfuZ/PH5JeLOs2xa7H/rj7x6NzjMyfU3cs0Afo+
k3sC+8KIYydgtAcZWySyCifY0Ce70qgJgcrLkjdILp2W6+Ol794e3s31IdQfYkMnGy02BBH9Ilyb
mJCEOwNADCZ5fg+a0K+B0lGDrIim7k5ASaZ01FrG/PT35MpFwFtVFEyyeSaGtmHHE5wc2ebYKTdH
ksaUqQeWrU5I8Zeg3X3pNqVzhyJ0y9AYfqWEAw7Y+fULgIup5nJRnSn6SoNbpo+U1ZeMJLs8Nl0D
9hu9xmvW4asi5hSvhsopk5q79qNk01DmO8grK9uTzBh0YjBJ2p2ta3++KF2Tp+cJfABcRoET+meu
oOXPqFsd4Ar04NA1AalNGOqy/R5g/ZJzd/If9bbSp4AIf2iwjYOd5mWy/3nxw4L8pzZHPqkLtNiH
WTomvfgIJAQg5OJ7nPlSN5PXkbiEMgBgtAFQLVg1kk5vubcSE0zSUhqS0YV+yR/9qtuIzYeA0SbA
NvWKWsgqy8N0CNT8lCHV1srddI3vkZ5mz1sDl4ywAQhpDUKtG8ZT9kZMiFBul92YoTBHNo6VaKre
ngeml48ieHn6QFB0VHwG68jfILK4dmfSpRlcsGKV9FXCu7RE3hf9rlBfjcuZKpUJPNBWfxKvnE+S
nxtpW0wkMO+SgQF1p/z++QSjVb+L/4LJWhx+RS5tveq925YdOp1AhCLnyfQ+GNpKg3FgNoasD4cD
Jlt7CECh9B7s9q1/otPh2t25ROwZYRp0dgjm+ErDn80JhMiPQziYJkOrUd5BCOV1F8BMaIDv5wYv
PyCnNz0VUh9LnHFw92wmA4Z4Mvy19PnppT3ONLUvkvoDPwwnCrE9MJmS8ouIbLoPetQvD1ePI1OP
qcO8p+KzWAC7e33hwpNxygiJ2lld44okq/s+e6KBK3vSdNCpQXHC3EjpcOO8dmtzfWzIruWzNQnA
C2WvLvjZ2CjUGvgPebgBOtyKa26yOaMAVUDRkZvUBH8NH2vUoFAQhfAosIMZlbra5E8hTfTVSWHT
AiqQdwGtWJudzy81D35tvMiQGCFv0m+5tTkxXI3w6d2n4fsQuD2Uy0fG0DNlmp7iCNDnu/SDZOmr
bNXRuFH+5YMf1QWc8SH0B42NjeZv7cVPjTx9tDmaMylhjwsvomYrJgMLlotxNWQqeKSVvTcG2HLx
oFBCT9wygG4rKsN9GIbGR8NmInMvzPm4UR8c+GxkD6eyK04dA9SbHAAf4BkS90U4Hj0N/JArQg5A
mWESqGMdZMlqqgbIeLC+JnEGwBx3ShQ94VHzyTvIeKamM2KL1qi3eIktuVyLIgEC53ip49qQfRYG
iXRon1ugTTTBKvwMTiZCaG6kzl4gsHp3JRXL2iCE7NuLF8Y6Ku/unE0KLgh/mgZUp5PrIxDHT8YO
5rPvSinTdu4h7gDoYets3pRWHKd8n2kqueDDJpDK4Dho5LqWaoiQuONG6tbMW/mAtFXS13F5BM/V
B17xW9EvOmQeXOCtIDkIan5/WDFjDNXO5NiSYd8giE/Q+HcMrfpnApXX+itvNAB5S3BZEWhdGwhy
3IfMI6p/M2lJcldZtSP9Y57UsZCzJ/C4TZ4ELzjEK931jZ5As0CiLrhukz8XSdXumCDKOgEHNRq+
cFhOXRdOPZmf9eI7Ume4ENPi/J/eyEshrE+9mkwBLG1TtLVRl+piYoadcxJmZ5Rfd7nMFm3owjQJ
8SEVRddU/B7wXZSttrH2kVcJXvPED+SEraK0VeuZX3n9a0sNBXRczplS6xnX+owz2Bok3N77BTL+
KgUuAx5CbF4TnVAwge3IWjEhUsKV8rjGYalWUgwLtT/TZYTo6cZnHMkf2n44KEXNtAgr1VdmTgjY
nQZ1QGqG2ijgr3+0hIllgF3khd/5k5mHuxtGNUpmj4aINrMOJMBiyEJr8fNmZgzNezVBBgeb11VO
BRF6efNBZz7988sZ7RX7GxWybehyINJmA2+gAM5YdevJSCtATLlLAEKuk7JANBfETTeewuSxwDHE
6UutUrtfcl5mcRfyHSvTLSlJxT4Nq4f5Onp5shi5Iibqenr8f1FSk4LXLi/TskBxIH7M+0ZrsLdb
fzhOrjGirBi6bJeTRMQ8nQjnuQABG4ZBkE4WkFvJ+2AlsVSt4M8qy2dpdciPhBNTCwYzPeBJbCZq
8IW0gyjXAJ7w6+7ekfsxAm+ExCUTj5JAeVnSeQhZ+wkA4nN8B8pr+yvmY7ForRfgyeCdZbzMIbcP
tgjRWPzjnTwk36OEbOOdvqy3wuHNzbq5YnejqbcG2tOQBfLnLQPKu1PU5VNU7HClJEjRKLmyZBgx
7ERnJedSHL2jZ/geDEPHvRAzBm8TazidHXsCbJ/aDYD7MOMplYAPYkBvyIPldRk8FSWjFVgkT6Qc
Rq+JeQEvLpMPNqJ7XBKn4eqPb2yL4MHFPOfrLB1mRQ3zs5LIHXC+5RAcW/dGM6jRX7a9iCRveB1X
kBB4uUOGGQpQJgViYOzKkfGM6zMbc21WU9DazFgdnyO4ax9Ud8DxOZbLXXd9o/lrYT3R5bBtCgC3
7LF2XKDzo8nM0TUcLbXFH6KsKVm/vKZ63QycuGabnF+BqdQGtSiLaSy1zLlSLfQQw4ybVmTiM48R
AbtzxwlQ/vASBzABPGy6p4arfg5a8wjMqvlxxSzixDx+SA3hXK+vymJ9SkjuNr7lg51zgym20Go7
KzO6c7K81vB3U+Ypk9YgtTtVyZnpe7ipMn+hWgy8NQYcb1KKq27DukXJpbYSEfgaI6MZ8Eahto8A
4kJbxG3a8UnHFuH5SG+mXSc/YiSZ2kyj2J2ErzJRK0NstjT9VeKkw3M+wlNVCcy5dW0gZeCUJcVQ
tdooIq7lUfoQrcBMKumotfZ4OowWu+sl6LDGBKDA9KAJ99o73kqK7A1qsfsHtp2LVTP04L8s/7qA
Ha2eLO2AUJEX6P2oAdSPkU3FcQKIFThIt7VskLaVnGo/f3OLs9irPIJURew8LCwZnAEuy5pbr4Br
23o+EsF5mbQlamSqrzKdOxGbgyI/zCqdUIP3TS598xJIUtFKrpq7rXw7V1C+adwcxW5Pkxw192c3
+VarNXhAXGBVq+onhGqXzeahPjDF1q6o1wD4gzOkHfRjxT+y2RTFBxaNiYN6syChYeEexc5uEF4W
mAGJTvJqmzR6K3REqQcqWWHwyYn6evWHEcvpat7QKePdK/vEEg0Out1hAxdjELDaJZTb9HvmcG4d
knSln7LGF36yqe1eoHTtnfBM7CTAIg03cxBgdd7YbIkG7ayX+3XNds1VLTuuWBH8mGPxgDzItkAc
+kUVg0ogFPtQ+k4nww1GZasrye53xQLEcZnj8ZS8G/FxChjVK6mp1tsEG3/AEbMlf47nxjqSy1hM
/I96OdGY45UvE4t6HZPP6k0UbmPmxzMiG8XwtOSjBiMvOWToY12F6JTjkwRC6+iQSdfsQDcoT1y+
TzOsIaxxL8k9k0CXXe0q+HbQxkh8P5db+BYTu4IOZocF/Z87NH8VrqQf5AgAYsh81iFkoN9qv9j7
J8IVkakP+KfEH/AsgZt9TD+B+/ok6Bsp/2AS4wsjTJAUM4UJiIyR1egLE1XXfCjSrEnbi8/2JUCC
ilvw5JemhhaF/30E3GjxR3ZtzRnf4/WVQnDstY5ISD6veS3ffRE19dNtS/NSl/LKpt5NVND6GUvR
DaoEoXXzhvBmCSD8+70ZBvbJuOfhc1L/9DbuVzB0MAzRLNYmuiAHP/dN2FMmmWnhGSRMe+l3iYIy
lWhg3hO7CnGUj5dvTfwmzmMcYJ/sGgV9ZIM+dkz7SEu1/VQS9grEYqwQFz9McF5E5z8oXFxPg17N
EvmJTfELDRsI44jyQtNFZkNIRKOuq1uCFc8KLNq9iS2l1EZuzGs9wczB9u3wRCi98Q75fzIngE/B
uRz+/iZ0MeZifb8fxtmeVMjHxcjUUB7ojnCQOJmwMDlWejgQa/chh+k7KldU8ba7BvXmANaJBE/f
mI+LRZDzppxdxVm+sG2u1NC7YlZ5efZWYtVdIh23TYbITA2BXIOUjctvDfg1IatfwhWO2NbrHsQT
L0mlH69hQapVwjiy7l2K4mW2yPZGCZD4RkbqzHoyqBcuNEWL58E6OebG4XMQ2wik6WkMyAMFPAFm
KLUAiDqE/ZooRyswJiuCtl7oe0BM9HpbHjuVBSgbGHPpA1raZ9xwwbGH8FyDuzmpt3aj2k3dS14r
bkmMQZL6Ep7F/pnsVb39W1UoqBczW18Jpr/Mhw+7KloGIHuRR99zUfxrFtylfn6q8RgLhUEIx0AR
LQyldbVjHj0DCgrWP/PWJroCqlruaLulIycdmycRwM+Y4Avc4LadymLXcXcu4uyzD1gw5ggAE3N3
wLssOgF3Mini2yEPoN4ItZ0seFnLvruy3qdB8RWZ3TaIb5qSyQqw8k0OXn0TVHV9v0mSkXdg1jPO
LKF7yZauZV5e29F5lYekH25SfZQktI2ZBfcYJ692AcowkjTm31SmGLonsI6rZ5nC1l8NumVAt8A7
FEFcNNbj8nffn1Msk+pHeCPv74djq5m8+g+2YB6o2O3lXNarKGXzpc3kVNsorDlYucojTcEqef4C
q+nBcTaf4AFFlJGx2/e+/OSTjE6v/ME/NSNDe7np7uE2MWjRtzEoF8xdzy4N4V7bcEehKW9D6TDL
W46w2771fSlRteyxiknhdlTrSlt5B7uQ1EXiMXfOOWTIwv/te2XmU5cafqGT/ZWfpklyjAex3VLN
cM7e2/zBvkfQ0dWTDNqjaPv6+iJ13qyuLyeta79ZzuBnrCzzNrbFfhnY0Haft7TibkLkMmAGd/Li
YqgvfO+XFCiXl/H4ftTab3llrpl6Bddd+azHbf9sKq9Ifv4DN2KHQBBeqPnkVfn55ifGrw0bbT7W
SMp2Z6SPjqqRFGeTX8xbHJr08dHLMUOEd/OH1f24qA05K/UUMaeWNC4f5kQRLK4bDnthbO2+jDUF
hOFxk5AbuIrxuq/7swA/hNPaFXRmB+N5YvqfdRFGVH6bsJroKzmQX9AZkvWPSCqUQ67hT/NqzPIE
LWdualZ7rwfdMIN5ZiDTheRrNrXxWn0kzryiWaIKP3qLzl0IlTcacF76PftDJFrRjh6qxsvxJ6xD
xKeJ1IuWpvtBwkk+9WI+b358oC0xOqfrplI8LqfnEV8C9qi5vVxTREbPhcQRx2sgBZ9GWExQnn3m
kwY5PlxRuz4F8Ww+s+eSEvhZg1DZQQK+SgUm8lTGxifnqiUMlcRunXtdW2s1ohDOHXhqUl/lxT4z
jPGqydnHaMyAKAppUMwmpx16TvhuFBs/ifauVp5GIUXnTeqCYMrwywFTtEQmGxkSo/DxeQCKujpH
Ynn89qDXxc/7e9Ju/TrhHIaf726C8pRSPt9lOqeXoi/rO8Ly56w3oSf5rPLReQwAPAsEA5rsROw6
9mdhYQ49U3OiytcVH4phzqKKh6M3IEOcdpxA4ZEQsMMSRu/htg2tIOzdJ/4icwBULC54FB4j+uMR
kTzm4ulwiCnMXcMkr9EtzQJW0g/HoGMSVKnKfxb2KfsoTc4mkdMGP46WEnkedyqWn9H+ft1GLSNd
g5F1WgBNkf2wQeo6r7SX0BzBvA7Yy4rNzRND2ns4Sg2lGx4FKw4V1SJYR0Y5F3YrCRezCSPkrjcq
9V7UH649zI2nEdrFwRRyic59ArmGfVfYiUvaWhx5+/fN/i806GJlqoBO8UFOQfQSvWJuqXl/ipk3
oA4h8mGLh56hv4+Xos6RKNxBe9RFKtvQ8/p8hL4adHWSFUxWgHH+jObJpNWY+vhTXwHs0KcXrtc1
1250fGBXvGNvgI/sGOCpU3xLz9S6EFKJr33oYi0tgoP3zCwOiMCAlgTpylgCViI4gkZxAY7lYkEV
aTZLQ16LP0ws1CWHyiaLlbKiwjZf3Kd2eIUhZ5aVDgQI/R8aSz4ZYeghXHvXaTzWWR4WZiI2CRFj
oTIrO3jjPIl/eXYXwPAClRlDBnDYJ/6IARuCsqBNpVRzeOFoEQ0KQDUt45nwnpPLNrO9hPuW6MQ9
zeoSAS2KVslVHJQLTnXKlUR2603xw1qih/4Q8abVeqc6xz4ikKRSaFj0F8fSziXjf2LdqqU5hOgY
X3X3VY1oXBXjDgGxI4NO2No6/stJeNrzbK87lW5liVLyRgyMq+wFDkYRdqtfMJWxUEJN211I9UGT
fCJTRSC5yB7vsMePM78KL554GUoGvENrUhWx04Illmc7Cxt3rGiEkFspeaXBQTaaZnVEwUO2fGVv
ghuF4sN+oNd6KOShzowdX0d/8bKsC040xmqqJhkMDLcrlCjh00VqLqcb98oRVeqGAsF8Elo7f9Nx
48NSl/+FdF/DyjQKONKGcBLnNovI+kL09JEhFV6txj9uVpSCVEF5NIm1vBzD9cS1FaJoZqv3fXSV
alrjm/IwH1V0Muw/Wot57CWyXmcYqi9ymF1EGXKvSDRcuUtF/NyrecajzrfM1KlRGdUxTWaa0Zn7
B4ahTLBGixjzbQUavBODcCvCRLfqcAMhDznfp3hCZnIp7n95g+ETgUydFEuvo27Yx8eRHWHwf/qj
ED0T/hgl88gHl0mBwUEbwq2gWkJNQLDMH9KOX6r9UadX2gdeCWtVyzLG90hQ8/rl56FlD0K1Xd89
tHJpttpGABqLjOUP0vCqy/ugqb7ezPcUCbWh/nzCZK6K5ggT6kxPW23m8kh5r6LxcvhoMJr8rwIk
eLzhIGYWM5UCHtY09xLqsCMgF00k0h/z0V9t45pUybDmg13yeL0zNeECyLFiFxWg+6jauFRBRl7N
6oTmy5cVKnFzEAXzD3fnGgnS+AAUd4xIP7uVvM9NTIeMIujnHkI6zAMOWQh2J1yZQrBKAQOCRr/J
7P+ZIrf/ptKMfjj6YHbWe/REMb+U3AFjJ7N1ZYQVGVF8Uxcbw0HMiAGkJPI0wOt0PlryMaJMvpKw
kTNgIkefpmrxmb539PAsQbVDpFLEmZol61SvSzulZXkEUISRVlCJQgGXBIRErlJuWA/U6gvxkVrL
HhcpCl0HOHeKjgFhZTiS0ww9bEHKUTmo0fqXP0mgTkYuYm3ideLTfzdJaDb372rbGALuVMK1pLBO
3Z5p6/MrHL6szE82jUZV5Y1NVdh2br044EoVNmYRc0Ldhf+quJYG+55/jF1r5qeCPml05VzEAQR8
RauvPwhqrmq4GJqV+qCGaaaD2b6UZWgyt7pYoTZLS0LHGYxwiN21kdjo9s6OMPbBK6J8NuXJifdR
a8m1DYAraXnpI6dVsEkCCx+fIvU+LcjwXNqaLC5h0bZxAHDuvnH2GyJv2JmU+x935t86PmGHOXpt
zIniwY4Hg2xL2XipB1Lyc5xIC4NVT864PojGGPTYd0IDU2NyCY2eXaLzyQsBrYJHUmklTEgcFxW1
WK5zItV/oEM/nPwtrgRw4qWKa/VXmL0UWPvG7+hRy2TSduWGNU/yPs4afCAn1vaMeA0aw2mNLk5n
JdRVfX9wSJvk0IEly9r4WjXkarUav4bv1mcXu/lM+uXIHJZ5RO5QsWuY9rbl7F/Si/om5ICJ5Xjy
moff0FJTptk1GvnJX/OHacg+cKJwmkxknhxrWSKKsuFSZ5whvb9dB2EY4lHCXyyfEB8jt1jvZz8K
bdVkz1any8on0su3VPoefIHqZxzXXZoT2tkabbqlBlguPHmpNFs/z3MFdor7PF0JTFcwd3kj/3t1
eas47uzQ4wpPkSARJ5ZjWLZ8pIB6FEHk9Y+DDyW2Plwe0aR77W+SK6t2NQKNMEhzzRKUbRJ3xuSM
AWSton9IKbh+gtSuTcGQO6q8eOL6XJnJ6hOleyDIS9kBinPLfnuhcBzibx8jyyEOzUGrQDVMjgRT
yUl+XCGm8ZSbpC2qo8Fvt5Alk91pa5Vw/Vz7TZsXe60ICUOhEw0l48EY52uetbvbWF+/fj/GPiEq
gX5aY6E4Mr4aQ3Xm1Qyr0PXs/+okx5IWMOt3Y6IlLHQIxYDA2o3rN+zqJ1F3xuYnqNkwV3dD7uz3
oGR+aIj2MzWNlkNI9TtIAHkqe/zT+crqVaN6e/8PFejzO5/7DyIAaMl4GKW/d/ytOrWKmls2wTbX
z/BbyC5i7LiOeImc2jAcY4VeLJgMvFjP5xHiZj6iz2Q5s4fYk6KLVntqE/bcMly7aP8mYTbHmRlp
UEQimSNCIj/xjMa+JiQd3eYpQrWkMaox1OeAA6ih1ZFwD3rEZd1t/18vjoEyYhsODg0V8cP17HLw
cnZ8uTNCnkK2fj4UPkhuaYuMRYwdHhnOnvHjyJe2tuW8Yp9F0JaRYEzGqaY9Ow97PvVFW4c9Y88e
egogkm3B2vsQyjZugTf9cpS6HCOJE6LBebdUDFB6FPsWvRjO3GNIJgkuzXjdCCMIk+Zeljn2AHit
KbnaJyxLAj3O0IJ5GDXeHxslF6RcdqDsni2vO6tJrZKQvKILWjJCEPb05XLojeQ04YMn1IZXw3aF
FMYG26Ocms/skkNAZVYWU/DhU595c9WJHVMax0OznVLi/LRuf8tqmz1Gv5+5dAK9JwYlNbgxkAM9
qao2D3enhaseIa1xa7M6vmvU24bxPo7cwOrzcoX6xRrl93CTQgaIaYxbRLkNsQ4IqFaUQRcb2j6B
egNDujLivS7lWrD/2f3F9DRIQOYExCDkArYhpwBrmIDOLayqHLHc5fwQnJRdlZffitZKKvxQYkmu
ZDuBzOugOZqVDNus9245y4jGPdGTuV7xyrAyTeXRUY+4bW/Dmb91UgIw1yOXXTPGdWBdIXqWeLE1
TbuLpvFVAoas62P8RQraz0aIE65Nv4mOglOzqC+a7Aav7+eFNE1EliIhAJOtqEwB/2pNtWuff/xu
nRa4YYuNQBTle7ztBP2znRMmTCEXWwmYJ2O/P8heAyAzT2kzxhZR+D5I+Pkgqh4czvx37bTfLjDX
XkLIiEm0uyfGm1O/kCsrt75352biLnsRQAW4+KOiNv3mY08zI+9YqnbeOSoQyqcOWhOT1P8RXthX
vQSPbEBAFoLxF/XoJtDuX21K4NElnJN5bjj5NZdbxavITJIOPHyQ0u1FM02H4zbf1IL4fOoo13Mp
jVCVo7WE26izKHjoY2xOIn/wO3/S+KXAir58iEWKcnZDtcLVTSXlIsAwJK3yzMcYsXER9uGCRsbe
kE9zbkZebp8WQXLXg40xN2BVOE3Wax0Kjtbe1XDDeFhZQYYZCx3MNuWyzhP3nywvylup/ZZP8hUi
h7yxgb8fkoRr4q9UPPSpHekFvjf9rptM8uZ7TaP2WlGfNFgEutZsgBzeAof/R+C/BirEHpyB2hCN
SNCACtO5nEMskP12cXHVKu+pIkuYlK2tqrkzZ4HH3VvCpAH31C+IovjKUpf/rJ5Hxw/xMs9xrdY3
xlw2psV6Ps7wKRbqasJ8tQHDGOADaYLh16zBQ6iFDcGouRmFYPkKHU6EDVSsOKw5yzpnqQu3DCj1
64Ooetj8Q2a5duoucB95V1lqRI4IPkKcc63FjftS7Gc1GexGjyr4SGWasGQj9sDh3DsKqClGcqeF
PupnPR53Ald9sPMtdVvdz+uwxhmukwWpEtgO+wwpDdESmsuXCS0WmgNPlyXWx3j+5zhZvDG9a9Ze
Z5BYrnouR//mocg+RkU3r1g/ecX2Mpz8vIh1OuE+uKLiTUE9n4dMztzz5LJ2w52IAcbKTLjk/zGD
qD0hJxfB8W5/bB+A/Sl1M0zfEfvT7qW5USczxzJfeOSbOOebT9N67G3+WQJUuVTGDx51E+M9xYqd
MOqH+LahfqGGrXvUPEcTb5XTxRL2auBvqJoM856bB0/Da3oH+ZIAUnOqsmQUtK89RMnypHPiiZZ2
w9qRhac5vO9p4tNRyXns24RBTkdU3gk3A1DG3+byctnm4FEvKS1+LCyIUdAq8CNkjpgHn5wzEipJ
2AyBsGQ8FBnJvfaWxL3vxIjyLXxym7XuUXS1XKz8wNsDVN4EZ5Vg1t0SK0yyCWXiEYPOWWwfWd/P
7c0wem7wSE+24msUUg6ksH6hf0W3hotMQKmSGXafkuV2DNqfwbieZy/fjwYW7BsQ3tlFS7A0mL5G
jROsfBURDJ+sETCPdULJDD5VuHHD75PZLSel4/q9c6VMpjwx6tRPKuw4gxu0yAoPUfSIW5wdPPbK
45FQWYHZM+aq20PGKbVQ1Txet/XaMcvh3YGxz/qtxcKG1LuCK/lfRJH4KxOE/x2WPuaBoGMOUjLv
MXZemKqfAJi48Xg3j6WDbGJ6lGxS1m8skIJJ1L3cEbA00ZwENkxo+iuOCVs+Re4vKHrnjV5xUnE6
RFVBECBCJ9oHREgfsObk/51iqYC5fueCKKE6z1Fo+ycGK2pt0bgEyoOTNaK9ymYj3Bk3GexelQZf
9NXbRbmsqlTR4JrE8IEkKxRrlG1Mg5vNREr7Y9Mhod6o46yCdZQWSh/e7H0rGUOh7Tq7LwxGDxth
ahuB6iQcDMJIVc7a0hw4ibjMaerfXakzfUD8kuOcLBBCp+wxfdIxpy5S/gGZCsY7/BthoUH99bkB
OXI+WFiKnAhPUoJVIrWjmXHZ1uFasqicqaGmQzx4qM8tYjwLIxGJYSwZ5ZeUTLWV3O8wULyVOBa2
4pWpm8VLxmeh3M90dJ09xZi+Xrv51M/Qi79D+HdFaD/yNVkyKedw+Wd+0/3QJ/8EvOWZblzNjBMu
THcdpsL48ofi/RJoAbIWnv9T6vyqri4+W0iOai6lXWuRNDbfWPDm0NefLVsYC2EGAodq5BH4yQLV
tq3EiuJiVoVmvx77xPH1X5vbi88UE62uxFrNq6IIIz9LS2NTW7KBBmTl1IOjz0Qii1gndd+YB8P1
yox7K1KEQr/o27rVMvOq3BMxs2Edp/QpgNY0ZCGWJmbjOY4j9gfkcdf1YYA0dw6cVfY5Ft1qYvyI
Ixpnm+ppbiF1Uzke1R+gbInSwjlmgaT3tDxKTjMx5GXCd9AXI3gk/zkOCG4yXRi12jN81SxuhUSR
eCT9TpPMngRdepEwV242khNJo+tPaeEGJg44TXA4Ms+dTi8YS/JgOE2RwuVnUAiFN1Ycfg2akhp7
Dv2L6qFa22WPu8pZFEhOWF/mfeL2IkA0k6pDPx61hip5Q5tayQ8z0ymzOKGM0SdR4+w0xLRdFhli
KjPrhTqPKJAQ60aiHh/GwW0P5gQldxCnrF4zyhl8TBu+Xw0NigoVwvad396Skguveewl3nV8FUnc
gBytBKSwJzaCeMScRpQaJ35F7C5vn5JMlNXxkvroUF6+KbmFM2u1kKmWMWb3ILHFov1P04uiloq2
zGx/NX8KCcvl4ovGbslK+rRM4kfRhrXg4fdqmTGyealm81Ax2K4/0QetJwC8e3hQ8hPP7+cLOvMS
VQeZsPPBKkEqO7FZKLQZTWzypBToBhDSAXRdKRJkn6SLowVTxkmf8azgQ8eShSBOSTkEZ6kyoOqU
WUQJS4wTqko7/qqpKq838vh9uH6v4CMHakq2hcjPjdcK4RHXwmzN20YQxxFLIIyLVy8GJnLTBTh1
4Tn0pk70bBHRR7/U9Qrduj2SBKS2ogKrxL1CQFgTPOiQPwW4kRM5lESuzcoCfY2i0DvWQupii6Wa
ML6A+xlwKCZX/B5EWqystktJ90+6t9E/XE+8e1epDDacvcRygqPZdkzxI+5bcB/e3dLIgEIkWICx
DTqlQLdVh/DYlBzM54+Y8EUQlQt2ZvDmTbnp+WHockg1W2fEt2TzQgBbNN3AvKyb1mBbEBOdRMPc
MgLDDL0kMwG4AXEaVpGp02gW0P32l1JY2ATgIsTNcI8tSPE7VQhdvW9QKOFaSDUfhj95uFhSeTyM
zTnWTPPS2pguPCyiAraGi9J18DkvcIZIzUsJFnPEivYFdmfyXuF5v02YdeyveCwib3FItJ/twWDV
MH2xjZLbzb5i1BuqE2P4+9NqDKFfSSKiLtJAKHec7+AOfOC2mfiFLtuHCluzN6Shy0BicgWN9qqq
JL+PLELH41tljzbMs+fTIQMNVK4WAfnCw7nNpngUVN4CrbFP7tphstdpOxLdZXEi88VNsxXGORv+
otenbug1rFsiQIUinVQJpvake7LdX3kts7n+ZIk+5JzR9heDZVbuXj/UVZMi3i142m4NX97peOUk
sv3WwmFklctG2gbr8VF+rw5aqVJt+NO2fYO387By0ZO3w87THPH20YfMT8VIPoAtyNmx2Vtz11j4
WWl6GmSdoqnIGHmK9U0xGhvtppOBJ53ClOzS0XWbfhd5NLDiAnj7vdAZefgvPSkSJMwTIRSd567F
l2GSkoZOOLEEuxk9MeBciHTv2R0gMwS916gcPSvv+CGS4zSsCzIOCO743vq+7bPqS6SfJg+qT3mc
g1alHI+cH8pzE/p2cRuHFibqDPHxdPX6VZX/VmZ0ycra2FLq1IY770PAR3PZoI4meA5XAKU6fS1y
9QRDEjprQq4pQhlssjH7NmNKTCfwepJdLdNRVRRGojAfHQo+bJQgj0GN6OOy4jLlAxJsAqHUJFy8
CXcl1FhWlYkNq5k8n25HAObOwlobGhcTRBsRtXRWmJyvnyqtUpYJNxu9PFfRXh/+BntEhL3nQGF0
Vp58Cx6Rg2zlGhxyWeZt0Qo5a0Xq73Yf73OmuWyyb0+R3BC+aavbRsnSDH5N4ubU+Eanoum2v3Ut
QhoNMqALZ/tAB8mOxNObfDmIHur07ixn6I6Lvp2Lp7lV+VMfKntBpT1FIyFeLePW4xU1hReWs83P
Ox5KN+V0SvqDa9PU21UbDOHl2XNReIO071LBEqgGvwI9+SygOtQJSHWjSNPb2ezjV2vp0tBmxZSr
7C0kxJB5PFayXSB3fsgNHqE0nYH1ZT7wBTpQ9VDQtIG1YfLf3E4ZJaJp9vWzB6xQpDRY6aVgmICe
sMJL4pG+wyguuq9RhIsJDctFZjQndB8NJ8g657ehuPxo+eYMvuFaI40peU84dWCAZ2i7/bGJljqP
Bzuff32anOvbsnwsNwUQE3sVhrt8q8GUEK42HYGuchlmkZdjFpkQhq9tSnrMjobGTmlc4vIdEcbe
2/ND6/FupFIKCCgZIGmVzoZBHtv6zzxKbdvHdNgibeZhGDs0A4FE3or2DYDWUEeggSHcv16RGu2V
bvVW5fyCywdPqqagJoO7QBJCJVPF5D5fB+4uw/AyYh83ELFn8GAxI2134V++r12IfJMvXZ8WQpnr
528TqtMBbwEz+GgDGEATy8pHcMkVyvD/7hJwkqVA/eKvi96mUN3wDAUE9GweuEu0YHqhLFmfLwMX
JdlD3518O8szRARQHDHUhYC2zevWzl5OwN5eCkBhUiZaQtWz4jY4ZngcXGGMaJH1XmYpBLU9il9p
1HpzRJxm5/BiGB/ntjvKFnBO9IZS//CAWGy9z7srXwcckb0O7hyY5iW9SCyIkI5gisUmFq1SRnto
pT4uo7CjT7N647+pYHjjNJ4QOahruokB9pD0cUEr/2mMNLTp3Pj3aYWPUO7yifgjk16I9ZbE2vww
fXlu2NROXMX/3ABTQxEmIrf6q0ZP8HR8AAnHXJtzKIxbdI1BKWt6Ax2HlmhBvuPFiul16Gyp+7ye
tTfFrhhDtlJRaTezQm9aJX76GT01vyjTW4FDmgzwLz/eXkve4FyBa+kwZptMcWHx7aib2UvKK46a
D3MGh565/v/gJ6eXqFcMXputzHSS3ZPN19+xIcuptH8ikxFAg9FJa1YG8dB5PBxmApXyKar8ecEl
BSS3E9U4LoGmfiOEA1/tZMMbFP+Sgbc1BRs4gEyN/2AqEENavzNwt3jGDgJqhY3upHp6LdAM6Uvv
dunvNed87HqehHV+pZ5hVy45x3O76YV74S4Ha6aKuTLKtdYcT5TA9cHJsfhMMMSmgPdmBT9ZJkFi
8C739IwXH+7DPBUJeRLxI/lCLM3yNqOPuPwdb+GGQdItLOC3Xix4M8gTsytXptLtmCV1xwktva5K
oe3wg8GnLngD/PSqKu5IDeZ0JgyeJ+pTlVBAvShCl+YqInjtAHn6v3bAVZ5MrsJpkPa354w3trsL
LVr3xvqG/SvDkXIg9wCduOTKm0g6dOKYHBJvR35FDrcfn6+VPEE/W49nPcEiBYt5vkVBaT8+gDGW
36Q5xfSfloxRT8knYDv66+E6hE+IzC6jo09RwHIARIKbJfrIWvOiK63Lg70wTKAOiwxhmnpGDKh+
YUCfEU+DRLg7Xa+/DpfEUzB2KhK0uposlD8jVkjMAxSTfsv6PkyEHi78iOwh8n9oW2iUg5vFErYm
zb9HTTCJ8ZdsOrT578Y7DZPtLZNceOrZ3t08upoa6i0Pd/zXkcaKmM+w2h7L1jYUa4/1iD/H6o//
idtcrynRMdqhs8sFJ/P74ThyFnQa6jIm3CJtVFmiglP0epjySV71MS5+Pwoyt8ceXcKd5eaiWxY2
wCBInVVhykEiVvoHlPQ4yxIdp1QNx4kIhxyXwODozU1Irgfn32PWIMmBaclLvbnP5d+OTEKJnn+6
3YI+FGbbXvL/oDIP2QGyEqhQsgr0lkrIh9bAv0rsR5MlCBWFm2h0X3yxV7U/1A0WFNEwthh1iazR
AU9MJkm3k9TEMu8rkgy0YQhFAkik9rwCU/FeQykEN7DSRgHGZpWJqpNfZehgbU6LJrXNgU8g9ZLI
hk5AanuT31sERspNr5p3MG+9uW8S1FfX/JErilBKZI+pXeoTGesH1k8+yXnlbYUH+0XcY0tFuEKx
0auewFIZWjuMgLAm5cSIKFGHfJg8A1wiZH6ZqdGnkERhQXATNyn5+OEapYRLV7eD1JKLpnNEm/gn
r1Q7MxVO89naJ0N5Wf/hsvw7CNnk/mPvB3f5VQ9JGZzvpB+/D4RZ1lDslZPJZrQvvzhFHOgb8DYz
a3nBX8hp0AqT5m466dLao019DwxANf02oYutg0xkGYt2yUoIAW8hAK95ignzlniXw0TL3mKUpK0r
kSWthulwCad1Oc1fl2YlawFAGNSVbz6L5ql9TJXY/eGfyLFnEiX3IbPgYFJj3yNV4JepHOfSRf5J
hQbhR59NtRjCHsGdYNhLTeYD3h6LDEirO4PnFaDfiFsJ+EVnwpYtMrPnFgC9PYvIBBnnH2dKPhAs
W1612vHLMRl/Va34dpdRQnHjfq4DssyWameUjm7al2QvG8M29jvJ4dMg4bDphdu4RVUIgNa/w6o4
2BerCoGlFAHiQl1bKKE1AipKmYteezbFfJ58SYo9tvYkUXyr1vNcoqjngUo8jnscwwu/m5Um13OM
XyZNxgpOt7empC2QkfFDV7cvS7BkdB7uJNlk+e+PSvk3HTliLakXliqDplEzhphElqgjQ/TbufnZ
a/KTDF7oZuecLPiguiC3PR7ajp6vQwWre3iTgW1A5xrvSulSwQN30OsraAKz42bdymFnL+Hv/kpm
EZD0PGlevRyAiWfeP+0NqJiO3GfI7Pos+4CVjULB5ZrK0eci6/PTmAsI2lgbGjpFnUEGSi5+Yu1p
cA5o2x2fAnXXpitOuHXl6Xkf1VKyiIeMo5n9+ncUX64h2fBVgOPV2KQeePqJoMpjb3383ThEy/s7
/11PdpGalhWMDVsBjibBOOPSID2G3xfvF4Tg6YDnkBDy3EhJkTfpTs0SO1NYRu1D7ABmltquAcrX
LAX6zDvJiECPLMzSgMemr+0G1ri99YIwIPV1zsms7629OA/8eIKO6KfD4xTmk9gM2FN2NQun8slO
96BTZNNKCbILS3X6P7vZmH3ko9lhOUzEDh2+cjLmFntusRIY2UeiFjETpL3pSH5xx/c46u6lzHN/
hTvOdpIYXxSoYCHMHXm+lJ01D3KUN9RYE3zTUzXq7FxZ/iC44FBns+IsV929JDIaF5K3rqK8BW3T
MtLYvCu5fEd/VcC8IURzOXyW6cssWR6mkpIf89vSEL9plFtKQJTJb/80//tRSFdRdj3+vjH+PMcN
tj9J13Eood6cldGRcDG+4YrR66if0YCzBlRxhc//sDH3t1d1P1m2ZRw8xfW40mYB+QW9kaQh7wj5
2M+RVEpEPIk8Bs4zAryCJk1d33kpvjpKi6YSU5zLF+KkgJEZj6Je4ho8ShRk8p18MOxGcqNP3V3T
CHn7EhrmmGucmArelXpN1YZVU4VMspKqfHZ0TjYlQqWMuU4igjfhjgvjCXasqG65i65c5T/4Frfx
blwOAVjVZtjy+ZKBk2h8qXEdjRNLf55ym3q5CWRgGJw0VXD7+6uo4yqTadAMpmnBI5Fkeu8UUEEf
m305thQO0xWp3/R20g2Pw/C/1pORdY0cMv8mF7qbdMS2jlaZmK1KwL64eWIPaMhndPMdC8EiEgIz
hk/V5yhgJchPls8J58CpsOCedxfjkOMWv0N4NF/fKHxqZpPlghzLUNHcPXTtiXQOS/Hx96VIDaGc
rCLGvKT/duGwqc88vUoADLUmUbul47KypubYQRVzBsze75Dr6ZuZkAzGgDlRU0Ek+I+dB9aXS1fn
IzXDkSvJoCuzAItCtfznlp07/VAJ8iUvcFFao1ZLvU5yaYXSRUyI3zzsRPEXfRsidJy+lvs28m00
HPFJLek2C6HdGeK4rf12uCRwxkaCnVPBUip5v/9fnfVQpA6htsvRf+i1tssBtTevgOnhJxDH/wUZ
8EjbMeGhwpkJglqqnUvusC6ZWJqhcyZK0kxZu7AijwGaeM9xfSykB8HCEEUQ4DPIsjf3CfbmM+QT
EoY9HWIZPwL6qVrrTZlfCY1g7bWj8GXtDMQITa+yInM++1NNwswgi6wrmEohicEyWe7C0TfHC4Nk
rA/oEpqN73eEjrkNGS1pJGtbmczXcUkNQ5gW7O6LoR0uwpenPNoKM3Q37vtEzvCwsGNSFmTsJZqW
VY4DN0BncbOHRZR6kDqh948vhxeD4nGkekS6Zx4gdeTBbr1bmVfbFCuFEY7xer+ea4CytBWaehyE
t76lXzFtAJ7lW3rhug4wDI0CslOmKY5idiG3u5qvsxbf+t4DCOnSHWOZZMqAede6qDVHkEN5LhDB
iTkcCRrbjB48u3+OrDo0C4YCcDJWf2De9ItoQwRyulRPyroXJRXq5XIrsEOnEzLJ8FDGCBGDeXah
9dfgwGjS9cC4pUm+IEMng+dVc3QcCAueVBoU0i/c9ZKrGUyXygx1bGHMHAC/Zp6wbTM/+ln+80WN
p9OrQW86J+0Owy8p0s9Pa8UcqgAAS4OsI6ki+Am3bFuvEA5x5y5RlBSI/AXehDwJ2Hwus/NnUhcJ
20F/hxbFJWpLGuat8NMFVhtIjbybtadNqx9U26njMZq7zdbvQYRf8BjcwLE8R/XEyIhPw2ZAzP4W
7bahjgq0DXV5CRGUdYvfsWQgLsXRQoIyrcJ23OzSGph+wqAVFNe0yZsk91JZTzN7qBIqxm/t2IMu
SI5uzG89c/Xu0+HvCVbpgAuY+rg7PxD89kSuBaQoJ9irxn7CDn68Pl86VqLegkccSAKn4LKcFiVi
1kkJUWFTG3HCxwL3S3zd8R6EbZZseI90h2+Ulxm3UgoA/ZZK1LkQWTfItc38RBMdy435eULFGVUU
mK03BS9b0Z0fxqa2qHYB7858YKlbbOXsq+i7B6FUBw6YqBCNDMGxzK3zoRKETB5VL+XvCfH7aIcO
ZksYTImroVEm3ysvwPN7hj0v08aZwUy/pebxv3S/aMLBGePXK2FsjS9lUQOo9Yi3ZfBbo2OYXTyP
2YbZbcsTKZI5WQVKeieCVu1OLNie6jdD+3HILzaFaKDcgob9QrV+o9vwJQJXcmqFsgQntHhqwYHP
iABWejN/Wt7+Bpsya5UplbrMy6GvnxB6O5dgSPIN7AhsnQ1eX6hgxDvRN/s54MkEZvJSYKOtK1o/
MabPTRSAZl3p1tbZkzu5p3e1zzUfozyrjxu3u+8s4lUuOZFXahGPo85LTVRQ8Oc5eKaDKzOmC+xy
e7dpV4dqzZ70dBYVy4yHBwqPS7c7/+rL55HiiNXMpou4bWLYy0DAlSJABrNgtqeiG1iBMLUPDHx+
n5IjdWi62IC7egwEDBwmX+RLNiBNqV5SttCjx4jyuysX6Vtj4aLSf9AmF5XFgQniOOXppMSkOWAJ
BBpVESj36aT0UbfZd4TCXpoZcUfEFl+ii6A7vuhfDGZvjxGi+cGz2nt+TVsG3w4kzy5sPwAVw0BS
BRXSu+3QIxWs7aWfSNzMws7iPb+guAt6XfFnj5SmXF8VY2iIVkteO8qOmNkNGbmcHbhVpkeNKXgO
cu4rtw5Z6GVWwQpm3wcyyWjBG9vAzVhNnbFsLHgLICuXBabWFSAGWfg9R9bbd/zelSYVipDzpoq/
CUD/9UPZzo5Z4FovBYAkBgG8O90rheQ3dl6rOCNUj75+bKLrTsu3KdQjEp94+ZOHd2Q8Niybjvki
0nCpG9kzXxOJD0E53j0Eatg4QMpRgoSfA5IbSH+9CpM867XrfbZWCn1n4sqvtsZthWGpFH09CJXu
NdRK1X+HNMfTTexbFzAs8Ehz7G2p7LGhxETsPKLKMB/1syNajo//wVFLHBQBUTz1ZmEiKpfF7Dwo
WttZLyBtpbZdqeLleGrOXIHG3jRL7csGwFgjHXaSgKiA1g3oEFUSt0ccBo8syEzKDXQrT8sQvd8Q
rzD9onrFyjwX7BypNWYVhIW2oV4zF6NTOCNPt9nRrwb7Roy3Cp+2A/I6DFV7SRWZmFGGIHVFsgvf
gS+UajqeRC4xCLh3A5afGG/iWDjBBLM6R7T47/F25eRJYrtuWZRGRscuFo3RaBe7anfbvxmeJSnR
zTiWlAZJZE/ewWHbrif6AAENuu6ObsqCvtNFA57YdbAtNABeN69lr5MJ4nZ4LQ3hyO7TtRt9slz6
WbwImuIlXVyqTQeksPZcUeOiCU1HoE+SLYQmRASdGcmFGjE+JeE2jrWtYYSgHLwEptN2SWBpxtKZ
ziNshD7dHYBt4SEzUD4PYLFhrepKErw3Bxrbj3Q3GtkKySHHNNKQ7gpESexXZATQxMI7sRH/n578
U3Fbokwa4aodVQ13g4FDA+ACgEqs/2DBN88nKZ9X2P3hdyUT8hXMNPTxPAHIYW95hHB5KQmmQF90
JNO6XxglxS8HakL+c/9hu2l0KBxKJojM09ahRFFrA+YNST0vB6pz9vmyjUyeYaa1O/H2gRwkS2h1
ud1Bq7B3WlEV5iaS9ixyaaKAC5ph8vyE6fP9d6Y5+rUHxiojN8Y+9nwsOYBUVWzeRPZYXVZ9vm6A
aZkfcr/qL7PkIdoYdSvrmKFjj/w2ZpjkpN0t+hKUJC41JZFu3aOEad2TX2kwjr4kcNLLpZvikeYn
aSg5kFHyubgpga8rjExgB+/zCU69N28HFwhby6zArsHP78Cmyn1S/XtFSAaOheO0WkEWFuCa7iE5
0EnTgwia/SkFbJtSgISTAo1+q8G61JtQJTEH3HKpfoNfcX+ete/H3YOW0/0yYh6KKlJFTUeKKT+a
N/WQs/VTX9+0Sy9EEFatKPT1XzNS3UXFJ7ffCpJBc6KA7o28RntAUBlgtUgRisBs4GWIbpb9LvD5
BEb/OP+n4xnRg+GUvkKHnPytqqccAWG2OaVrg+UzlHdxnYm1oUgd+eaukHhLOvdiL6vYLv6fQ7Sh
UkguhGb448JUkMvMFHyl6wLidOU3Vje/e85X/XSgvLcWgU6exe49MvvQylkUExyPlm+rnlUOatFS
xXBIZUp/kRth3lB/hBtImgvsJSnKpHaX+yos2bd5ygiYlogpMB98epU03Da5YGOeKZa9b9jEUQHP
70MFZQO2RqQ+HcKHgu+xltQxX4vP/kjIDzrpn84Hnj25MJjJ7nNrxq+cclax5gHRkcHTrdhi2Q8w
JRWjPpsfI4dmV4aaN8B3UUVuykZlMOwNe9qG4IDnxxYmMN4edCvWp2j5Srwyl8xqn9hzgOhSvRIR
n92rCWJgjXfYDG0U6HSO3YCpiYFC0DNESeXVBmZ0eGBN2LEquSYSAcaYfXyrUNQDgWTg8UYLb8mh
q+A9bcG2Us2FPuZ9B30NEF5NXgS384j47WGykFr/tY0rtagcYC3hIK8idYXIr9zeG4rSgUg8GsgO
z30+tmQvOOLWtGPOWIj+mHhgINvPmwNMQLDWX98URka2huf7PERYEhIL4luZYZMOqoonDzdb+3QZ
f8jexoNhPV6f/tCRJUh5DWT/wopBBbc2WtrolP3scRvXHRqTYQ0VN/fUffXdJnIs1dSos4pyTg5q
OnqE56QRwCvYXsTsntDJ556F0ihh5GJia9cJvljoqVzk1a4Y8boc8AXFhgyS1NUkIfd+qFrZGok9
PDG+EVwGjtCKlGlVToIgNhmTXRiWU8DhMP4DLSEvGQOyrAzPFTiFnreWwdGX/Q+65PsODuLNdR4u
jPTnlGLRBNkDoXwMlgqqkodSQpAs8twe5JR4QrdcSywCUsoB4IbtGyptlZgjhdaCST12pI0px191
dxjxxt+PcR1H1KF8veOX4AOjtaeA6jUFn/n3fHIdr8JcBM7G1krCtNWPXSoJXLo0wdc8ACu/hyim
o5IXC+H2lumpbfeEZKpeGPKxCpKqa1FCVI81tAHAwFxFY+f1AsRhvEE69tvWiP86RYJLHcHdexmf
BRz15oaDbycAJxZSKa+QBTcIeB5TqmarZtb58WS4yyvOOgC1+mlAO18gtpWHGYPBvWVhjlAaJLcj
hehHTh0Z/2qv5pC6eEoBhoFjgOMmK+095mwTPT2rit8HJ4I6ckmzlZsTu9h2LWmRWDMiGRGHmIpu
nBRLfiTc2gBQSowEr/tAfckWtBPKLmr265GTremEBEcNby1DtvmbyJlXtohkLBWYviMt3K38DrjI
pOdRgrglW/kVFTwx4De0Bd0PYOMkPLdbgOYLLz92mC+XC5KxkwkIJNm+2tc4Rq9uNPMISgmNgXnm
4nPLue6lPt9ExKxIiee8J7taflh8Et6LzU5yiuCske8vK4BxngiGC1d6TQC3RnhalCpfRUwfp0c8
PO9DtG4nTKtuQFd1tGufkZJAU1ATM3uXzROOi7Bds527SJEhc6EDerZD/FGWin7IzkabzzK6k7ch
N/eWPxWfec97bRUCc6UMos6Cxp8GP6OCDlSwOaE30J9FTZSx9gvlU6t3E+BmTdK8d6zJJKECmXml
aceTU6VYCBIOCzGDnejVfa+WBRbrUJvWC5aXldruQsAa6LmeC1LSZKiAQWPbi3rigfrJfH2f2RzM
BBvwRv7iJAt53jWEj/jHw1QvlkHafTakdSINhuFYratliTPdxf11u6TpEcQu5SKOMVNOv8m5sLPO
GnllDpng2BvNhuw2TGWNrHZTlRb1nglhkqlPrb5u5MPhlYMMD+mfEQmqFvymctXvANnbYzAr8Hmr
4h6zsyijRrLi88pE5berCslv1cygAxTVc4Vuht2UmiRHlWSo5UQ+tbx020dWo+sqtjAWnoFuxT34
4kGsHxDfpp2uk7/Tov0EEJazSvbCb6cs1vDEEW14LM6vny+5Mzp8tzGkq5ZDVLu+5UsSloro+7nq
jhL6HbPVSPo5FXUa9MXNoO7+2Xzyw/FDXLQzX1stOUNJOplj2qbQuViPbr2ZlzzPGuWdnijLwHTO
5GiVpQyPhtjNi3T+zEEz+UqEjwBGE7GHRBASf53tQTOKzUQTHdJutKzXqjkSJe919wZKukD5KrGb
J11bedeCVoAm1z+Zj/7q+H1ywZwXaE4i/pE5LOS8YrO20v0L1wNF9gzFuhuAE7bzua4n+mU+ybsR
pTu0lsOopenMU8DJTj2Er582ma500N1FA6XSdF0dPjgbjmf5dncH91h3cTlLL+hliDr5p+KEhk4y
eDhPmWLHz/dZAbaj16hUa2CoexQTn22lxKi9aDBaO+HxJjcXV+OE9z1nKKcjVfHPSO6Hlx1mkSAE
x2gqUNqfgWBIqpsExhVR3007esMUyKh13q+qV8jwMV2PiUaOEvq/jlv1/1E15lmoiWcQRtnUoMpV
vUTabMg8yYvdBSNwlRY/r1yCXJe9XHzzY1U8yrMyZmQxgS3Jr0O2i+Hwrpj6U3JfIm9kW6QDvwjN
WCzjcsSAUa/u8ctHOrbVhd93PN2Jv2HaQ2Ym1vGr9e5H+tqRqZuk0zGMyNug1ia2WYbauUzof4f3
oAxS/C6ZYdDXywLu9BORCXkaqBV+S5NiAGAaaYAiYRCHSv7gYyy6MGL7qyKcQ80s/qQiX1n5WtX4
y/dutv0XNiiYOWZ1Pm+J3nqs5Iu75+AS98+NvIZ0ksdSfal0BOsHy6dR3kKX0j1brOw7BNvAXKwS
yg69R5o6ZW0BS71oL9BwJQTfBBj73yCKVhn7GlPeGo4nsevlsVtA1vMEjzZJf1aZEl6VnT0KXb4t
O4kBvc7o008CnPyMQVn+8gL7oewPlryZ28U24ePxl1UR5xH421p6sbx47tqTU20jHjxop44Tspb7
mxnAjuMqFntDF4M61yr3CY7S1JeInA241T2gGdSOhpdrp5uIywwWpqcNFiqPJQjz5fcPTdKHoQsw
4Wr8P42sWGzf2seuNMH8TJI62hqHS1J409h1nzKw/dGhelwX2cg8G6vEiklPBdYt79YU3KPyEiDV
pMGm6ygoFlOjVb+z9Sme/6sR5/xOfQJAKtt77XfThsHyYwathE+u+c/YrJAdDGIBqI8EqqB4qcAE
HQOLATEJOliWpBKaUQaATGxn3Oz2cFjExm0SNV9Azzu1cmDGgf4wXJ3T6hWtv9MThgm4/OsnLkfG
K561PNE6nKnZaALmrTAH/aCChWig5F5pKnTLqORb4lHGs5TYSRh4hD8JZRLwZWo3rMZYsGwrdVFb
ONdaK9knPn1HOiCL5jyiz0qboOGi5wtK7GHY6ZhQGt6SDk4v7lXqytiL86+sWaPyNaib2B2rXlCl
Fv+0oR5FWWgAMrTukN87tVnZw5cDSIlHnzX9+NxO1gH0Dj3gVdo4KtH/oSb/tp9BROp5vW1OMfdJ
xKbjA1Sad4mdUYj3ISG0rhmn8sEydu70C0TM42BlnepHzLgN9z+YCPD/hBAvZegM2V7COFn5b4/k
pf5Emg4aGG/nDU/y5scbQHWdrOT5ABgF8zZ1KL0v0LaHn6yQt1rqt8lyD5LZm3HM95Rb5lRZyo00
gQH9CcObkSWUtUU6iF8bg5pYeCzyTfrm/PROxd1RVVbg8rlme9yOv76EbbCuqYDs5x7XoE39b5df
cx/+hg2Hbf5qviHvKXeVvdvyregx4te11OmMyNU7/yALenXDB2hWfJvuDUpn5CQfdB7HXd6rLJ9X
i8h/IQk/irioUJ5B8aOzHTnZ4SOkW4bG/DAUv4KCfO/zHSw6XNo60+iB3f7paYkWoVklbNUwgsVD
6ZMnNWg+XDvzGhSmAM+Nv4ix8qa7TVCS5xAE2MXRhEdAEzovYd81PHOySJlOBW+6tMZL42ay/iIw
+kvpKoMyV7RNR9nPHUalLrHhU9W9rUdKu/RLydk7zhClEmMYGblKwVzt7K6/Gcr8vYLdnKjMp5xc
0b8sdTNC03Q0bBQhDmRTxIPEhLF7/1yBv5enG2nCgGtlHxE1h+X2sZYJ1ba+JA45vNcKIdzmvIy0
nuhsb+BIsT2oEONwOZsz3I8jMCslFjobSl6I6ctHZsM0WMZV3lyoRgLotcD65lmBtbYNYUU+4Fcr
udNw6xu3AajPU23VDCvhLgrjvybx9yUjnnOKIVmIOa5Wl3O43jFbkSPWLRVLYT5/+zV0F+5NDv6X
AhEWuwuUt7WAO8aCUqVd3LYGqsL5W5pKLGaN1luhqPp/EbIxC4JZgwoPabrHeVmfxWGVMbpv5Yvj
8QpbmRCL5NYo6FHcrGKYtSI+ZI0qE2jGJi8HpUeopGxS7eZorAKu8vlwIOyqn8r1ioRHoeTqn4Ou
UE4+W1ykzckClDrQWkttNGahWVBTAMQbzLqPGCOODcRkx+YTl/cCx33ROOeOPglRuFmZl+KJo+7V
m+yWcWX9kjomaI7FhWDaTFT8E9cT1Uy1JOHa4UQF2Ag68ZytYr2+JKZHh9qGZ1+1ps3xOdxYM6Wu
gfjeKDZxB721zFSEUOaNyOJIBrdnJAsKKtaI/gFpwFt9zG14RT18CDEMgrydGTmBfg62eaifKEDy
SkXz9ODB/5sj9vtyNCNxE+OTjtD63Ewm4CF0fjsMm5FP8goqpi8LsQQvSnzGsFJaAkS2fKmrlcHj
W7Mz99OuqIGu5gPc/4BOabmcF9+pjejD8aKRmWi018sue2itPsX/J3TyhMPbIhSUbz1P281UMvja
3mkZ56JTFfsl41XL03N8WgSnlY8K0apAXN9KvJ9tFAh4oHEeNgE6MLzJ+OEMItQ4XTTaAm2Wi+0l
PVKNOiF1eKramW9IbL8zryszau6V5kcj6oReP/y2gx92L82powOrw7jW18Jz7x1jhTMlorUfH18z
IVsqnNSDfuZ0IuL2dAIrfl7nfy43WAWoHrqYdAIk8oLOkB49RsUdB4AtfQnxcVVuHJ3KTqev3/la
cv+ELUnJwUrP0mgHcQ6JlP+UXbjZ2R2A1gfDBM8GhdXPJUFkul7xAR/u5XZwB6hbHcphukzAjKgX
833fzmgjg9RzWoriRTb/ua7WpfBHNu5MIhWr+pSDALpECaj1qOwjAgcRTlJZqOUhreD3cqGtKFeT
Mh7hZn2oGXNoTbuiJnNJbvvDT4SJOLhGOfKCzaG4GS9bOQ+ZSR0gohVrcW5ptkcVfR1290Jsp6Qb
yB/LQSrbYJd0a63Pbl9sBNPgr8vcDai+ZgRoBLP6C9/py4rR5OMImm6yIqSjeIKi5BAnu4W4aOrK
ycYr8oiLBmQc1iTMpXkI+gy7wa8ThcHQnKIYjjJYL7TlrWx32Z+fu8+aV1Rqo8NnDEkQ/pwG6WyP
kFXpmH87w/mMVwS/ihBQIvmJEmIOI0x2Oda7La4hGwoQB6nMMBdSSU121O0EVOaBSGny5m+atCPt
JzEykTkoXgll4RdeGgdfCoTu3Z2LnMHYHV3wLZ7kP/R+uvT2W5vtOAdz+RcNM/ne3JI+mwSPgdEf
jok2OYoSvPeOcvo6uc4QtNZLryBvlnP6T32lBkmWoEu0G/+tx6BIDukrLgJGptlhZBU/Y7e1+QoA
+N6lY8NBq0UlMeuuL3dupMwqOAieFm6YcV5ZkmLxDTjKRdbM6qHWDmGasYbaAAw11unT/myvYiAC
fm67qM2eywjd2aik76bxXV3+Vw/WQr6S6dmlrseUOSWFyvh/EvkiKm3YTdo50T5FHeCimWpMmVHY
Cw3FstxuNs1akRlVUxVqbhrKz0PLbhKWa0jP8BSs/4DHZ8XNfM2Bhy5aCxO+kddlfR4ZfrgSF6bW
sLSgAeRJ8zH7fEy5UBg3xYlrntwVECIayx+vKj1uzibP1bUYpQCPHHpGqJVwnO1by6kUl4ybi5wi
bK/VUDlTj6/TZVnzJDuSmC+S//PepoZTlpoDjtPrLYI2GjBBaU7HWHCdEAT8OJuOwQqTnVEx2n4J
gFQ0VeJRBgpC9hbp3eWsubDaZVzqimajItoe29C792fnLLXlQT6HQSpCFcN50lEDgcrZo4RdcvKW
rTHv+2FmNpvEh2+BnnycyhOIRlgYjJyMN2Gf4cOLNqAJBo624Um8/Hw7ludlafsVBOPCx8WqjEyu
xhhJsshoKPodBxmtzeymfSnl9lWnOD0Z/zTARR/HkEfzQAu12sblUOkFXbt3PwRWA/VJUXg3sZP+
0UKJw8o9p5+ST58r5s4uC3qTMdlhvEvsS+qhenzA48wVnPTnUfw3lfBm6UWdl2+K/WMGXCmW7Phq
Rp4icBiUqxcQK7Zeeq/NVobq3PKKzLyRP/KgBBxF6LykmZjQ3BfDYM5rQqKX5FO6NnzjEhb1lAuY
PrPBhTjGcz8y1whEwAgSxfQaDh26EUEwDsz4Kf29bBgQ1oVFgEtz06LxDguBqEdVIJhvmGJ42I8M
j6vHbvrqv8XkZUjsGZMDo7neZokJ3N9EsTLjWlgPhlvIpFBbfRl1r+h/DFcl2h+ka4V2s6xTnDM6
cUNPTQAtKPAzmcgi42ClQuIcU+tQ+eoPxwaZjwWjCPdMUfCvYw5eRXDtMP+86C1+r9BYajWJ1MVW
zOvHHzgpdUhnqUdKtWhQuGsMOIxN+8Gw9E4eVe09wNtxXidHFD1Wp5hFqUJWe+caUqyNnXbQjAA/
Vq00r2ljsJUqJLhmgW5G7zeuBkKNtceSEIa2wW9AKYF+mbSPYPkhT6x0y2wxrNb28Jp9NYhc+B80
z9dD/2+widsLJ2njuKWl3Ygs88+DbW1vmiYvqxELEDCypuFbemiqIhP4MHLO0atbLXvThTMMsyn/
CTfQHKtlB7I5QXQYQWoK7Qmm2MB0Kq85raeNBnF+0xugLiRfBb7oyWUokZp2FBDXEDKp5I7m2+eg
sY8eWyP0kvp3hbf3NfJu8H3dd6+m94fpTxRo9wWjIW56RC0syWWHZ/U8nmZMHOTTz5iW9rZ0lUyl
J9MVAj/0Tqt/l9q9qvmOv5vqPvKx521MHa1/PwJMDL0krYcxDTSMX63vDRJZBvlo3n+VLQ7bsslz
lBGpX3CVrlHPs2iCb6YQvlaTqKiDtXwc8gO4K+MrPQUk21KMyLh0s1Q5/d9kHAMFNWwKMltrDttm
vgVijNU5W22pgB1o10yPDOh3p11peHggWniP9abBTg651iF1dpoml1kdchujrmI039PmIz82NQz1
KOjJxacRl61mRXSmgozjAHXVvWzzd3PmyiAZ6BQBGQI3IozayLaqCvRQqgO4bchls4HyJDw1xEkv
HHdPVnV7xeWne1RRhtFuSHAKgNeY/n4yW8/2vvoyOvjdeSjh4bDVu3wSJmMvSWJ8dzFddLufo9vs
yvnpxzJj5ZtluCg7cJY5Uc9qcSlm/6Z4wegGM6UA1LVHSPMp+80Vo4fCKX5WajRmos0zvWwoq2kP
puWG9G+K2zo4STqpcG2AGwPUq1C8kviBR52vvOQ45bQTwQgIdCNyd3QcetVU8x4iyTccnNkvRys4
so+XDLIPywzfech+m+MMd/tN0NC/X+TdsPgoLy9X5SEffR3G9KwSZJsBpPlv+Hf1FU1IzxLb4lc3
uR/b2YAWfMR+BO7XK7w+I6W+RlAzDJdHkRNvG2D4ZQhFIY2WpeVGIQt3Wz7ZHSiAzwyCFQcVyXx7
G5mqLiApBNMS56qAPdPSZw6uGCx0GdSFE4Phi075MOl+YYel5hFKM8/X0Qz/O5BZgEP+rsNlN9n1
SzRI8GmmIdFkolimhaK3nsQS5YPiAv0h5xIo4C5fRavEvB1Q2y8wgHpCT2/IlD8C/Eupy2hB5X2Z
eUs5Aa/GTzZ/sr0d/JkKkgk+4vp/j+GrcEKB47FzUtGM7INii/8M1wbyCYyB2RLGdcA1GdqsOQu5
vafxakNRqpogn6UOPwXs2nevVfEi8nnbriPSzogxzx8Ra34wFUkjiQXnlfZ3oK/zG+QGBToxal6S
vHpDsd9UwqE6lwYAc2HxAjfPvKhNDLyvnRbKamqt59xRHYUQlNtzP1J2+uCZfHA2CIhh0uZ8aoTw
tsRvvIoZ2POTtM+7HuB+dF58Lyn3StOY/kIQw81psVpm2SCMpd4+SUshXX6/3dV9t6xmdpuuZdrj
oUVYpyNqMWp8Gw1lyubwgoW0prZqbhj9Q4gVLCPSkWdQZKlM5Q7rgORYIV0HvOjhTAK0+BhWQKEd
tQfyuDrhx8ibvEOX/7IiE6fa74yolg5yuMpFCbohnJyfzw+7lKjO1JlskFy/wQwlHTMBmTgsYPuv
D+ZZqNnsfZUdGmq0bfuvDU9ya7JzeVFgUyfng6RdEFe87PQGbCF2vjHdlji/EwjEV+txuULNqoWk
v6YwcBHbUeBShMGq1F8K09GmB+Q4nVk68tJLoLa8YthKaswGctvJJ1DNb5OWf9Sa5yvLj8uZgpqo
neEKAe7xjmXv4AiWy5GZpNU0y4LNzlE8Bw+R4al90oR35zKQHey38Rl0SIy8EDeIYnLibdwOC5oN
JG23cqlnneMahfM0YLQnEoROtOfhGDBE6qAelAtuG48ziEDCOmq9wy/q4fuLg9+MmLgKQ/R2VFFq
LxQbUH4tzOhpIqE/HP5g6IYigkJXvlmRNexAfT09cCp4i8bDTXzQAarApy29rKBj83i4uDAyYK5M
j7Zp336JrKFvVm/d7oZWHtpafUWtkG6k+8F3Pwu4m6C+KEp9UJ552z+FB/MKknBQGYNsXBkKWq+i
6KXTqnjVmG+rWnB9rLRCcPYSgtqOQgpuctKzwslNrsu2N5ToJKmW/EHs5x6UgiormqGVrRvyHz8j
bTzGrnhUQvrB6W86pT6tGGNSiulHWoJN3RI1tlaQ8OplxHEWWy1JqOKqV4Sw1Gy4BkWvhfdelzsg
ckjFuiu7U99SzLwnM+VETrjqd3Zfe/2Ik5OqUADTxCGTplwg5JtALxst0iJuf/cxva92UBoYTXQC
OY7/Oe3Chj68gIff8Rk4V/IE2tLKOS3RIlROZG6L7B7A+o1s3H+nFAz05SZAIbygGfAhNnsJlufn
H4C5IySqeVGj8afcuy5khds6Sr/aY3Zd9ifQ/fS7yaEbX91rqIdO47Hn4VtnwCGl5VEaCPXASH/9
jMe8cS0+GAI69PG3II/z/8oJjfqPuzYtKyiutRZQsgQC4LVZpDH8omvrX9BHykXivU3hFCZM6OMB
ebLRXbP/F+Lk860wHnis8fp0QCmjoBsIjx2nEkpmQPGnMgi+nawc6VugjvgOazxpUXdo4938S8gy
eFeqFBtmhk6ntb7p3C3Yl34QgYumW9NcIkublxej8bza/ht6LcBHYqPqlU1g0ujI0HKTyIPDmh1y
W/jomJHxJBrfijNly5DB4CAaGzKBmQiflywJZLICbfHuxhJR6OfTwRdEZtxLcSgSi2zZcvSp0MPu
TGGMCuZOyLQnP1tyAWlRZbsYRDbO3thoQsTKM9jm2oUnEsCklFLoPQ71fvK0pPbeFO9GE5khHO7V
u8C8BxxkZFeZCRWdH8A06HVrhx/BZzaORfbrfRiqfxBFHtO6s+nFCwDNptpRzZ7kXkqjY1WzmTEf
ltcq0xu+P1hFNVqZrx4gkxuAj670Qtb8kHs5jO1I/tNUxuNJC8ZNvznY7Ttu0ZHmzFrkJAG/AHvy
RKonAdkuWuEG50suqCWe+aGWxaK1tb/cYXlCeVhuUaZgvTL7kTuOg/93OHu8TrUdkPJljHGDvbO9
k3Rb7Q/REI8p8ZpsRiUCBNUyQI7oo3mFVO2rQW9/vKyD56lEkCh2kXvhfH+UV5akCv7qQj15l464
P98YN0grM3FEEUSlYQmCd2/Y51/VJ/rvOglbAsFUQvPwQiNVUsiHMLIGzAM6tRvJY120M0tcmCc/
hXmd+E3j5+IQtwui9ThFac7n0OJLvvnSZTDSrmw6oHPxnBmN2ThjGVcICKRlKfyQ9W7/wKnHo26y
hl+gqOu/075WEIJ6T367cxpeDEHc7Py2lh0IdO6UOD5poPGkNuQBT/W2znJSzvId7cGlI0sSjWVR
WivuD9Huox6F3QXaa15yTglW6ahVcSz63Gp79tOdhKgV3AwQeU4nttKsPglUfZQNmLwkcbhMm00p
0T9+s4A0YL9Hatr/84uJj5EcqOmnC2KJnkE0Quy8PBsHNqhFY89cXiFurL9qgGvH8F6QlJQKH7Pc
YpXZ0NvgM67okNFhI+i5CRxpAlonANGTEij18+Jaog0MtCwYOiVz5T4+KeeZYPQQPKPXNqQvMnmi
N/n/VTgFbPhbjFUt/ebz+ats1Jb604SlmjeACF+fXsHnblirq8TqPMr4DUsIK3IlNAlXdxiC2+uJ
hWvr+9MrfrNzL7looIzlz/KI9lskWgREzdd3RNP6FG7AwXrWjbbNaPiUZQ7hqEWv5OO+dof/myuf
7N01FCfBmtDxT9XczSwQ8HW4YuBRNH4SRFb3zsdZhCUgzahipJJS96GJvO7PV732QgmjeetrAT3n
+kcsVUoSJYdl2rlLALUeXiUabAF0ItykjbdLftTx9oHFYdX856Kps6zffYI2hHVUrKjSkOXdGX9o
0JcJUp1elMwFqiUKhwR6/fEvHITnC0HRn21eC3VTx9Olgx4lvulAJJmYC+bZ7jz7FIVDqUBZgJ8p
vXjw7icDKnRJULjCGurZflZK/TsAJDHMwoFPKWXfZJM+1O7hj3cpJNCBiB2EzM/DvORbYPBVf7Vg
nDAQf4adisHw0vmLcT0DUdx147H4NXeL8npPRv4vGuJxeH32hIFiq1PtWf3pMTq6QkwLZ5DDY3Kd
i99ivNe9Z3+JMUrleMBn3WDehPkoEwuvNmxvxI205KCIDWi0fKp2NMvlK7tEgMX0TYrO7lVix68+
pa5xvSXiKUUmj1gd9OlOlPJo74UEASYoaAkRSvjDmd/1Ks4CWxnseMhLe7U5FGm+nFs95vlGh6Kl
84Bsq+rcA5BHVWIuivbr6NIQMjEx8kgZp61/6tTTXvMg1q2hb38/ONNX25UXWhLP8GKKpzQ8nslx
4UCCJef7OA18jVvl1RXXbQa+y0SyRzC5Gl4Qpg7Rp4DkBDVpnSYTQgMBiLUXjdkWuksIZs4e8M4O
GTac1nwamBV/Pb3WJqSs8vB1wl0PaIgzC/iquiuxGkTXoq47wzndms3Obx+wqHE1i/CtF9Wg9ftr
3Y/EQtH7JbL9jZ2K8ex36ERPFU5n3n6OdPHnFTJe1mSagHvFSBEaVxcMknvLseIwSP8iVVaH47dx
cMf6+YBQeSkusiEPkUvBErmMC2EVLz1Aw4ta4Cdx6CCnp8V6S7MBw2SxMPLeLS3xzE3V/5bjkHUL
vACdGS3W+Uk7BKE3ccInEMSRq2d3wPcAD9rq1RQgQnNgzEAYp6Ch5cuW6wsaVio17dr1s7FnEKaC
Pfa9axF4Yf4zpjxJnu5GnAUTBw1elriKtK3Ow9rwyhlLF2exr4wDbghZztjzSchkCev1o4vCe5Fg
p+0Eu0SpXaZfmS2k0a84sZqVSTutLBaMMVGq+dbUwvIVwlKfTL0H/3F3uuV8BlzJgUTDhYx1phDO
ww/N9IKdr7s0Kk14EFJUyWSZgu1QWi9qr12KqzCgZ2+aafvlEgrulCFUCXWoMmOrBNK0mHuj6sMe
OxWe/nWofpCaYXr3++HJYtgY1bM3Xc3Vz0DgSL3/UN2GM2R8FQHsJhODCzDcG2pZaw1rJt5ckupS
TKN64++g/fT2pVJPjCAnaOPJ9106sYqQaHCqpzgpmZbr3POkKdctWSe0WV9+IAcouEgAoMc6kXvs
dKsI9iLhFR9XQIgiGYntv+vQJ5Ue4akpxD+H5meJRm2+hW/NTEsoGBQVfjl/BHk7xuhqSBnUqIY0
0gXsT2eD1tBBzGjwctpaj3LCgRHI/LolvMuCZ3pCS+sScGAFsVe34LoQABNKoWPIH833xtlDmuNO
zLHtLM6zPIjaSCgZIm3+WErqgNyNPsr8/M6k5WmCOmyCPzQyiljK9nMJlyFD/2qtFMzqZBbWaAvy
pOTS20GpmYwYW3yKY/HNzTVNdWpWFqTW2vzooZmgvhHEB2TGdyG5rtZnx4eFK6CivFwpY+8321do
MesLFl6oPqTgYQ/UCuk/MGMkc79rbk83dAhvMXkzF9WVRzyeAnH/KbdLjBeJCqUcUNUhKxf4rM7F
JvZ//7XELkFeGCUS2xeLYs0rfurLniH+9tKlgwc1tr/+y7LwvO7Tgu3nr6A0StwkGhVBy/mDO9dO
iNJi+ghRugTkh0antmccjLxs7kDyj/Wl7CHLXBSlDVex+Oe+ea0l6nVcsKXFnJ/EJ++dB8tFrzFJ
MfxD2xHGZG/DPR/PajzVNZEOvbpJ+puQACNZy62QFHAxUs9anaCz1BTcoUsCgyVnJeCPYQP+YHPU
d/Q9H+En83E1qkVUtlYigAyNLi1gBEBw1XIewnxxWL80jeidEps94kZ4YoOTS7ZfsGQL9H/YTkH7
2SP3+lL1Sng2RJ2nSnvTYHpQftOAW+UFx06hMrlhQdzxvZtSh1H2EinpOePZCGo+o1LDlEd0DOxK
bdugaSVH/DiLc6VsWhLkiNDIGJDSmU1dsIoTjxS1h5+IhBi4Bu4gAQoEUWo/zuRdncQsM9EAH9ra
KJOn/aF/UrzGbgSXH6eRpDNT8sFxujc4ZRadKgmP76B9NGS0GkdQU7k4KXUhNdorrLJIUuy5/Adc
XtJSbb1uvRSWIqH+dzoqK6EA9V+xbbC5qIWuzgnFsGP/UJnqjWvyqJ0L+pBgIMQxEAO2dnwb45q2
WVFMsctGKwEgtsbTKWhUQCWOiVKeX4Nh6i0DyKZl9qvNbVNaa9GcBqQtD50o/cJAVH1mnIKxU+NJ
0piEoqQ8/Q/+/WWiqt/HRfUG0O5SmUyHlYB7XM5hST9Adjc/gGFRver9CWmw1w7AhKMgCVzhfzRB
+DmVvcOgpPR0bqx3v3yBxp8JxSiZZpgyZ+m867p1o9HS1n8tdmlTUbCVb76T+DQyVmr6SVggwudt
xQOOctV2Abi02F/Y503iUBts8pc1gBzzoagbS5fMlsZOm67ff7a5KrXk4ENR9w5ahrwj2vPSbiRY
ismvnlIK6ahKTf/Ro2tJNMS4trST8zXIT1wxhz+VmA5ENPLNk3obnSIffTVYkzWmgE05neNGCtOC
VvaJz2pbeuSqf9QAOgnQpUBqJ550V9MywgQQAPwMx8EBuPvJ6D1ga5Nv8KYZ8I6Re9JqRwK+gdnU
3H2cv0/OJQA9qdVU5pVA3Ow8Dnf/Hafu+a+vc9MjrOuww2AxDBOWX6Xm1Qd/SiA/4m4XEmhvgJUL
6YD/3RiaA6SYoDSe4E0tt2sarS0ygyWk4sOcQ1i7OmiHKMfyPq/maRzbcDSwgfHNX41/0wBoKc8A
tyNEPFwk7T1y43nAizr+HpyMc29RwKzJoG65b6KCHdxWLt8pnpF4uTsUfU/3OokASeCgVsXTCaYg
1NbwAkS0k2rEwTB9GOfqZbJI+M/cb6Qc5yomxbnPgnW0cVrOY2/JB5RjZDHAOPV9vQt1+B6nAaJG
TLX77fmiwbT/yKj427rtjmshTAtQj/YLt00uLeZTDvn3q3qtPGx+m8XyttG6oq9ERjnR+14Timul
NVsDdd1dutclFvw7npENVwQziQTJlJbb4P1zCTp7y0IKqhG+2UJ9j9xtvHjTFx6X0MKTjhhZJEFJ
DcIHYw/w8jZMoNSDkTqAlhVIlWLK6Q165aajO06Tw9UIXhHTjm/5HjYn9LjPMN0XY8g98yTMobIA
1z9ftGGIQgCrdMHVVfJCD7KECV+eV9xkAYA7httGL4naGmlSaza1yA3MTR42YGf8gGhfhn1wW8WF
UAuYJyJzMmYgq5OKSzXTzdHngW+FFpWQ4gGDhtpwHPSDeH77EBJb3dZQtWyxkfK6wGM1YU7NYmOp
XC0u457sZfp+OM4RlVhsoiTFzl196ymulDJubUN84gUsdpSNL9jPD6n0JZ4ErPvRAd2xOpKCwxFm
aeIE40Qgh+8sX8ka6gdIE/JhU7++MsYpqX0rZu0mnByx2SVfTCQq7gwMJMcJpRWEEPO2ZbFTNyuW
y72aYDdyOunwf29+twGIJIWWNCwKbt8B6ZlHsxw/NGD/injzIxuyg1l6PTVO7hYw9PNWdLx4IKc0
0q6wRafTgH9BwHVlTe9ih+2CxO0VFx9VUoOc3DZQkjd2eMc1VpzgmGAWgA3sZI5HHXEtFgDodEHg
Ax0iMUVWrNKdCtL5Vufdcqrls8JJjmLzVwYkjrU5w2UCWFExUVR0ewU2kjHLF/k4gPY3hEVBF3JD
2UMyyA94f//bU/T7cuNTkY/I5xXah8qXSr0oM1cpAP5pHlTyRQVcWo6WkJVTPw9tp1bap7DbHa0c
45Bi9CjhVijeRsQgsiFdvWWLV4cbh4wDSsV5ldF1lIzaRQQabBrWCkVxsT+TTPvmPub34+QuEpwe
JPb33ljlZGTzMeLWb/QEiN7E6hYN0doL9u1O0MhecAvSbypPZVgHGvZUJu7TJgnt/5+ClpA/8i/u
B01s78nVKNGaByJrLtBSszKcO+Xr3GdlPN+Y1VzzIRX4h7E0UyMtDwgC3PInasJcB81nw+fP3VAk
8oixm+nhl0N1GPnbWd5+s6Dq+bt7bJUjvCEsRM2SXufKsj/d1AdTQS2PY7DX1C1/sY945RGusL1W
XM8bu18Q4kZm5s4vBBM6z41oU2RQrqBQmrPB9nwLd8Yno6CAADnk7Dx3Fbp+PcftSjyv36VblJ8l
eiSJvGox3ZXiYgPbIz8VhrYHijbt3t3dl02ideBBiUfyuPdsz+qyINlTZ9OlTKEACSToPa1UU6r0
KrYNOb4RFwVawldXrkN3l1jbOSPJtTf7WbW3sJYmutbkGvuMlvvJyUlXZDRML5alccJIr9jYDYkx
Nt/lecnQe8o3dwX2cjqXzu8JwutEVAO65HeYMAQqFi4PAS6HIBFZ3n+6/m5KXM0US45MhsLrds92
It0+z76njwOw6QhCAQy3a3vdoh50XPMxSTnGsVJVcvickAXi5kq6WAqMMA2DeTbxC/QS1xvlcKBF
ONIuBZTRMedOIYIW3fv2WVY+kJFT6Htj82z1V9gCcZYo+jwMHnABjr2DOMM1XXcNzcSmdzf1GC81
t7CuC9TQjk1TBODOpyiYAwaRBvRmZrE5fg1//LMRxfBXfAFDDYiGyfuwtxSsseamVhOOLpGm03mt
+o+eX7h9dquWJT8rJQ7LOr8YgS6RFtPor/bexs18do6OciZ3ApN+T/klvPbVsAWq2W24dMsb1dlY
cLCwNSlMPRQDi3yTjGJElYVtGoNlRpcExN5DpuEBU935ItSYtunnHDlUrZwePBFXCZ7t/je5q+yc
Egk/JX2nuNkmtLl19x2//eVKrgcUNvSlSIO1b2p6PpqAg15iGxAHVjdrvhh521vFIlMMuhN+tFc0
2jT3BW1+jiFd1cxcaBAQabKYULGGWcCTrVaur7fGXkajFf4TENLpxx1Xh4ENGdbREuG13EXK9UJ1
suTwzqFhhcznuFW/PRefvi4Ie1ADFFp73oLLcHxSXaswaAHJQtlYHxXzWEEA/DnGhqvErgiEAINa
EbEKMt7tjwOibAU6vlsUqmuPB6skGXUmeVYPNKyi7OSaAggfu8guGEf5XO7sYaDPW3UWCVLomZWz
3tLRxO8nFqwItdSPMYZXtT7MPUrojV5i5xglrG3G6X71NYRi19kyA2XIkzcwqsj2Vflvfrd+HWHP
M/de04apQuYXsXaQw93eRQw1GUlSOzkPjXaLSwYDm91fqR0jn0KCm6XZ7uwcoMxYHJO3GXmHKsVc
xlMTxqJshTppCHsq243kylI0QTtNNX7yTZXoXmbqeHBafRRmtcI+3aR8e0VJ5nwl9HcrMFyspi1Y
i4551LOsLmBkGld/QSIr1uxdR/fOmerHNkgyqWwp039Fwl4Spctsv6bbog1ANTgGfptRRz3RCbLi
gtthjJtGOS3OKI7AzEDHjYDBI3q8CViSAsPGNSSJ5WxjZyE4Vk+wwGvKK1Q8r2GTl8+8QGzZxXqE
9Uf0awzy547MXoW7Vrjx23x4Rxqh1csXiQVqqjVMeTXnfnNhazAKadP/qzpq/5V8Yj9EAY7N/5gs
+Klqnha4qogWAxH1f3RqD/JhpsCRX/K/IHQq4FHQwDIdSIjx0HrSIscXKpZeXCdbZxbM0jhg+q6B
qLFkcRhhDr0HR2VRoFuS2WT1TRdJ4ePV/wkiAu3FRi/2VkZy2A2XJpFLkUeorZUJxuOzjB53UkfF
d3gvUMNFIUlLQKapR69hVpoZoKlbfqPeC1eC94coDe4pSHBPhAhwsxdai/KAiAWouTD3MQjtz67C
2qzfiKgMOVuzIVdNdlL+Z8EV/bz0xZ6SSli2rEyDsLftZsoWnOzBEOt0xrM3vPkU7Uhfy2T6A9o9
1enrgA0YjLqGJMfkErefXZRpxWcZ2u3TWt3kNIHRbYJmKxs6/NwWu5b8gK0QFehRhqChzdu2GixB
x96sPNs0G9muWCftG51GUmK9/jvGfKbfqfnbmyXO8XP3Ev6x6AJ3H1TnSEOhZIZF0dN8bJsOL+B7
uS6OVJYiVtQ+ig6Hm02QqX3vF0e61bGcHZcTWGnylW2xG6zCugKt09v42Vllq+1Q+gVcK4bqMiCQ
idTz/fnGK7d8nndWzNKufq1MQJU9V7DXmwjHi+z7YYmEcEj8LXIxzgoFmb9pj1+Ywcv9x7Q8XyL5
luWmUV7qk9ovrHM9qqGGgiK07ardBlVng1+9nrnvvk/APTaMTAvL2lL1xMtPXfMqWRbT4PIIbG30
j+T3gOLdGb3Yb7eK8kqEscd1dK+fgae8GCc1R5++NFzAy3zidsQirlDVXbZOkkP1N0yi0dBVKZg2
fkU8LCZY99AxFLqFXlpWtJiWfOFwRITs0Q/u9iSQB0OeXhnzroV3EIjvJ1gwtSwWabfz/1vdW9GZ
g7kmYU5lFnztPaaKNC7Hv6oEMB3obZUPSQV/5d1/zUgoBXNPFR+Pvsd+aBjndDcOzue09wz9XlSp
iIZKJJGa7qFu71SFuLxPmbsAjRbWk2ofxBfag1s0vlJxJZ3h460GE8m9HjQWXvYMpKy8yulL03kM
x3KpNtEvm3i0cvdYXLSX1I50oxjWP7C63n8CUo3X5sD4zKI2zqgzxkEeBAlkhcAmjkbHz7KIj2KS
5KXOQudgddMM/LEVBGkVgjnDlOSAbvDg9Mi/PRl47Rtyix2R/o+eKvP2KbF7ZIU/sjbU95J0qQL/
QDvD9HDrq7/Fm8WvRlAoiGhBF3zcPdMOd6ZeubiuxwhMYJNge0Vfr1GQQW/qorSfaMzb2miqBEhQ
kATQc6vumikNQ/Fkns0BaNgwt+QfCiSEUZCtbSvhsulN9BBG28bGxsNCqXrc4DfhkV9bHtZPRzP9
JzNDCnkDQ3H5kun8H+DsUDmIxKdOmbN0c5DmA098tM8gy3jQGWIf+sA1zxiw+xzYagPl5/Wv/Xtn
aq9cPj01KnfQEh49sO+SyrbcWfiuAUeIN9N9Vsn8j9/aImSU8740v7MBnWPOFdMGCTQMlnKovPfX
V7JucjeAS309ND6WERIfmm+ijBhSEWoM+2L4fIBMzecCvfTJ9XnomRXhFk3UrNKQcfPL5zxsXQtt
J3jyg92l5fAYdtNEQ8QAV682q+mI8TYuDGGnfnnn2eK6A71cDu9XxZ5R0inr1/tJQneBYj82gdRQ
HKGNIzW8NaaiBFHWWd4n2oq8uUzCiMPrJCgPXSDrf8DTRirAPQ9Y0GmCuFn+KSkF2RUP6cgS0jmy
hXUfiG+PEFonW7IPm1E81jc/ON2m+xUTCiukprznbUXDZZXBu+gWdeRWqpucRj70GwJI8D4UU+MW
15wKNOmp1vITYJRbnMMpMMMMjpw7tO39/z+cIHjpgypR8LRHSujmeZ6thuVv4Ru+wZE9m7rw9SAf
b6oIdW/8YxR/uCTb8JsvLa5mDTpugsAZjBzk+SFcKAC9+hgwBc7RNoXSGZCfojEIDuSMfSJmT9AG
kY6UYb00G8mJqv5RyKo3wU31AiF7UHRmGtLtZ7lIBuVqu81H0MsIGZZgRO2qzubtfBlRbfGSbA74
wqO9PXYteSyxKPSyzbb7S4jyutKSK4DGZPlp7M1BFSHpMHHCt2Xz4AMrO/RSFQT3sBwpZi5cZc06
eab/cyPFFqHhRIBVCqd9bwRMXU2Ov4E+RVa5u2ICbnHbRtMv7/n+dMK6UYMpMXaMv3k9qGpEX9YS
zezJlLSwYr2GO2fcMU5xESxlWDscD3RGjivLCG7lFGf/hw7z8KZ5zmMaZ03i3fmx2XO9lm6+GYzX
zyibAypAWg9waqdc+8A4toXyfk0BFgVJE9zgbympQjGEN6w+B26bccRzQJbk7hUCYUoJFj2vYVNn
51u2eRhyiAM5hiA4vIU5NfNw3OBnTCCzGkozRBLL2u9uD+dmCe2f2ZregbciCYHFTFnUV/0WySfY
PnOi2rSgPemhg2L/Ekzn/f7naZHGXQcH7MLYRKgaCGsDZHflOnlx1JrDHW22ZiqJojV64gFlsGjS
krwLMFnz/CG1BVT6hRsNRIinq0QhhztT2GNaoIchcY6eVq9loY0sBbyJ09kqZUt63VRAhn2FBch/
z40uAuO4dmMwIQhZCOBWPO/kNZXS9n5BepaYpCkC9MBCKFGPH9ZW39x4szxMpCKsAweOdHApy75r
j8O6lASX/6FugVKxtzPBVGVn0tlVaOu29w5WWRAhQme9aPczHK7ZMA8/QQLFzg86B40JwXTbXJrT
n0drjFV2exyLKvsSFSOfveN44HlckwzfdZTp6y1A3lpdDvd+kJNXFdN94QN1diEdE2aoI6wRDjVG
R47dpmdCmmD6/1Mn6XwNLmCAalYlRfqZyiBLkIDjVjDFgny32b5+dTEHRwIwn0AjXniNlfwZm8Fg
cZ4Cbe3q2FxBPO0FrC+Ld25XOrwFtYWWD4mDDoHlLDo2bc1vU8cBLrHfmuNg8cKAm2rTTGS+x7po
RCajvY1a3pn18WXRiozrVLksAERGje6xwp2o+LXWuOyv5k62NrGH3gXpkmhM4Lm8R6wD8fiE7lPj
AX7pDW8ZDpFGST8r59rvszWXGYBkM7LhvY2Go/jTHUSEMi8HYCUrJq85NpPGmkiZavr7LVlitFxn
XrwSzVLyIz7qsvJETNiJJZATVhis9ZugLDFufqjwI0/wmpGpxHxVx16R2U4x3K2UzpS1KKSEI16m
VH0chfVMcxLZjpgZU/mPbehp0MIWLNdwxbZqVGCWPSPNtp0Lo8lk10zoBvx7hKfu+6M+yHjSQ2/0
6ijPpBVNPVe+iCFf3rRpJEZNOKsUwU60M7G5EInxAHjLLiEuhnoVy5mHz9P1q73AjOFB92/xCrW/
A7X96yfw/TzuGoFtHg+Y4CX8Cn2kf12bWcdxIc1BuHfo8N5l18vFrgLisZ69zsGNyEQB5lkFTCQO
H7BEANg9Re9bcbW4QWUN38WMIJkhm8XRleGx/OEazYRcdWevigASmpVLm/Kos96Yfro47qOb7pwT
HELRR6EEyiIG3H45DVuhkrvQIs7nUnjStaMDsve5fIeEiy5qwWhWzPFtamKYmzCVTzGD/Z0sR3Lj
SVQ7eie4ArH6c9lxA90yscJqfySyVBc3L//+yYYsA7ZFZSVqt/Qe+Nygl1nTOIAu50oWzGQTzi/o
HPt7r50xc4E0fvJPJvufq/9RCnGb5cuIBXX/8xw1juGTXN0YvfvcHVHfXrHf2qoTjWosPbRhG10+
xEZP216ygFX4GoA6bLrK3Ic0UgABPoj0iCYltgxJ41/PHan7I91TFk0su2uqZkX/6GvB74nWH42Z
x1TruaOOTmE4Hav6Gm8ViZyjWhL0MioQ2lZRZmyzrLUFJT6s02MPhFn+WSyu7x2LHgnjfP5XvZeO
lOoOA9049czukgPLBeq58f6ot4E0HyrJ3eYZ8qetQDg1l0dR15mCm6aJNpjynYmSAvTHBw4K7L8c
dkl2R+GqbaQBrMXi+NqHNfh9IlnN9+SnTVU5BQ5ODZO4atix3Cy7bAlfsP6EEPC5zqsXJ4RFeWMT
BpS+33QksIEDNTjWr0Va/n+p0NdDV0fFCzncFChixFocKmF1hw/Cbpkg1nK46Cpj7k6vN/bwulTt
rVH6nhdSEYirmoVpVft9b/ESAhgTHudloRjIU/tJ907nt7vutdbNXxzlzShT1zzOfSvD5m9zr6uX
AldGm/lBcKLg1mdkx5xI57sUJo1Iz1YIb9W2zd93X0QWNbVV4c7IieOnddAuQGOutkVgn5u38Qyq
/hvh0H5MOG/J2pigckzod8OUKRLzMPX1dFaIBThexVF3kPDpqjsHBRFqDykCV3k4uzuj3kJVIQFw
f5eI6e0vt9kb/i9UOLGGz8di4K7MIpUrfTNsGUTvf7/wZRmdvTJu1Y2XniUycnPNgH177CxNzyLD
kmq5bJvxJjPQelWW+w4djuq0e1Sn/DR3pMH/63/aISJeUEbUtpRVbJ6Kt4o5Ln1BJiD44itXrtUF
gSnZha77mMzTf5qtYJByBVMQP2xQy0MqlaA2K1pAK6pGfY3RxbFgmSGCXCTk54EwUhZHz5rB9lFp
OhxZ2WytDHv+BmfFtSC6QwP0rY+URc7zYAomj2oPERBTE8QK342WEMm7Rw9tLlLuoEfFZqHB9VUe
8t9WfxzGKhbzjMCfmFTNm7qc5wEI0VZywFW44+1gZLqYzjkXzb1pA66TfQ3yELtHHKmjY0x609Pa
gqBCGFhLkxZMva+5TcGsM8jM4kdarCR+RLXSzFVS9pUJhfaNMUyUSLPbNTbsfbv2/33kU0TbsNEp
Th6IRK1+k8qHxOfhcpfJl6lIs0EhVRYWQ481agogcm22XbUo4u80pczySDv4fhsWLYLYrxxaGMEo
CrHHAtviMugEEh+6Wh0pyXzTOr23NQrwcNxuhPogphgABw2xtHJeP3uqacXnla/Z/xnVCOyK802B
fal4plr5WT0RvESpo3O/4dpi+5cv1/5hkcZobSSBG8DJyZ4Moyd19TTUAsApTNF9USA/skMEEJy0
aLu3XEazOcbTNFV1idC/OKmly15pYsiSze6lLU1ZXvTCMt0xzl75vPzFj+DPvJVDxmme6QdDjnpC
HPlcbp3zBjJhS8BLfBHsNStzLuTQZElq8+6rGBpG3iJ/KT1w1ruNLq2Pq89VZ+KNczK5IaLzEh31
QZU7s9L8aysgvzyijBBxJno7hfq3OnSjEphx7bM0z7PlGzPSjoo391u5etaboUPh9kz0Kh2m5fMx
QwjZyLErgCz2FLXIi4nL29R2TaJm/Jal/HYot+wU4w6Q0QGt5RFTs6jqyKBxy0G1kHB8pogxCEBX
saVqLiATWsEZqK1QOoHLstioLxB/lIqvpQzYhSZYzVhqTcivT+DrBwmTOlX1fU3pkBi8SXGuHTc1
mjqpRzk5oQNb4TwqlJk7DNsqx91GW38AsaAhS8bnRcgIKgFQafv1wUf47yxsYZeIWcsmVaTQ3O71
SJyt/WRAcMqHZIfEZX+neRG9uW6PgwkzgSJY62bCExn7UgbqGytQDYoYZwaZWkUXTih36tEO1R2l
h1gZm82NSPw6xi2yrVPzQaaNPIk3L3xnjk+jyL0jDFzPKj941AVxbPIj+ddfAee69wLLLklckYpB
8A5Fs2jDFFMhUzQo3Gi+QquVzAnyncInKSMwk1+QCLIPMn2gbRgYiQq93K0qaRZTIwlM2JXReb+R
0GMVxVoOi+meZrd4QwbpTupe1Qwevb/RcRyn7+ELcKNTlXVbK4prPbEMxf9iQUMD4VtzlEAGQNCa
8fCT8GUOW1hlWH/Zl3nqZFFYWEGC+SE54PnYCZB7XRmrDfTCkVHkNc51foG2i7VyAk3Y/8PqtBJ3
nmoKlkH3y7AKANL86tRuYHeN4FUbecrZdNIgxSQdmqcpZpny5CcvmXHkVz7cwnV8xc67IG1az2XX
ogLysc43+e9m0Jfb1KmacvXldLw3ym1JmhAM80ch8wTO74jVCV1hoF7jMbbCYy18Mb2TzvVmqtkT
A08sBp+igdkYGWN54mJ/1R8ZQ97vZnpnyr2bUWIJF3GAG8YqPKzI/rgaUJptqVgkgSa0P8tlHGgZ
zcfHxyS0kOnnox44brkrzPhznODZ+psn1MAU52rPIr704FluSwrdjR5B6U3DLeya2JK8J6dmKEOl
LiyooHoSdVnuTdwcR2m388yATPdOK7DqYqvz33nMZwydaa4SNdlQxFd8PC0KFDRYnu0rtON0/xeL
j9a7txOGxvt+cUsgFDfqtdEPinhiYxFhlmPpRiKsQUju/CKUjGWkANIrKbTgAxi6o+0WMZEdQZHM
4qMxQ2ygq62q26XarWQmf1mmXNtNx291SNOLG5+D0jVTJibfVmQ48dL0dTO9SHRkfhdSF8uOoEND
QX34KbkG4QK3bEIEhzDO0DeVLJnaOoXoiu+9Wf6ArcLSds5HiT2vngaKM4fFiQTy5q+5s36RbFkn
T69FijHI63KFKVX81+4d4LdyW+bFFR/sxAJPrsx4cykllY34GrBh6JIjCrKHFt2BtQzth2+QM32I
T1Iy/ulMo2E9qc5a0I7WoerQSKMUWqH3GcE47DnX6j/5jJRQ6zPKl31GRj5zLyNFYgcIVxBvqcyM
FmSX0TzqiBrgIkPZO6k6FyzdCkvXWn2SRQHbiK+73KDVfahsewYNh5HA+8+BwMEUdmRzKO7YljZX
T3HbLYcRmth3tBjkawuEqG6vPtGEUkWqN3FyapvKp/uOaduD8t3bjOMOC7pb0z21NCgz5iul9nph
xLgililO338FzCZv25d2IVFLKLsKQhHsEQZqTbmDae7Y+RR3/pClpULmzqBNcE88PC21r7PNQWGT
889scExNzba57lWkWWKBNp482upHtRWfwaYtb2qae+TwcrHE0gi9dqMltT3+7sPHZgm1hbLcgtV2
7MKr4MRPpBuvKKRy/LWD4glH52pv2eJl+REycI7ONYWwzLJbVZklcHqiTtE+/Hnl8DIqroYanHZP
EMIshSVQ9a62iVr8S5mGx+LqiQjAqF5Ovkuq5yZd/bKbSafTxnIkmqpNbQJLItlOo3B3B9WPfz9n
3fWbGiAsd3ckGfjM7YklTS+ypLInf4YufuY8NjPaxA1MKRySPqXMsZK5ZCYRLdQ7Dqh1X/wbYrlq
ynvnsLvVEqc4Hm59oAdQ8Jo5v7ubVWVDaGQ8jJg9wvbV5f+zzAoTcp5ToWGw/29MAhCUPpxQXf8u
U9lODhSHmx+ZBCmI1w3pFWDTtJ08JhGtrjL4kRngEh5zM6Op5PntHtuULp3urOdxx7QcesLXbC6Y
D2SuGU76qc4miwsyn/bwfDvvNpx2WlrZ3ZdPEmpN7KzG93WLnpkMjWMax6UH7FfR/GAizoQREsGX
tIIWDmLPfEdUa4z0UcAamFSeTNp0z6l9Rkk32GAa5YoirHuv22crIBN7dSFEcHuN+o9SZkmQmtiZ
j1BP5njeT32lAn+9lunDk2XuDgvl1jjtQdzW79Q/0CivCxYLP/zP1WBOPZ+1/PEz23QRDi1gYVT7
hs7X1xHIdiGBdja9XEX0dieVIC507d3/7GJgoCREW2ClsI6UpXq3rK3z5hWv0hGnynlpW1uAX9Tg
fFdzC7scxERnOzOjKvtTJo/AwaXbTED6ytBpxkF7KM/gmrrIpxUmN9TCCPcEBEnP6B2kyJbdt/LX
CDNtXjyeTqPCszIXywasxBwuUmEJpqcUSOb67i0Aif5E3iYHxypDYOJ89217R3yCjaNUDxEQQZuR
AAXMWZ/r60QY+RF2caR4veZdD5nzibO3//3lMSAeKFYy0EMkpEPgG+DLjJ1FV75SAPMwMcXfyYLu
r0mE40+1Autu443WjaWw4Isy+sDHnUstW4abqy9QL+7yBEyxYSk6OI2YVfpGrqZsRjdBugqYZmqT
kwQ6pwinEirKSAcm2NZATu3++KoucS8LSghNWjhfUw3MYJVBTDfColkZK2AnzNlr/XHb5cPCuh7K
dAMOA4682aKt7lAMX/Hr0zWNriF8Z7FOlwqR6cArbZJaDOykG/aQeXKKGDcoqrpWoq3whY/+GOLa
TjratW+5604OSADsi3gg2OeIZS6ia86VnAKep4GXK70ZjRhmc6MMi4DAA6NrLXrw+Zk5sT2avS0y
grirfUC3matnTfQg4JM+KINI0LZ90cvB3AHjkL2qxNCYoRWR8vh3tVrGoj3YjxeEqZ418z8eGY1y
5mgLgqxAHOuKbBu9MpijmLha8ItmJIt7jFEpDKxMLVNG9dI6R8heS8rGU1z8F+qv9git0l6KFW3k
DIrumJjl8kY4Nan7P2b0SKP3W8ZPFON4CcLWImM/4VkCl2UEILP3lugp/8nYQAoMJX6LyfTUxZQ1
iO04NZSShSqwGvsmDFNWmXJJ4zdafv/pAPuxZZHxH/qIBX2CMcz8fukcC/ajAizAvSawctzXDScu
hMvUq5IAE9LMU1AdNkgcPGp0ITtDeP2a6pEzmgy1u1tmizyioINRnLDPpCeyV1rjkwBw0iuLaFWp
vhm0oHw70c8PRJORK8psOTJE5jzV+rgXyu3typf4t4WxVvfKrbejfdiUjeLN1EYoGYl18dvy54Nk
P7QIH/J493+cecG8aD3qzToVncpkTrS4VBUFbubIotOdZ7m+WhbrbzRAQGhn5c3K3yG0sy9vGqgs
uabAp5J+21fWFq6ciP2FQlycuV9GKXiDGKgOhNw5GhmWoRhuGVFEHzqucbwLCZwaffid/m85O7uR
vi+BZo+7fmfI7XNtAvxWLiwj8q+EKrOXiflUgWHnnEQm/2jrMPnbWJQQLeRemsGx2IrfrmjkGOAy
djKnMLhARL50cTYmnk5f9zb+wW+SX0P+Vbi2utLCsNg7RAMT/N+tOiJJOgWcq77o6yHT3wc24e+z
d3DiWtATBVduPMkrozLhDxOts2Ys6I9tPbOy5wbj767dDoIAgPljRhgXjvKZQJzlfHetYoGe8gJI
1qKyDB3UHnv4spJDVuFmrDpHFOZZhSIl2fcHOzLW8LEiYN2RBTllbbrncC3FeAdlQplH2Guhu9pA
lOwIH45/03Rz/9zrFz0SdnM7gPZntlBx+FXQFSlSp/h/unKDrr69sjJL371TX0fC8lkrpS+krnOX
RoB2sNd14ImW/fY+vlSCr/w3EcTuoChL65EG42LC/gkWmCmEDYxRzRsizvegGUcDS1Cvy3vifHoa
/coNpQQ47C7SAW3LvoeuPqhyI3CCNNj+WObg7MvVeDuu0AuFalITQZasCzP02h+eJLOE7a8Fhugz
HUj/BjiXptSSUEh6sraDLvRQdgZXSHH7o+ic6ZN+V5VN1TH+haKJn5VT6Rwe5nGKLchiy953PCEx
jg7dJc/O4tdlkPWaBXP/tk4VbR/3blCCgh7/RFs0VhjqWX0Gz+1UVyIJhl5KPui4B/+0tvfuGRbH
bp/4JaYolmHUyvwROyET1lv2fYlA3j2nHyjTXxjWsgLPBnUQGmxYqzPk3IZWNYyLYgbVcg2+4qX3
9GJ0W2vCBFPXKhQiI0mUInXMKzYoIW8XwvuUl3DgKYhKLABHMaz/bOpbf0LswCWum37b4Z6pOm1I
OMdxNbqCQVX3uYeqyULAPH4pjUYFOunvOv24svlAAcLmhi6feyCAO3fRxw+O2M7eYySI3cA4Mqfs
zzyqi2kyqZJk6ZimeVgpeRsg7pX+inkmMRRFKAhhmXetfYZReYl4szO32UGwxoa5IEcHP8Qr/iX0
vvniie5p3TTiR04H1oFhGOPkZXECcaQuFc6/waol6/bgxxaXazRsXiRpaDYiKQaLl6GPLIw1u9JO
UY4xdXtWit/EMshrYXuIEZwqi64TkU/Zn8JMbm7sEu+IZL/IVlC/SQ7eyMSgz+vSlohl29W79qwJ
JTKqdOO5vDECCCmWxPUTZPNXiQ3rShojQRjb51JhSvZHA6QPwYA18p7O/OQpxpPqFoOGe3MCUbFI
b6cWihFLWIK0optb5w1ccvknYqPDmnNopALFApP2D+uC6yg2Vp+b3B09VhIkODf5Bd3WDzNGQZw6
Js65An1oFjC+bBM0kxFPGkrt2wnWsOoSeoIpPY16bwTMyWUHxJPHzmT+48TKpXvh1Dk5piOVziyJ
WySsvrj+Aa5oujyeWccWsoabE4+K7qwfVLeVLWOUJZ69fHbGKZ9MY9NrJubH0s2rxQyp2qCd6+bd
8pHcXScFEUJiVt4XL9/iQu7i889k9lm7e32ich+LNUutmZXk+vsVzYOQy07Z2WCpVHaa2HCnnky3
I2V2rSsUyRZuQZMcGmd9f6Pt4q/Y7ZHV23bkKY9rNrmwRGqhuqHybu+6/anNAVHPE6U69G4lErHM
mitCEFK26xLQ77ZS3NEDlV+yZeb4uBN+4C7IH8CcJ41gAmmhR4Bph8yBxLu1PKTEF6a/GDEHocSi
KDryP1c6L5/RVNyEEK3dvTga3QVZm8UzBEgyR6LPpbuhIYnVQIXqkWcH6nEESuLzdyWG60v0IzVR
RdZJ4VNHaErRWlxPmPmSY98qg/T+Bh1anwB6L1rrADtc06UJMsn8SFOfBM+0HTrUHXi6B1ZuN6vq
wjkP5lqfRYoSoJo2OO7UAwx7RHSSyh+ComxzGUCoRzEOQ3Fa3u5FVJhWvtOUsLldWm/m5ASwMWnL
YwYLEvb54FhuMOlYz6TZa2AsYYsZFTCGhW8dmlyPBcvrn0OL93OU3SqDnXuhTC6t8ihZ/GHMP2pu
hz1pCiHdEpp4IDfUAjnMU2K5Pjye66Yv39DUvlf3vCAvC5gUzzQK7ICkxazI5LdJD664x/0NqZtX
wow5ofugkIYzkjimfQ1iuXmxGmxhsWwwWnlmUJwANhLgpVbQNHuDR0ccWHhKlA4/HHJWeozxrRz/
fKT51pl/sKdVzJUO4GUbNCKIHpTdVipFK4m+OMGvdFsSjqi1UHjLnvo0ijmyXEZDh2XMTpeD8pR/
w9YV3yIYS2dyoWFfg8+SzgGz+FwfS50VdK4oO156mh5NdNddJcP6ESZBz0Csaf6pMpCIiMuDNy5V
vJF5pVFwy3TEDAKnLw8aijMqWCOFuBXEfup32o8HUZxY+5RPQojRVfG7zdGwOunBsgtLF1/GYiF8
0cTvHq9G4INso+06HELRLT+7fsTPd123jm0HXWl9zcRB4s7ycZwhep2thEDpwC9SgMzf2mX+/Ecr
yM6VykhLQZi+Sn8wdQ7xgZtGUTkaJyti3Yr2gZdfzo0nbmQYoZUsuEisFuD+Y87y4syWI9GJZVP2
iM7UwSQxMlmgin4QgW/h9D8DiL0XXbGozcxreglIrDqpGtguPIZppxQ25R7q0fqjToZiP2GUbD2g
mmeqt5K1Mab+kFUTJTzWk4EdGuUVBehUpd1FytJNMHPDUoeqDN9XA1mqdQzs692lI+a2MtiHlPwG
H5yxnS0O/bs28EHcIOWtliapcS64S6knPLsSsE/DhVvINuXWNMTlef26M5Q4MLP5ZxHskp2fFV6s
0N3wSjq9+YNE0NkXFERHwYKQ7C/0Xj8ztjwr3tzOU27y5VTTfI02j+DLN6X8m7OZmy5VYNcVR0zR
a32j+3Dsug6Tk0LabSaokEg6T2hDLz8TOaKJEn+GuNw0l2W5KN0e0UFDsbAf3NWx57VFYzUYR0GY
iEGYe1eIGHEYAJ4q/0Qq/092lLv/mWf9VeFkjWOZ+jmctGRFxjlQKNjUmL68fgxRsyXDh67OO/rl
0A+2BRLv+C9H3HALkx5R7CFyGD1YfhPKfBnzvDNvvR0XxX+cqDRaX8S3TdS3pQmSclTEw8X1O6/Z
tAZoBsLjoE994SRiR7pHWj0sLu4F+kSLFrUrgoit/7ibWA9jJPNwS9OgM4l57vrYeWPutRVPK31g
LwIBXzn6e+06f8W5gdkPvufZl0fIxv1jtkJen9T6w70vfL6UtcbcjuR+z4hHZIlPOyFCYUgcxONl
fei14+xDpRMy01dKfkNLuk+2ii6fej88Ya+igt7T5d7sgDoT0AiGpbHFBX16Uu4TIQh8Cxo+GfWe
kU0Qx5k0/mdkXGKRh0RoS0+UVCfx9Jh5CaRoecy7V/tO0QTXObKcCF/McamtunX0FTBiTd5zzPez
/sNg/teeJBcemTPRWZSV2XyHoZs9rwxEm6RXsMLwnTIiOYDLiQLl785wguT3kpsw0AAOW/Cu5zls
+rQ1hLWRfQOibd1+zRt2Q33gcmQ8v9+kQXHA3XDaoIAghRbD1NsrRUG3BESM/CsE6N7j/vTry7vs
EUfj7zY9bbFr7g7vJM9vC32GQyKleRcucTYV2wPxpbIlEkcBbdfKlqHEyTdG9gLZFiwxkmnFYZoN
Il8F2+hDVi4vFrebIlcY04FiqDha58Gm59LqRjFNN+o3yBg29SSYAY9OwEOaip94sTiMdih/ABZ5
EKzsVuufvah1xCTwhAbejvfSLuetDvPGX+9UEYfnDhQnF10P3QQYLHby3peNUOnUxiIBIeYiWtQm
ULvXtIkk6uhyciiklh3M/8k0l3czDPX6SjLWMTTqSF/DpVxhRXpvB2a73wUoOucWIsFTq8alapRM
ByAVZdTZMP5DVBs0KPbQ6rPwaTMEi4eXoGL2nZcuWPn9RrYkjX0mHnRSEJ4k5qt6d6KAJwJ+agFB
GxwM5dtp3yk2HYhngpC0bsjgVe3rz2O4i8LCBZZ5TNSYPkt3KBXjNLDKPf2mJ9m/gPxcgrV2paWM
SYbVG9/VWV57dEYaLTKp8rfBr8wDvc1QSQwqwOCYsBj5HzZYZSAH6uyl2SvDOkxxAaKtJBm/xPj0
837JXH+ggHnqqA5eP1i9E0StEqzvfWkTReI9yn5b9V/qrjVxqB+Knx0v5KYn21S5oySKxWe6EjKk
I5Mb+bkdkBNFQ7ZZFGsmA8rzMtITh6E4CFxnnHbjk4F4Zi+9rwcqqB9eSE+CRWAP+Wqqvg6uIKiH
mOTFaD4siLKdGLYOkvE8+rD6kafuW0KVNPS9GxcKS+1Fba45cXwC2q6QdKfQevtmcDjxVlIsujvH
W1bXDgopU66geItU7xVs0MN3e8hmsKINNVJX+7Ix7jOsl4X1OzNpgc3/eTDlTugm/pTd3gcamyef
XoNdM1nlwLdGAr4nTf2IFhkpcB4oZXI+Szjzy4lT0I0NRAEalQT7sR/hbqFoeY2cgnSac0/Cpqt6
PxmjSxVSD2wMpk/1odBgWmgsp+nG1fhiUpA/qg57519eEdLAtRttRXXojxvXhRNjzTbKA5T3BQUp
XZ/M/vdEeFSAUNFAHnHsMyAOxixO3GMys4yfAbfCg/RkaJjQu/Vcmi/QyzDd/tYR1s8sCzvj2rwS
CDyBvll8j83uPEIjQDJSNFQaMLeWuBgWrNsk/7ZjzdHEYisqiWLA7v74KzCc4WKLCw2/KKRWuIcF
5/ShQaZoEythJ3UgHqTMORdy/ctvMZ1Ekuv/1fmLPMU4hOXOr8tMRARNFtKvTQro/Dyrxuy484Vs
sV9Goq0N70jDxdArxwR7LQNZl75oAcLL212EGeXUoY2Vb6fEta+FZzNWQY1vS+2CRIptAOdZud/D
kDQzg4u3B8a9ZX1ZHL5VMQWMG+ygYEHv7RVGqsNF7qfEVEejNIOlkXZBKSxcKBmkX+jOgJgrYl/K
vNuKWQLRfIDE9HcZCRyhGWTalmaAuBsTdRx46WnamUDPbLh/Pq7220O2uX8hnnInpl+7dIaoGqPJ
D45PAt52w6wWJb7DzbpTSlMwv23o88b3VTeZBcMLPZDM/Zjyw4FZvBYIiIGETyHV/X4XqtNxGV71
WnkyVHVJ/4ekb6If0JLAU4zYrBV0Ahwwl/H5GmIjq040E2dZRWdoE887hPihYFCo6vaz38MddDUo
gPJM3QIf8eohjbM+Q4muMgokhd4lE5mjMlAwzGa/vqMq6r6ho8frx3ZSNs6iZDGzICRi5NdoaAux
P9hYpKe0WBzQMAnX4Hb876Y2kDL/TaWCd3pCMEd3rFFYYtuSbmg5ZvErnMhIB9fTK4YzyezD5fOG
rTtVnZSoS/IBZvL3/NYW+7qMaFtN7DT3/Jc+2wUE5WqiA9N8fwyr2PJsY+XWwZ39vaqo02I0XEDu
uUiuDqBhN6/w9W57COeyMRfKTffSCZyGG5YuZ88p90Agoe4D8MNEfOf1Z9r9RRG6590IGE4bU2FM
a7XLwC+Oplv2W7U5HwyCxNeyFF+hGHA/SejgDOZXJsxWSCN/JEq8zwDpLdpobxU6psWrgLu4xaL2
ep5UCwy6XkL07GK7B5JXdIahh4bv4LaQTNkEDzBx999ZgPmiCecenCq4jISh9wCKroubd2eNEsWt
qY5Ind7/1p7Ntmf+tDvLF4OMp/MVVr2CT40hXEAregpVXsW6whrA64i45H7H7plhbQJZQtjuZjla
dWZTPypXwGG2uBqWyAXL4viXHGdedLTx0eSZIWsoaCRXu/4IonA9A6Lz/cqTFf8MS9NJ89lv5Mj0
+gUwDeS/YyEA5ZKkJUssZSK3CGhTszMX5BsROlKx4ofyAzvFrB0FvKEQCgM+Mcx0vdfWJvnP2Hil
q/MvtjdLwDEO/tQCF8vGuoDbBuOFm0cucFNrLqEanDob7bmte5YCmG0IE9ydNwxTf2MlBxDCyqpa
eI00GhvnIp4fr5mhwLWWpThaPV+jKBUQSukMzJjafTAXLxIeb3kcBLJGB6XkBT133kYf9rux15pw
F8hHknpWGsyfeKpHKLoTH1248O4uRYYczAR0dxK3McZLqk5L2G5xsl6v3n1ymIvLhGA/C+n4jWOl
Bb3QDqyFZNWcMG/uvMr8TS8x2fgMAotR5+W++aKMWoGk3kaPDHrrb37DsKKKSefUKw2nMc7IyGav
4IpEGp1bHulWLN2/jZLVs4mz+zDrWC/L2+dBuulc4kg0eBrIMLRYUq8uaxhUUBfidnN695YLvHx1
FRfnIx9v2K53vHmNKj+zhqhqVy/9f+2yEZbW4TdDwSUoZHjwzNvM/+Sfe/U4gymdK6RUQswBsGVU
bKS9pumkjMXpmcze+VwnwGDv2uzHd3ubuh2CtpCuy/gDFfkWVbs3oQFmrocYYc7bbchKQB33HYzw
AcSZ7UngSQWi+h01Y39UNqTZtOOgLHF0JM3q5T0pznUL3pEiHKwpkingG5KoIWc1BVXieuoQNp7c
7Pisnw9qymrEclL9CCujKvQ9DfReH8uqRli1nuy7o+WjsTsRk7UUR5plnY2KnZZHL0WfWl8Fvw7x
jK+FJ9BOx3prioQ9YnMMh9Eqi4LerdXMkv/MjxOBD8+D/7RKH3r2cL7qe8vZzm7HDpEKVe2o7QHk
X4y+BlRWZ+0+5AP6jFzic2WHfqLiZJXRq9ut9+oyHTKeb6TRNedfifztng1EUF/wLducyMhJP5qP
I8FOvgJXq1qDvmGpsup+K5NR+1DsjcqYpIhW/hk+CXxbrN1vM5OKpc2xd1cHXH9T6+9UuQzUMluW
Xl4Y10xq5jCCgxHNXJp3E6/zWc8Cnr0YfHX4Ra1Nx0E4B6zmbWFe3CRQsGIVOTAI/kuaEI/yYXzI
IH4sfNjPg648E49HxjwVz+OfwjrmAHzdO0iruiVq9lnhb4ymNtC0e9az1NkfQ+xJoPtKYZ0Bwo2c
dZkoqm5nxI+N7mrlKG0JpaPopO8XPAcFqW5wH9NQTGXo5AXOumDHVD2YZ0WdbbPlnHUSdLzqAwlk
yh9g741nhE+cPZ+bgfy08/JTv35ci7KxMhX9C1PagCxBr7aZ1WMGyMn/oUxQVx/Uld+zU98e3Lbc
fJ/QPkQnbGPvfrKx7SvR4t7CID9rn95dKlCFUmbGcBgMGSeZbmXsMKuQ4JHUMk4lWXwGndfJpXeS
lXOderr6KlZ5TCxNa8DVmuGpZvz4aFhKt7I1BvKn6yIeerZsTMh8HDOXgGIZ/gIsLM4NGDL8gwAZ
zB2B7ekVEqXg2dviZoeZI0v8IWHMNvEpB+VDcLOZ+rKW/0qc41zYKuhG0nzXH/g7s6sAkVFwKj2j
aApyqd1j8WAjVlg2fBb9rtG8q/FxAKCfIJ78SBQcoRgeujAUd+8lekfdMaRGs5nb44rPIrYzoL/V
HyC0wfG2pEt66CtARlbQGASq23yUN8ue1n4ZkALUaCbTAt5/Eg4A7loPGMOTkU9YwkNOuCb2tih7
8V62Cm4191UroqI8j9aCOmw7VWTMcXfDywmrYCgf/zUw4lFexJ7NH4CtIazfBw3CgXV6dcRykABs
ui3mUo7N9Je3jo65U3sLFcOHYavf18Uwix9yUyWiCRE3f3ESRVW18qYghgKK5GaO2+MxnHju/aza
4P2sFrvH2l7M1LpLqQPjdtCyFcVL703TvHv838fAw+xjAS0MjOoXnqjoCVDhkvDt2/xf38LCDwBc
fe+GRMOvaQG+GFVtwcLq9+Hv/Q/Kgq+vnQwsFPelzzn9XECROIZ3P3fxcMgF/ALv++cDTj4yBlHI
N0r2Hjuou4py8dj2c08PkwgPC6Gz3cnBiUI9gJPybRqygfLjfJvEZqLAD0AZTo+bQPuoz3Ra+lWw
q3EykeS6uhp5dW7dKFZX/2uh9GnrkRLg1alwwqh2It+dAY1MRzF35L0GXnjbCCl9zRsnS6yPlHcR
ED8p1I2TSSCpLERh8aEBzSvCQRKBj8aZkO/aPKWwaBR/B0bEoAgnah6I2elHencNj8VyIhjM10R7
g0sgaRRPBQn1uYDwhpog6rUrrkPt9exFAcMBtbNcfpSZvlM2VaYRgwcAn/VdRb9JhQZhX7TDhZyG
hgjKuyOwwOYOjru0VrFpBLodwrmM5tVAgYTPC1bH/etvAKDKiJGpzn9Z5ED32xQXL34/5qTqhsPN
Dlm5g/qZmofcDyLK9vXXmkOePPI+AcHGD/AiJ2oBuC1yuMUN2h5CVZcrc2RjhNjLwoHd03RWLad6
rkGyLzkp/YNrCZFGxB57t5wCL/Bk1bdNXH4Y+985vFDMtRoNC+ZG85uBSKrjsboLQryxRGl73L0K
SHATtA45KLcQBGTwbDgBGVICaZkEeAt5n8K2KIHR1j7waThtZaFd+ilSirJ50gMG8Hvc4I3SiHDf
Epp6ERIMucECVvTOvxqs+4QGJOJlQaP1bw4yjYI4+Jz2mF16+VnDjhJaKgWpZelCcgdmU4qkexJD
V89Y7upZTaMuVlkOfPjpM5l+ZPdQGR9Ff9rMBCiP+bhUqpvs38ZcwBWhsBHW4e0IFBPToJO8P1tK
YTl6LhB/vg2NkPKtjp79r6EjTwfJOuqhrwMmjTBgUDS0si9ZHilW9aQni3yk2wt3SwCfuutXzQCp
ghfjXt9Kw26rYiGYuiWLv2Q2LXokAivJLkorgGT93vcvI84oCZAkIw6GKpv2/dztmg2TQlPzcjaO
rNANaM9Dx97WUdtmYt7nkJ6AttjpGr5LgUA7Kp8LS4SJ/aOUB4WpUcv/aMMjoZU6ulHTsl4HRygG
cB/wQYZejQ8nX+KR1rwms4vMjyXHttWbegP55Sh0F+x0C/4pkBqbCzz5zKDpOqvHoI1yuEvrMpX0
NiIY821Sm0GJtbpvAvUZQ/s2MSx8Iis9TOCA+qOEWhB2/P5VnXKEbStomiEqIHRX4ISa7jLrAOKJ
hqT0OsE1j/uweLcpvNbWqFdCVyxje8uX0Q13cn0BSETwnyFKvuzNoVfnFAroX+hoeDjsQah3aDAc
XdVAdTsE3nyzRFCoPD4ci2EanWFFH7t9ZmuL5BgeztjKzpWfvEEmvMB6dDhPZaaQJKmxclkCM1Gh
KS2uLXW6BRfKwwIeMcRi3wX8Km41bpe0fAwfKMvy1PCqQAT2tiYITE0KoyzPgTb7BE3FC22lXuy/
CGGvcaDmbE/g599e++PuxasRlNb2EkXtRDq7hPlToPhwynhqzGnlSLyGt4KmI3zOJehGyNQnWSZo
ODBxqENBqfhRN0oHW0iIExEGBEV4XVXJV1ifI3boRkyXGOCp0xP99IyF4vmWEATikuw7fGk8cDVn
vD4OYHvNmSwGOYyQq8oveklYYkaLxqGTTVpR+lvpZpdnYLOIDZ5GXYGu3mbj18FxCMAKDzecEvy2
0J6h9yV54Qbp0HVXuf8ZhLWJaV7JqQrdDLW18aslIlKCg6Ye5jucGJVAKf2sI1hASnuXjz8sZrDE
jROJLr5hskwk2R0mkM/tcFVylHUBnB9XPsqWiarxE1jq8Ui/mL/hKHuMN+3XV+/tikAXwsjiMmWD
3QAgzqp67OiFYHdI1s2N5S8WZi5si3NDQcHTF3dWAACG4w0AAG+RZ0mE5RXgfv/tw25VAKCkydrz
/3YYLb3iZ2j9eS+ix88ZE+nCjviryZ/aihndO6Sxlnh8xSFBvCEnDzcGIbcrJkGG+wyObQx2vAeT
Ua7um6h1qMj+k0AHJ0cQq0MjO5TRr5NQ+irAhn9vjYZkavpdQlYXL8kDZqK4m/jnzcsEAI/kO0LC
Io7uy5Sl0t3Z0Bv+ruaaadXg9c0zw0S7e7uUVU3NF+8bQpdrTcsr3X0qcLSa0bMwWTwlhQo6lpYu
6s075i2XybXmpdTf2hXaKQeXONUovKSuReuILyXtOqJ7Qau59YWdeIVN22e+9n7uCO8A81R3Jdlp
DJbNtIR1XVKKuo/jwDXRiNijJMv1YLunVjrTvvlA3LG7D50zM8KQqezGBbkSbTW7Aun9qJFWn/UB
n/oeW7XROIC42iKDVKcjZMZ30UyuwV8/Xv846KH5JVxVjSokBRdGR6NXkLE+bdqxWQKJaHS9ARrN
aTd29y8/OmASQXtUPHyqGy0DYU6LssH0CsTE4pg++9bGNofgz+1KtQB6q/gqEiQECfTMO0eNR4er
j+5RpOiAU3EIW9Xtl/H64/KuCZGBk6kEljlTL794E9FlBn2tTGAh+66t6+k/vE/1CsifHyfw+i9V
wEXPotEov5EnIOXiIUMjngVdoZk9n9UB+18mmqBiVB8s10zgR89KeHI4Erjq8qRnqrFHx0TMA+fN
hwR3KvqNtFcWVTqB+GK1PmGelrkVzPj738EU2bwbWuJKDcVu0IcNE6VWCU67+GOcJJKafrcik+re
K6uXn3yiDrRjma4qGEHzIXEUdgC3bVc/i1rIbbGZz/gt5UIXFTlaSBHtW0dD0I/DO/LcOgHHZD/4
VN5A5tpersdfVB9Y9VzSuZn31O9Rouvzy2wVWx75EhoMYAx2N3Mv1G44Wyvb/SLbalcwfOaWsXQe
n59UPz9U1jI9QW8ojA7IkUh0uY98of8qHoSgKHJkXWbMpxgBB9CAtbR8p5n77H9iZFGHgO8Mpn1n
YO19xryuNkU7UV1s+BgualL7kE4ylb+gJNuD3V10JnQ2IhWwyOoECBS7OsNAl4HhZy5hc82mHdte
mA4qgWDzzdqedn1gJlR9Jde4OVre0R2NxpcNWINZNxcpYJYDHkze1r+PSfcKNGE0SdSdiAIDTAy+
Pfxqxtlogpv4mZHbryMxgqvujaKhT2W1MzymEFouaRXOktkKcba+73zKf7AKrJTJrEIHxNAQpDUh
S0mOMVEYCMMYFkjNImsWWmnhzMroy+MBWODs1Gy//3iAI7KRXKmhEP6dqAQ5sy3+T1Zfb3TsTPxC
zFhb5/KyGyCdBQPTTgK8bSFZqvqg9hRxOoo10fvle/vW5vhBflK9px8a8viOwslC5L7kzcXEQ7n2
U5MIfMRRn8WbzQYgXNozCOXuFxoNCG3SM9tC/7GJwGk6hbq2nyahkGBd4DEF7EHfgqHgu9yL9jPx
FL5WaUJNRuPOYO/hDGDfEOw2JE0H4iewiYvx3DsfZjBsDuxLmkbH8RDY96RQ7UZfMePUNaxh8Bq3
QqbCRx5FjYkEPvEGTPqizXeMwjYwXuytph+pA4uYNiclyskc4XWeDuRYL5Fk1VbKCEXxDNf5IoQq
mFRBj79TMumQZw0HEOpIm5T1oWAxxoityue/F/PGl/Jt4xi3gRjOQYeSSoBLKOdrI89z6TIDMgs3
gAUPBgw2VlBZxh+yBk5boS9QXLGtPZbmu8zNStahGVmZaQuPH9mQ685Akkbul3Gqxcq0PwyARvGW
WtCG/Tt6w4BLyLZuRIPG7OFq1pAjSBXZudFCVPjObbveAaIdZ1YcxmLea1utAvPeNWXtsTz2Raou
NJTz31POU1HTxRPGnIH5EY3+ix46Io8HOLo3L1fZ7SGNCRYeAQE737ttVNEF2YUfNNxSGjbyIioB
omDbIJKUDyDCtIOnuOhBGu2qisq5iFPkcA5fTfpmXbMBD6ehlIMhKLy5dqdxxuJL5jwAJfLRXwEh
F9H7+e7ygtqECS3Mvkg+/jWlZ9kn4m8N0kJ70Gkt82j4i+RdGh/z4pMgwU6tpZyTRSZdi0QMZile
85l37kis8hxZr2Vqy3lJGV7sMaWVoC5krHAsjufo11s+HDjAh3zszM4Rqi7r2v6Sd1D7GMerxQ4A
UfwOh7sz/dPOMvEtziWeCF0bhkO8YGak0zKGgzkOPPJXVyKssW0krDgDDrRnxpnnlbhPfqRDboZO
wsubpNTv3y5kzwgjB3OBZLpPbegbZImMx7vXFARYYonGHQ5/ctPa3a/peTxgevjkjNos9KxJokC1
nrGJXDRiDanx+ttVosWVhIzS0mOJSzokxRy4DOrywUdLslDsmx9n0mPX/eV3kj6szon9+NckF9Fv
ZntUF+M9u+bTxnvdgDWtoDzJUIdjegJFnWlToTLXpiRyNLB/g4dVb/D+Khx3WnOnS/Cjwt3dA1XL
p852uiGwSbpBlXKAlplZnp1Nigce806vX0VohoWUDqkX5oHk4FAr9B/wEUusR0gBMUaoWn2y+2+P
c5Zm1E1LWMrDLQ39bq4xkbdtAhGhiVKUnePcX3u4HnPhejWcBzYUCK7uEZf/CADX+3B/PWJUJxna
BQqYVJlpSNY0Fkf/YCWm6pNuFi0Y4n017MKb1RTQg3XEXU8bMCe2rIiNsdUGTBEepIHbK+IFpWpp
ev3iEs9pTZTJYjJ+d/FxogV+o9/ephUgjSrrg9Lc1zdn3u/6nFawQCmoKCFQuNsqmIlr6o6Ug8kJ
qYaDS3FbkCB3JxGurethCG9Y7P4b/phu+fiSxUalz6tX3Jpzzk/kC3ZQuTxZo77/O61KtOseSb/h
dc4oX6If1gZAWc+zMq81WuPsshe/XpPUSjQLk4u0hhHUXg8jRyO+o7f/+H6yCALuks//aDA8NtKk
4XfzhJAx3VhJ3tl9Ega3SRiQxTRrF4aXjc4t4gDTErhMMtHlcgUaJPmUP4Tzjm7m0xzj7MkoBGH7
+EVSSBC8sxviIC9cI1n8WnZfnW6hNq/0G7MfJqlLuZcwuAgJ8lQ31shxDwq3MUx2bzsDYL3zcQTB
QhLDQBfLGOio+E0PFXsegyPyIHRKe5UyYYkVLSdymz1wtP1LPrBnmd19YEFOhmohzckFM2fQU74U
NrD2x+zQb31u8Is6rNLzWAzE+/HsE4w9uSFXw6Z/KEqVLAniYugKJXZo9LoxEaax8vpqmWNAz6ZE
5rxg50sDP1UWknqHxMt1kI9jnN+KksiteL5QjVKSY9GrBJwn/b2g5VF+PBqBYfJzL+rQPlTaSx6o
39xJjs3wGtm+pFSKPFjfwxn4h3/qJSp/Pf7QlPR4oBtJu3bSAXhhWw8j84xvLJjMZp7xqlxRTJdd
Da8ZEETAqq+VUL9T5ixzPGYEhc2nJiNdKUjg5ESHP1/8O4v4VTU8SVicPah2MnYy7YjRhw32kXzJ
SIPTFCI0r0T/9ylTDD+Wq+UZ4aSFRqiAlziCuHbRTb2hZOdgai9aKkutkWpmk5YNGHqg5AXq1yXm
f5u6VjKI5+IftyC/0Tsbr8XRSdK8tzFeFOZ94jppAsod0hwH2rVJy97dLvAgAK3Q5P12TGLDUdzW
Yfd41I7JmKkOTaF3llIck/dY8fQA2xMKASMEro4pl3CUCWVq/OgrkJti9UuME1ilqP6SU90kUja9
AgQIy7gA9pJzrjqSUgP1LIa6Gfr9K7tFBZprdYNrFr5aLLcbEizvVZHblId2OUGXqNEexnwixG7y
NsqFCrY3y1IefpZebrY3rlrruDhr4IBTBvLO7jrtYI7Md6KHcnpg00DO7YqbXC8QdbeKnCZfNYSc
5LjZc6mAcytsuYCXheFO0fwKRDBst/SPrLyNEi8ijR+AZ311blIsQH9c0VGovvX/CD+9KPf+dGvv
QC9DC/i324qNgwOgmIbrgh5EKLj0xYof3sCrmPQUOosdCYssiboTNGI74hjlbla3CXSlk7KtMVh8
Hk8ZfwLcUaIJfHop6x8DUaK/U2lz1zSAzCLGO4RFbWpEGZC4aDluw4MQ1JC3i/GoFgBcWdqb/zzH
wPEWt61lKTd38tAnfKg84yr0B5BISvYSuQIUja50yI0BeRsmaCAz7P2n6nVe25E0DAPKp5iQmswv
k4WgtijBvl13Plr/xkoqA6Qx4OVyA/zuoqHmCE/7FJftwQXYlv7GMU0v2tmEi+OpVJI/QGyKRA+K
Gb/9dn5FAOD52COASzNVeJDhZs9o7TrlPwlfuaNcevBb2DN47D4pHEmYgQbNET7qpsdWOnOfOkWq
cRrTy6csF9ZFpVoui45TLx8ZvT+mpA8Bo0rqmQfW99FJyz8c+fSfOF/MW1BDM6iHC2WlIJpqMCGA
wfRq8xu1KZRPGqcH8cyP+BoE9l4CjTICdc8x5uiGmHJqDOqZ7TLmUhQb2eTJ73voWlrJkIVQ0+aP
7kE+wBOfDSFR4tu7PE35Kvu6l+XMZZjdiggzUIpnH57qU+YupNaWJjvCGLAVuzkUYWmM5l5EzF78
g8s4SDtNXog3jcPzyvAMMPzNOMGL7ilIM3NeJLkdhGCsAuOqCqlNna8ugOsaNCDmEU8ZQ9JU7HpR
oFzBm6JGWoWYVN4OzvU4wMLh8IvxZKENoYalaaruzVTtHtznpvPuRL7LJAYnckJ1Lr47nPjKsQ4f
Kxcs1AywkzfThPuyAzMysJ1XjLkB3RUdgK05St5jhf5+cACgJ5g2RH6CMJroLl1AS9vgqT0Rvcvq
K+fOWxiYJZYj8TIoB+fsfI61qNCXAnmE9qiL1EA5MU09B8eOXbzKue6roOb/o2JTF2siWwMFnGkk
4h/zyYiMFDxdGgF+T6nfo4mJQpFjQHEiFaxcrHAeuOvdIo8DIZ5pkIKlZGBOHjXnq5IkGjWKlwUl
awmWDSJZo81L+PxOvC1GDQFVOHjJXQbXNemZTmL0IYjiFGKJWg8K+Ca402I7WGYUlm8o1vomT103
ra1dAK/4vCMrrl1mEBamS7IFo9Ou99q8YiIIwh4jlyCl9DO6NA1ro7qXT1IJOX9itlMeV9rIhGa0
u75DufnCDsDVOqh2lRJt0tZ3+z50C3J69m+agNHGR70TJHNnxnZ3Ove0tQQG6qC/dTxH6ie2lNLy
+hx9veJuBv6PdnEe9Hph/m8N3cl7D1OcbIrYxvdIQg+JSdVilzH284llHqnu3MOskCIWdaCDrHje
m9Bv6KCI7WIbTwquA534yG3wFNDBgJpl4OamVufpfPYkJVJNKZ5DoP2efjuQJn8K6Py6vT6UCpcM
IQ8cOLm/uaXqO7hSHTv5Uw3/wi4xrONwUxHC39TG1L4hHsYMi9eIuTsPzMoXvE+UVvo4Bvlqsut1
pazlWy6FBpsual8zc/8/RqJrwxd3yDLN+wjR4hi0lTaVJH4D28u+XV5uNj1x0UW/ZqdOrymvp1i4
vqcp8/5/H491kcVB/mhEhACBYrVYt0cQ3HofldBpzQks8zckHEbOg7+eVlFjEuUy37EXB8eyq8DL
yiaafpk/mbFjmu8N6WunJ431zrOuSbgg8xATiEPIXVS6R63wM4XrF6txsPgHtDGIXfDR6fCDAFW8
12RseqJo0qQFygtKEgmFqG4CZnDK0fUtfbx4LPO7HMuneqQxFDxC/FFwpbYfetIceh/y8ADWaN1F
1l4DP3ob+bnZw0FxJW6XliDhwAjjUl9BGqr+kW2PjioQMqYdgQtTYfAr18Uh1ZQDNr9zxZcTSJiP
bnm1doiVqBkug+PkTBwzJ67vfaBoax1cGT3rxBPg49Q++RzGG0kKZ7iHyvYMSTeOuweKDhBuxPhi
Y0aqW0DzmW3z/mKoYlWeQziUDc4kb+IKQ+doUH39IZq/fX+vXT6d/fGqwUpCbBosoIDzCBJOe+n2
1ya+VzGYHVKKHKExzf8Rcvty0IhWxEYKQKVGi3Mx4HW9ld+jrriuU/hvah7w3oqDHgXwL7qi2FYk
3POagPcRB6zle24FAOmiHute7IKq86J+tZN7RWIIhlu6ok5DUaWv99sUb/mW+R/UyqbdYLR8LzLM
owpvqxGqVWIyJlt6x7uhmpTgJ3Us41hJe9WPrNb5fyEwJxMeiE6PVPu9mqI9vLIE6cWJ943pZWR2
ersd+7GDsImeD83+GkblINWImG3HbfJNAF43gJtbpgwXihT1LxXoUkNBE46WcwaGDyUWvFuhtf7y
9x7CP7kzLLw6MnbOrgmdkbLH2/wa/S7dQ7W2u2nRHqtVVm43oxzcWXoLlperWD73hn3G+i74iu3G
Z7RqTg9sW1mMsrbcTeL8sTZaHy3dCFYaNu9TORtWteYRFz4qUXGSw4lZdZZUnzxFXtSssZFyUIVo
BhMaK1jLOQLxLkAqyUbZT9/UU0M3bSFkc1+qwGt1MviaxBUG6gqNY8NKL55d9yoKAmNRAGYWLcgf
to0QKOhCt7iZBFxsrE4hrj/8OV1lvMBu++jgPvKUHbyypicgDoJpTle3KpvT2dpWjjdQw7kRYdAG
n+PGlpcPIZfHPMOzm+ToxLUMFpoo7ppswzJ2lPheNukGHdLADCUpBFA1VOUVhWniEgb6n9P/fgmz
GrUpDHRaqNQGCU8qrdD0bx9EhmpYVDplQbeJmg6u8Uh/nA8mjdyGz+Fc80xGtspNkITj2t4Qkoku
fQd8NiLW84HMfEE2LhxVGdlNQ/9/m7T7IfTcizS1dp/7wbjbtAZObhEgHtUJ97GMIzwmQBC+rh2G
qOfhxpA4/w31bc6frSW1pb/jflfyPiWrunC5Hg4EG0CJdbyuNYyEcIxdrZ9YKz0/cJIR1QV5CqvV
7WPo5/Idh0pGjLFaJVxR1ZE90cE02oSsmBNCPsxsSYe8+FJVfHaf72kCd5yDhoygYz34Jfjm3xt7
C72rxroii+zjxI6PdGzvaMpgsaWg6sz12gDtSsXE85xrDLkBywaxESgmNjKrX+d2u1DTVrWEfa5x
L2kMX8lYg+XZCibwdPZMexGzeTFzQPWc482cdUXD1oZnY680nCMTH4/0OvT+YpsOU7wUt7mXI23Z
wmA+oJBgzbg7vB5eX/UijpTWQqaJppTgI8WpbtBMPhIq9JxMdy6hvxwzdA7M8uWmRDYaEcnjOuMN
I+iz8HkLaWedqshlyh05pDaUmi5OVC43q+br4qo7PnpBUjvWgzKejqrTqszlKCiPU7sEhey9r4j1
eof4pIwZW0bML/n/tnmR2M/xDnw0/Is89Fj7kViyqk5UxeKQDiUy+Ee1bIBWGFAJyuYZEXux0Z7i
nAEum9v40Be3rOA5SJRtnmhaeq56J4KXi8WPeeD0WoaCgwbUfvGClsQINv+A+GSkaaFhNfpIubZz
GrW7g7Uplybmfeqhr7qvYRV0JFMZyP3CqnO0FnsgFNPxubDr2DXOtIHRo+v4i9kJDNNG55L7YNsu
WghxGOeuP/l2Upj+UsRMstE/5DsLZV854OgvgzbcOA45uj1gMsmaK9CNF2C1Z+ly+Cbb3rZOaRch
GOATZMS2TM6gIxWC1b5Znf4x8qgk6SKiYS0mJrVKIX7jdYGGrVYn58OM6hP5YUyVv5yapBy9amOn
ee6sdPx2RdNBkNEmV1FkyvK/bhWbEMjfNn/yA/USjGAo448RgnQDaU0hvgqtxybB4OWG0UvLkUYo
Phuqj6lyawIN54Yy8FEnAhhQPWZKCsvr/Z51xFjYxY9hhugx4CfKPbIZeFoYB827SERHPL/+XsQA
rJUnLsmIr+i0hPAEfeCsEzB3pDVtG3Qshete8Tied8obCMQa89xdCD/9H/thJE7lzysHXaVHkUPZ
rCcEpSACs6FZTfrh1yPgkiHpFy02lh7932Wfkhchnsui2hgvwcUsJv61KNxa/+HNycJ8+gTi6R94
Bp8wNjp7rRquyGRz0i3o30OslQteL7Ya5Zs8CxuAYRuzvy9y+yKTpCMmqMFHqsplZQHERK0hBh5q
wcb/jVNHBgQILD2DIeWgS9jVuV7nLumwLx+EITdeDYbQNZE8/fmOwIKlzuKjdKvAPVl1BfG75cdH
shmOlPApQV8HpqoE7E74jDVfDOjJkTGbSxmppkIAk/GYepd//i/3UmAzRkKOclOagK0cEYL3vBmP
a163eXXxL6NlmQfYbB7ubpk34Kk5MMY8QvHoPYf8B/IwHF7wPs2ND2LxEOOwHj7QZwSuo+0PI22J
LAXCstN1kHMr9mxOydr8Vg2kuXi9RrBVa9dM6S4MZLZeZMG52Z239hBJ5SWYgRIIiHAL0M7VkUz/
C1SogayxRKE8Z3CB+gicWeAGIIITAV0w+z+wZdin4qmqEv7wL+sBzCLEZvgpZ8qbVWm7rQM2pGUF
kp7+y3d4pQ0xCN3l3bDUoj1l2OfnsveAB8v/WPf9vW5hbCx1cCJloyJLAYTd1ABnATCDmSzAH6ws
m7so5GwO2VJxi/c4XCVn73oVY/CGgVOU+MttKsLOIrxWD7QZUzgkIAKse7nvtkNFjPEwRsVSpvyT
TcB6h7KYe3FMPDJnF1BEcr97iTVIArFMGYDW0TWbKal3umAvLYVjn9r05tVjHqRh/6CVlj/E1TMj
WHrAgCT2BN6ZVAhR0qcGJcK0A1n40w377PaR6uLZT9iUx9aGl3BXwouc0+xHZQRL4pSYRN73c3f/
xVSpGDM4rEL+zSTTW3KJ2j5I0bs+eKru6Le73gH/08ZSLIt04jBFvR9swH0O/+PWFYJS3T/AkfN2
uggeM2rqC/2C6sNjaJPemtL5zqCl9+6VXAeCH1HJh2diYLgRdaBChurrd9EHq1I6q/xizWBYuAZ8
Z2bsnp68b00hYZEKJPcqI2JgGHd0Ve/uXAoixISyrMGdVMySFH48PTLrEveJpjvo55oV6ra38W1c
wEqaqNBWVShodRfqaGt3phDIbPKPrwQ3YoqG1OJ8kwf13CJMIX3vlVNuo1/VxlNzkzxyH4bL1ZlV
EWeyMSlZEGzQwyNc6MSPqlITITr2JJNufBuYl0iX6SFhSAYCePdicNoWBfRRp82jo7+fQX/+Ya1W
IH0JdNkAOcKMX6FLGvYzsMUlxCUNou6qXkFF2PDZNwGAgotz21tWY3cGsRKR2/57jHxHfgfacJM0
0PMSMoYxEaoQxrK1oixA4NvTJJGgs1N4YVU/sCwMX8bK3JnrtFn9gbbfR5/18b7nbqfTqFWzS5iZ
Nj/rr1pQWV9W0Jfs8I8r0f0+Z3KS5ISZJc596CPjL5jkTeNPfTnyTxn6fUg1O6u8F7E8qClJZ/pB
Dzgu9sE7BJ+9V60KBLzeA1cgmcZ707YRvQ1Z6DLTu+B2Am36o6r9ZUdfyZTc0D9Fp4dLlAp8Lgcb
eRkEQmyyjcYUKYLKohZWvur9Y4VnaJtsvxtCIutLh4dtKN9GWu5nrTirkD96MmjCHUe6sBg+MsTI
FsuVRBLdLjSLZkQa7HzbZwEjlKTezaiJtbPy/zxermidil9ipkAdVbL19Eg3hiePWEEdOjLBZxpP
znx8OGkMsJpNDMZPcE0/DN47YwTvYrBRiaceK3C4fYTfPKJA8JvI8KR3CAelGUy5WjgHAvnrw6fa
wnHkZBEaWwsG3dxVujlqb7LhZlsCoYlO4hhkfZHVwsOsxYZl2t17BtFHla7az7WVwieqd4bNJ2HZ
TjpjGlxFLbz4HXhjUbsOJ5FRuh1GjTaTaSYEJsENorJOmWpOBq3h0rs3Fd8MwPR/r1amPyStG4uc
sJ9TeLPPr3bg+YcMiT2B+URM/w1Y4V6hXfkt4yW7aYgXHlmIZDw+c4uBpGqYFtRVWxETLWGwGM40
l6cDgv93qxYuurw8afbBqrwwdcAV6l4WDoNn9+yKBjs+dY6ItWZ9iTVcAL66fnz11qm2SlNn7Egl
+oF4FmNhC1/Vs4M2cqZnJJEbnKHX8aJHDiBezNXMRS0aegpKTH7zzdiSDJYHZrB6QUZCbbpTJQjC
8sjuu+1XE9OgRvJkB+PsZcGQMV5X58XfSf9sO08iDsYCZq3MAObjxEodM/QNX9z2n9OePz18Qxlv
aZYLC3Qswgnf059gZmgyXff2bFALqiZOCtW8TlPmthddBw2JP9epqJvsiiy+rxu4iN2ujgY3O/9O
DUPzQkHGfLsUuVZVPWTwaDApj3tt5DhC2p5H5OvpPiYE48u+67vEMn3e8lJM9Z4vEg/Yrfq2jxCk
MzfaYLuLKmzfXX7HjU0nD0O3pQbdkGdJzB7iqVYcTv6YinRKhCck2mlph36i/EZD+qFDfeSF6tgw
PYQrgoOLizIG5RoW2H/PUFYMruBF5ZnzEUO/652Dva+DJ3btYLy8WGhNJky0Dp7qY7544y0ZCJE+
GaEudrrnkID707ou0hb/S4E1XcocsmiVtiHJ475Cm6gT4Nb2wMT4qtNZuXcQ6MidO05sZI7zYNQJ
3D9+TLNDT6u2TvSN6pTOr3r/uTdHGKTL7tXDuN1djbf4rUawRME9scGv7WFxjxVgCfQh+FL3BzcM
Wqt8Rp2cWa1k2redPkPNB8WqE7+X3ka1b0d964vNZj18z0DiWVgjWz2DNmPcPpUWvLY/5plY1AiP
GoBZWRUMonMAxnRx9fqznE/mhxzkhzPLmsItoyLbtkmy0dYTcZH/amq8L3ek48fAxGdAJrSDHsCY
+1ZV5s7ygWekZ2+ljAC5E5JMscNPM3FAnnITNvCxLN6XiEunq3iyNHFuuWJzSK0G2PGBhji93lyG
LzSkzaar2Br/yIcGLuBKy0cPzNcwoZuVGRVwp6tJKnUvnP0zaGPNXbkSho5VhpIkqad2U7gUpxq6
yqinLVDfQJqPxbl9R2N+hc0q9HhExR2/mgbYYsqyyTBtiptGTzO0MAASjTs4pUuVNh3t7e8ESWqb
zddVxshznTJ40IFvJOWVaOuBKumFsURwGD/KIBclwSHjTsOnx2hAAiJv54IVj0sd0HfpJk1+oRc7
RjPboNw3baIr8bklWG7mht9qEx/h0PwnSSEn/nGe7kMhH1yBJFxgFCfUckfdWv9hNDd1PNB4R7WB
yKiueorzH5lWnkngmMqbO4FXvu1XuZEcmYFB9tmxnYmaTlE3aRQnuSEVZJyvXYVjaQfUrImX6NNK
zsEFZ/U2PBVqx+GjuxzqN2bklUardj9crBTwlvYq+vgIbFSz4DFKylr3gj14+fDKXlQdGUEn4sJQ
AuXsiJjgi3bmmaJbOV4VQ+ERfZ4qbMzwTVXH+fjUQhM09I79Dd1L6uL8h3nhEks8pr8Kt6S+UVlL
QfuGSWvZJINuboxWOprNWOFsNl1c/szH1e5BrI4Lk8SnbdED7WojNlXnzsvc/Tw0dxn5JwYpjcP1
s0R39ZPnqWj5XYdEwWZHdNu72WF0KpduF2cSJJNHsK2LJnmRti3+a6KgYkONh7JeC+kP9O48sosc
am2YP3WYT17WDhKdL0r6zaCYHmAtRVRbN+Fhy0a1BlRtnjYXR5hIP/cPrmQsQLfZSEpsmg389Jdl
R8rFSre/vK6sVgi6OW49p5u0AFVA+6J8Cng6f1RohXKLjxKwgVNFUrbmjMS6VvYpkD3L2018/A1d
MYC6QUkPvopKmTeE5bCCphh5xKBFN3wD1V8i+BOm/Ka5D+J4fwI57bNSvkAFtVpI6/cjM7I2BtmL
3aOyzBve6y7Z8600MiJrIsh8N8yixAQ/bu6jNCC3Bgwbp4D81Y67bTMj1R+CapmHtYDAEf5VZX/X
6l5MsUxUMfx13y0tgKRc17+pbmWVOigGW6nkkozIpMv86p0qnfCV+2UqSPEgdxl/MQXBjJfxH6KF
QX/o8PpNEayWBXmKfLBDkKT8UF1xIe7r1hh4+iZFQhgM4OT8Sd0KJI/bxytHQDtQPAyRVrUF49x8
QhSwQoriOTkSEM2RUg38wgImsrLI7PcXUrpTL9QyZ54cqyXaM+F27ww74KRyvUMxjjO0HMien09Z
O8aO6GSzErtUGBZlvnVk5CiIEy4Vw7tEtHk34NqA7pqSKCenJfhSfLNAOgI2cnHCIeQLjxo6cmrQ
FsF/Bj/5dzR/9gzBcdA5YzUT8gZj5yL4biBXS4zMs9JZPw9p3PDIQFwKU0o4A+ajYTXFZbjevwNB
bR/+NmfUKMzezlxbtwTg9TiVX+xUH3vdYuiJ693T+qAbpKokRKCawJ2y3f3Gb6dx3VQB3atJLQKF
nRhS3RRKaAU1QkExONOKMHr4GOiDCDD9Di1atA0iOwL8fW27UiKevNKnSa/paRrQK6Uztv5jMqSk
OaivDZWA4T1BTLwLPnOuvpmfXqq8TlNqC30QHL4gPEixxE/7fMWE6hOB43QZLy0oo8Bw4gD/+NNE
RlHJktrNeOO4pzWoJFgd6spEhrVybct9fOh2aRNLx64EQ1lZ0tpEoXGl+M/ixR2tSu55mB1kYO9Y
vKxF0MQSJ3cZ5K7syyKsWpN6Hx6C/FB1H66+CROyLIrfGv7tnFF8LuGtxKnmUzEYcKJkYPi9PXRM
mSOdJOQtlrNv59Q3u6dCkirzJDifmvd31W0ZqwCMFiUdUU4AvmmY5PuMZeIJgfpVoquAtDeg1b6D
xDa+5udy8kIg+IVGxoL8zCpUN3yvS4rd/6XX5wthVq6dpKZVgEP+fiX4aDlihJKhMCkhHrlikSxS
gyO9eoDQNnZ9rjxJ+8/RXtAMvB6TBoju/oE0qtb6KodshN76/aEogBMJZm2K+3+y4lemeORr1jAl
hUPyAmITatHk25HswGR/sHtqV9OwOXgxzv456l/B61jeG6t6PC9gsfrs8N5j1cNYZAJmF/37N8c7
R0YOsQQi+7IG6UU6O4048GHC5iCkUzb+/vkaMp9hX6isKoqjdfI5YLNgvDtsLTN2kT2A/grLbywQ
7IPBhwLzzh0MpaIU8p/iu2FMpc3/FDQNnTMzNcom0f9O3v8yQH+pCq5vmDhJfH4T0IJd15caOXQe
sjbpcKVBKtYEzcS4jxckbrK8ofKtlpDen6aK2+72jcnQKMPqVV+uP9MDzdgI8MA8nZ7ep5zynK1d
kAgh6GFZL5YzKp7PMWKgqZ7PAMXM2ulXlphu3YUI8Yo6g1hbH4yraEY7dVePf1aszlTxk6AvAjV+
JB4wuJQvERQZfz+FRRLvSbhu7Vb4VYMcs/rFDUolzKSy/qSuPmyuUftL4huO2Kk/GEWFIqVRDmUf
pE0oFP40g1WP6pJgHuRcuJJWO40/fvNopH8PLYXUqkbfriD5wS8HcuCm6qzPB15XRshEWj+Pv4+h
7UonmdhAqmVA3rxUCWJMhJcd8E5RJHxcLozR3e/SCuGvqNhxDwTHOKplEfLo/PVY1oOiRbp2FzME
5IBTzPo/qQ5rvMCQ1w3KECaej1DSTQVYRLRhRT4vL6ijOWL4adOXwcO6NA3lCWC04JjQbMlPyRnM
H3oZYlOYzDnXWLfD38cfJwwJXJkfu9vftmrt+PIpo1e2cKnw7jIZ472bpSh+xMDq2fvCi84KuWaB
OyW6htoW2RKg1kRSbXUZOWXXK4dEM7vrkOK3MIyBZweq/EsASY7FcDfmj5cuZlbxkHUc+SQ9IpVx
/8B5zA3JZaMe4+BvXAVJgiudTvLae3AnFtWvzoIKK3Ud3VWrjUWwd2jyZai+6RcyRq+CJ70YI/Td
kpL5c4ZLK2JHfdjVZKyRK6Zq8jZDf01DokjiJ3hSbemHVbaVzAqcXJAbzlAbESVEd28BIJzFp2Me
brD+aluq5y2s1YAlbvjUSdS7h2ARiOdWA8K1i/ns4nHUCMmrSdrrGyIwt92QYpFOnm46EcaDV/BZ
V9++DF/8RjnCmHYZzMx9poJTr5lH7A9DygpndYl/+/Dug/13Uxx5StjcEkbTKco70KrdXDeyoi/U
hSnOwC6MiWn5Afs8BqtGTITLWZdTxO9UwH3PZfMSdh6YlejsAZcXiRFbexwEMEAOguU174IcAk28
ghLdN6b/mCMnRub7/S7YJq2Da8AZKUenJJZHIZkEMzVdSki9F/Eye7mPgZvMNhZ1BW7fpP8HSm1E
7tUwq1vNoZrSXHWluBLJuqwDRPvtdr+HBKgNnGVFgUzeMUyAIHNboeBYTUgS9obnGUtYTw6orqVa
PChd8LeY10RqZRtQNC12HMvRWftmcD8oGHtZChb5+NPOUCTPMX3t5KRWXCrz5u+IKTISAfkFq7/C
wXyeV+SWRzQudUZJBLSJ8uFJZLSs930ELBfq0ZZMLNxghXdGqtw073uu95iWKgxLS1NR4v4FtJ0I
DNmTDfWJEwWujgVNGDNXFuBWhcnaM+Rq4PGo4dkQ8GG9IjlGHGN+TtuFE2ybceuuwH1WMUBdEK4p
3KOqsVSe16nk8tEjuCFGSUqc2Gm4pHJ0Ugi9vuM3aTwjS24CN/tehFeh1i2r/UInFXza1hntGQqn
JKD2BbVEnd0Q55IjWtMXPh4lLcRdJ/w3gZIqQaJb5tzmrCzPwxglM5qw3mtrkB+H9R9mg7n315l7
UtPK7MKq/50KBnwjv/69/CrjNkNWhwnDGlm8QdJGlWA80VIF8jwPlchkq/X4yZqhB3XaYHRsO+gp
RbEeB5KHDPZklr1kguLh9f5uHPT2WcDdGNCYCg6gPEf4/fW/ys9qnbg2C2if+y5LTmavTISmW1AO
RCN6BbyL/j19a/M/TyAOMvFhTChqtOPNRnlcLC8J0cZjbuOJwIXdwSXFPv5lUFZQp9R55Zn74Yff
Ddvim8zsi+hRO/HJGcZiI2wie0uq+jaa8eSpEevMwuuujdeyD/tYUS3M8DZt8c30NV5yuKL6aptw
gr6RUUJxq9XlkOcJsu9hoAbg0k0X74P0MHahWf2UrsYMS0kTvgpv93NdWBQbXubk/IDhW0lVWM+R
IuTr011wYU3+TipQZ32aej6QQyA8wkPw01Qo5dSD/SHzHwco09mxvRz0vgGTkb2wLLp9zc3LvmWd
MG3sb06uYb3ionOegW3gPWj6k2r84oY5samzKtkJHYJ0rVuJMXnBMi+T236TBgqusVIwpPI/sVu1
+Gc6iq1eb2vAvqLzbe7Gvo+VxJIMjpOF6siDnOrUw4sdwXZuz8m8VIkqwLnvgkHyfoL7khtCcX7e
cc4TalOpjOSM9RnM12x1PLcaVdmWFgWEL84flY7nbv9r76O9Hhid33yY+Ot077fqcjWsOw2ovNxC
QzVQSH2caYGbrPPT+/CSuP2fTNNH+PIGkHSwn2MWapFuRe/x8hkdF3z5rG1mX9THsyN87ahn+ocz
RKlfSQyKV00IsL5LfNlgiJt+RVAcpXGpR+YkIsQZDgobdHYdQ1m3j0nYv3PRrtttsajy0me/bQuC
oR1C+eFixfAW4VHQ07qW4yLAlYdUFJwdvZra2vICKrmIOOYlLR12I/GHU+E1UWnEhrrqiwWkGH2V
BoOOhpnsQCrkb/1V1lSjENTFy6qgJSil8W7tCi+MiTi+/1IYSSr6OJ1xZWdL3SiSRixN4uGox/Nl
YRFEKkg786DpIHeWHVXzCv9YX7lC/SVsv5rvTY8Wk/x1neVD/2xTTh+PcQtCd/tGfI9FXZEO0z0t
t+YE9QCt+kb7fH+9LYrZmo2W6Gb1KjoqhCCRe+a+AKcIXrudNZxAvHgZqyBR8s4ipAezSx5j67xl
agDXnvEq2iDstwIeBnP1OpnJ+ubRx/qpQcMXFYSysDa6Aw67HPX17WaIyMAfkpmX8eRtmuk3W97T
QZoYTBAglSzbIZFzGfks6oVLRUE37sn5BLamqeS0co4NWep4SxjhzWAmL6sOUslNulj9YCiUW7U4
GwroHN9HO6tY0jKjDkRPeGlq/RX7JyNTOhSrNbwRX6d9u+wRKxLHOuPYcb5YcDGyWf1m9KLbbqcf
ELKQ49zpH9bonergpstasmlIIlzoOXC6pvOCWQmCo7DX6IOm5VxNG3fWIWZZi6Ms9VcrR9mz+DuK
yF6ixA0QObeZVr+vcpiNWhkfYTMBqth0l624N/H/Ojr/QU33JRFJEuYhBkY5lG+VnlOlLE3EfqDL
xd9yPyYaf4AUdfNjpYQ32ofHW5aKHrOKXrfA6XMCaKT/PRhFc82QdXGVk6BhrO+9CtO8pDuAXT3X
9T1q77Q55F9COWOtxGoGNPiFBXOiPJKg5TS3clD2JTZsTWTcrfzwLlFNlZDg+ij0DLHzGi8jUNXw
tXybYjQzQyqvzWNj6uAq87dFw5wm90x4/DtCED1lehn8rH4JdBIEki8BJhKII1pZNNR77LoJ1p30
/jov458BygCrGYmkESc18A233J18LNq95JmtykKrd1nwyRELnM7OysEEgpYtWdUBo1rE30YljYks
+tM4hTZj8LahirvBTupvT63/JbwTTEDIurgMfnq+pT91guoJJfc9yv4WG22F8y7kyGVCYhk4isQQ
CBt0A+MO/yrvojRIiPnX5AJDIE60Cb/0MDt3oTr40Cpxe8l3HT2TKH5LNCNrmCbgXFOmZ7ANraJf
JweJ/4ucF9DKGxu15QaX9258Ce8cp2+Aq3qV+fA7Xkl423mbWGu8zDHMbtbTbcl1xWuF4ktT07nr
sn2FYe6+Cbg5H0EtMia3xem1JtQniKnW/Y+IbHkVvUy65+LwtnLSaJw1Oj6vvOlRjmS5i2APKL+v
bqpwhSaNZZaUMezGoqKUsMXsltAgWyNjLp4SphYnzsEmqtz5q2WSAh4XI0R0x8o5x3ItmsNH245S
VJRLh9DMTC8Puo+iHjpBsLV2WnU645206IBmLTBLQhEcNqvwJ1m8tdqCLjuEbEHxK21IO7IOa6fZ
/SRznrrir7caIT6O8Nmc+ZjUGSM48FOyEHLgGwnH0ysnR9Tgcpp5G6CcpMyMU0C9PlYinh+IA6kn
o/WTGSCVJPZwSyF/EcOfGDO7t/f+T6noaAKm1JBGQm2f7t7PBUGsbR7p+ydoFv/7tZHbDtXLCizC
qNMylcCIOn6my8WXadNGpuyfn+9tLynoVL0YsbPy6gIC2GkaKW1jiqDcZUo2sJrvD50mJRqjLpIs
oJqsC4eYIVUQDgsf7n44yj0MXnW4izXhNZbwMXlx0PZRzI3Sn8XJXWmYKDuOFn3hHs/FGwLx7AWv
DMSWvyROvB5nEXmXg0+XBNKzK39Z0Ag50xe2GVTJiAkWTimXhS8tAZi3VJ+urDpS5/KCU6AJeJi5
fTF26FmCSoSPXObU5ItXV6ACp559GG7i+1K/VTxH8zQJ805rGcISPEUwac6bWrUO2dS14oGA+HQo
ueugU3Rlgwi6NVdgJud9pL8OT20pn40cnz7zRYHgWOu1t5ADmAMGotSKyrmZz8HwRe8i0kV+vmBR
xEjrU7Bev28Wq3XgqCiwFl6et2uKwkaNjfLGk/YcClIE34b2V3toqOkt6Tf2ATqPuqQJD9o3qMC3
s1P73MdrZcalk0KQM4beMtKhX3hDpBGoKKBDjiGPgT+zy7OHXDo1KIkRbq3fVDEWOQ5IRh6Lji+i
c/iYXx1FQ2GTUSwJ+y3aSqVucJfsApSHHtEH2OzLsPoXfYGGmhbgWek+wed6gzxt46VUElMFX7o7
9W6HX4OFjdXXq8assTXRNlKGLXfh/ozYPJx8tMlV4bEWKb/rebttZCmzZDKhBLv8Gw6Xk/yKAFTH
deZ33F6pN267U6PP7Ua9ARsP2Om+ZrNr9xJSAB5I5G0TAGpqcZbmqUcfvEtcv2hmjWmL4I+ZCYVz
Fy1De4oe25gJMroEcRjp4exHO5f3gVsMHvIMJBmOrzmSvJUNzyBMdGdpx/F25wN/ajrZbV78Fmq3
5LUA3Mv5dcwmnkn65j0I2m/Yd2eQzzIWvkzO2zrKROYfsxqvTCf1qvbHmch+1hBHmS6GlMbzxPWg
wN/NqtY0i72AYL+roB/aW7T1D/cWu58L0ye0zjFLkbHTHEly3iiMiivsDoM6Vm0t+Nq7VVeaA4Pc
uhoE0CWENZx8hmZ+A76EW7Rc/BRaOVQPmX9FfFdb+mWGpJKbaItRCXHk4RTEDABU9XcZUhL3yKWQ
5Va3qsbar7mMvIuP09H/6W2jHK/QDI3ZJY/Qck1TtLJbxl/kZ5deQkoFhetQbKJMsmG+ZMYRyU4y
qeqNEgGWSMA0S6f2p1sME2qRnEeMogmaiLMJvBg1zyG6fSbC22d+y5KfrKLbYpiiHVWXjLOQ9m5U
MAuZkW97VK44mLmXRQvc9Agw3eXOVWYI+9S84uMpj+4P9RHk833IzD7XWOAj8CiR27vpygGbzKtW
DD2YfBz1XndF8VJvEe+Haz7m6UZ2jM87FuGjcMx/3GW8gMlX8uYfypN1pbf53DdbK/O2V2rA2KJi
3DJ+HgOBNAJgxE7bpgPhHtHj8MZJ/rDv8jaOVH8Mbj0SAo+X9x5z9DtZA4kmGitu++NHalSdaucE
6qFboqiijYR7Q+8sKCJhbSV86qFN9NtdJo/a2A9crIRH8mMBPzsvrRbjjh89d7tyPT36w0jcKHI+
qhSr6wYoPwscItX+Kbpg1iAG67FzHR3doJex4ecYv6SvTLZqkS6A8WOM5047ZrG5ASHYfL0FHAAJ
PtxkOkqyOV++7MymYl001ycSm1pouAgWEZZdijddF7bCRcPEbc7p6/eBoWgOnmTkKZ6IZvk+n7Uj
FFgsVyaZVuLLM2EAG3pgBAsHMjHCyn8aQbek6OHCAn6emQaCSupWv9MpNy5FSBDZx1YQaSkeJce7
fQ29na+xKTG5CCHmeKt4NrfGZVHPnmtMOtjj2Al1INQHr/k2wMCyk7OyLN1TFxPRLMmBNUVCJVly
A+jf+UA4JWr7ddKkkvgRz2D9BHvRRdx88zNRKViW8Y7Ui3VvvvHQ+VceN24+aqljYz3jO+nIbVoK
hd1BvMVf3HvSt0EydcWM7rFkhzVjBtXsQEW6xNgdb45ezZ0FGmRLF+doy14Wn4+DoG7SPfseYHNO
gKGd+QklHf1oD3k6pM/nRGmV6I8nyJyDczn62QDQxEJ3/oKM7S6NQ4eh+8dMyjUn5jRR7WPfr6ke
ofxdY0eVWACASe7nx6oexrJVgNsWmsyAjC81R7O2aE/bCB4b6egn/SGEN30uWOBs0iSQR55Dp69L
qOMVm14vCFZczOKDVSZgfEh6OjqSZhdPSs5Gtgn5vCNVJSZjNg6etqLmqYbffIw51zcv9RQ268yS
CnrxKqjv8tyKYp83h7JkeRDWXeOntmAsZ61VBA6v2RT82HycqpOiVUuoucKpXqJJqvU0njMFGLB9
jew+eNOAS04NFws+m4ahM/bdJlxC1ewZdr4niB40hS6aTgSOiq8vgMzVM5U/3e11m4wDK6tXe0Ug
KqYBZFxAh1Lr1rZZBNPSrs6Zbd6bMa5+lI24bcvY8jE1FlU7O+JkT6NmVokKD5irW9Hup3CI31kI
IFhZD2HenNiMYvcgrJQmrkPiEWoOOMmH19cX770FYuDcpbpJWdIu7j47hifBA7+z0GtR462KcOjU
0GbjrZSYEGvYjoZPOH/4sGLHzl04VrwGP0tHNbsheg4HwoxdDwXp8EvDscmjDj0CNr0tE3qFyQis
lIXFxG5lmWEF34qZIPgeguEkavlX5HlwVltW2p9V/YqQ62xgoXsdSiEWpDG78F3hEF4bf4JNzv4q
YAxB2mOTBfMMy+4vMiA6AdVLzit+bhOpgcqxiWT8eFbpi2JuXnvTcjZ8BC6pkPqXqCXvQ4Nlbo9p
izCosCFd3D3GP2QOUUJpQh/zzJNDLC3oX5anD4jfvg7Yb60rEMYeWuW1DYpv3OTSFst0BwCzFbpY
/VsvSk8PmuYaqKZkfL0oUlF0ChOxG6CyYVHmCxtsiVvB6HJ2Fok9QXgCrpLNUtBdTMed65jxAA0I
NG0ZAMPS6UrstGAs59Xa52uOZPAUZbTaf9s75wfkFZv9uviBQi0xD5b37FF2wrwB3GoS+a87KwvS
bM11Bycu4QJB1CDAqUjo/5TWK1u2jtSiDH+pO1MCyewnmu2tovT5T/0BlYOolrfJnu52paoDhglc
Dw4UnriVMZgto7SpsMjOAQ8rNYrdlPcrMwAv639w7y7MWondiFM5lxHD8sWwKbR+LGEdgDwQQoXU
YFy2NjdnoflfOEYDo9aPm87DNbPjyKJLpvWrLd3WW+KOZQciw9wZ3vmH3HWua8U82EyzYXCeU0zz
51K8wQfnntVc1cSblSaeGilmgglkcPzaG6fYO+sXqwfyEha0y6HI8w7MDROIo08Kzfaa/6NVUfgH
sGf8HKzHd9/yhO0915TYnJ2bQqk08a74/QOrQxB0XURV//v7vHYQQDuRHIZc5rGFjuUwUwnAnUnA
faIUndxOdWMHIbS0OREoJ0D8ruarQnNG8NjyxEM2HrsGJfZAHYXPMDy8ffrzmG3AOG00fbxPg6b5
LhA1nHsFPSQINg2GEyH4fb/s5EZoNYgO9XVwc6/A8cX4FXymNroccBwsf4gIdkFzVQYaROXCFGxg
uwo7aiCu9vOA77ERNtqASAC5BqMW9OoUnWAfE/hHR+2BfU7V032lM6dhsz0fALQdNKy6dJNjX9yX
z2V2NRgpU52eV8/tE02vU4Yx/BLUMtRNoOW0fENO9kXdsqBhdQGvY3vNB3ILb6rV5F8EmLmuu4xQ
w6RvNJD/hPrbU4Ceby7uAy1wQhr+JGcishkQ2v60Qbvy4uC+XVluKGSAU6DdBiuDCouVs2Yh+3qE
Qhqpfbo76akrqte0oVEKGu0ATASsmrGA00ZHPS6+W/dGgEUejC+jCXIlojsBK8C5XtaDRZacJc6v
SGnrLdHxrtTH5T8x7K1tJoWA96KUjSiqJKfUclDcyl5C/2rossqcyk/lbMWbAQpUg0VXkZA3grGm
1N9GmLXmdh0OX5o96AiRUWe4/D183smaSutoXot0ar3DWvCFaZ4pVHUmiE+cRfEVKftKXuQRX90o
KSUGwer/Xi73JaCqot1LcuXOXfTyA+vyD49aD7YUnfzXXNEBimsJt4Jcy2bZzSckCK0Z4C5Ra0el
x1DfIvKU9wy+USHG0nAwNtPxh9XO0fARsGXhXMLVmLacPfgpIoUSah+kkTZSeIiCaj62H6JkoL+s
gAK2y3AH5eqHk8Efk+7KSEdTHrfMcFQSYYLw6PeiYzpPMSv6RCQwxsAyikgJb4AA5JYAPASKQeu1
xugG+m1pKLErxqtPmE+vgVqyJ0dP8e63r376qILI20nVapgm08OS16O/LvXeej/BNifQiE+FBonI
vTHW0Su82HDpg9gf0kEBZpUZ5lsO/ybUSG9O6iULh/Ou4vRwElZxcVLCaeIvFBBscVXcfW9ib41D
M+jgvQEuWlST7a00HXnq0qZbq3xPcitpYSeOXjlJZjGfFYDZbMa01t5EZDAps51a7/qTnHBb7KaZ
Xg3hsvcWHyRV6cA/KWLb883keHqJX52JcbDEWNuqKapbNI9mgKzSzb93mycadKauVgkLoLeM5P3A
A6puMBjaqFWtrl5XP6rhvEY41R3cctfYkVO1wFXVw9K9Mho75X0Xt2KMjkavXgZ05VP5pERp16tT
/cbaMW9jcsPhJe5tR4hsR0Mn3FhF/mL3xH3Nu1F5ui2jl0jLIdMug+mtBsl1I8mKTgjJk+eGIwTl
lTk6BL/VUlF0HzsRg4CeLce7fTD/bGtLHmwxH/cebkpqKpzmjvWu9RCvEfEvRXTSAz09p8QlX8CV
X5baJ0xXXYbaC/KVVFt3xBQmLYHmcbAyaaCNRQYI4u/QTy4RuHlE+jPy4CawtzsQ+0y9+E/B/KCo
Gksie7Rg/nWvCYcctKlesEH1dajMRtyI01MWFGHV3aKjdX4JmPUCeT0irqsSHnFb/KOZqL+terEN
DHbJNMJz/GJm1CETSjnzGX8hDvkRZc9+9P5B+uOYKe4WIOLd/1Myb1P7H+psWzEiVleAgAlXISYs
t+WS17TZGLZNtczYAUQ7MGDyiWrYWo4nQ2HKODIDr6HOXbkTktWD42Qc+bDbg9YD4B3uJOYCgUC+
E/Jk7xGfmQV+jdnMKJAYWJCzdFo/kSk64aOqbI3RWFkVMwZ9jXISXNicZP/RGoo6oL5tQ7gAmJyV
6XBsEnof+sIyT6rJqeIJky90BtsJFt+VZZNxMIxX5bV/VE9P5Cy/r+BSmuwsacG9Q05xGZF21Bp5
dY5kWWLP++2zjxu4HQKVhI5bnjmIneYngQzQWn7Er0lSrjxoXdHdQhQ91fXx1hgU1fWXJoOkPf7R
/2Ctg/iO7kXIJMFomVBfdg2dEJo7WFR5LPIlpBMHTHb5sP8Xjmis9gZjCkFdAcYu5smiEQw/GU4l
MMxsDr+pY+K205eTMpdz/5/qLWu0cult8uRFbEvpwjv9DsAhtCSPEk2DshS/LUxL1TUiBwuDf5Tw
PIMTm10cLraeydaG0zQFUjTSMB9TV/44kA//08JM3L4SSgv3h/G6u0R4EmbOFlMcJTgWjhPX4+qx
+ax9vh9nn4rC5t5FXTmnMqgJ+EJTPJjEoxWLhAbfBGEZ2ory5loQKYbzGBXJERHrlt93fUKpTp84
hW/SU+U30XLffDweHHmr1Hd8UszY/TBAK19/kQdDJJ/Ju89zn/yUVwS5pddzxsZHBRtiUUPb5MJf
tch8lXQ38GKJz+E2zU9uMeddQNxPJjDiGbbA/lPvxKJzQY/g0H9ZzpQ4i60Y2clVP5IGTiHlwLvI
MywEANI9uil+9faHAFfBxoNbUaWMZfC+56SKoFOkYm5DgmO/fB2sAXfaW+fdHCBWir9owcF1s+rB
OKarGjbQbK5qDCE7ILxMVZzN2avrxyVCD2XnoeiF03p7kMZLwR0J7IVMNo0gPXbev0hB+efNgoJx
AoxERNH1grwfqM+6NhQ2U13V4pU0FVLsWMi9IH0h0lysrvrgleBDfbtvSBJqF4r04rRQeE792wsh
bXCtLk0cPFZbwx2Lg7QO08BLxa7Px1D19ZV/G/ddL/sgj9HcdyVQABxotrJf8L0B0UtEZsXBS53H
5nRnkxfVQBUm44V/UP1Mqug/K90B+uTSRcQv4cm6NM8CXVbwtbhRNRVNI6ZHha64ykaFgmDodniF
3Nb1YcXCALqv8bLj7CBt+P+fIIEOYRMaYXjiiY0OR8+MHW+TURZQF5jWbC/NetxYrldjClRiSLAT
dy2eCQT24+ZNSCKQslsLFxX8VbkQWuzMpnhXvtLl16PzsZ8/HWnjGKHRMIXeh3W349dpSNTL+Fea
GhhTsydY7a+ChrI2SsNF7LtwC0Rzz29izf74A+11jAkw+iasnAjUZp4dqUjrnYo1VnBR8nTtpTKb
0LNi6SAB7b8dIPKn1TLB5R/FD+pGJVubwWtExqNWW0ND6m0CxsTQ8+zSvGFgXWGZ1Kgl7XMpsvD2
0YViNlWcPOnJ6DjALB/F0gtTiQ1jAQ7S8lBWTk3eJEQG47sQkkt8EZeflpJOqpCh9sYagRfdvKpy
30CKmi6A+VW2Q3XVdmFXwB6I6o6JXXefrWbu17GCHzz5vcSdOHPhvUP6qAbOGbSdKqyA5I7GhHfs
v1cisN8Wh0Hxf7ddmMu+Cdy3NJqnbO+8rCH6/z0NXloemKWJF+wW8ad4S5LwPOqBeBZRWFz0ftbF
z2+Zv3ESKKn7k9h3HymkT0hHq59H8Nn2eXhLNHTbYbHEPJyzVMqGunzlvGX2e8WxBtB85lan5da3
MzUOiKWsSa/Wd8s3QLoG4xvObXC4/C9RV4mftbonvWIXLcuUBNzgBOshErYO2K/ws2R3sn3JYWwD
ULnQPRzY9OyRPzWN7J3IU1qmHTgAV7kP+JkPYrklDquHEDk6+tUp4HZW5D+i6M1ah/5uXuNVTRS7
mfhiWqWCYmzC7/N5nOV1sYUrlewjzQ50Kzm7Yx1lTqLJrhMFvcOWZmosDcsr9PaftAGEF8kbb+Bh
1jaXc62SRP2TYxPY/EO9ccxQFgKVMDSgY2AEIUY5pc8L+Lhe0PXq4Jr6UT5VGFJssGWpJO6hUuns
4YCSYhDSCeA6RO7HV3WdqpR5iY560UEgMAPgjpSlos4Z1Z06aXkVTJhs0qEo3KPFgInPl3vH37QD
KgFrufblZRFXOImydkDsZ7YRLxZcRYBeRIqDkZHj7XELgOKZAqf3cSdI608DalkZnJvu07VSJF18
CvXvmbbY2rEAdUS/s8UEKKtJq/QGkvvHzai1Zd66713Jn1GBLUw+r7f+EU7cXL/djN1YhuSCgVrD
BddTTTLg1Qt/asUFCzqWTUR8o4DAJUMDkGAhFnJ2zbzqeg9EraioG8OCS9eRrNI/I9Hvd/R/dJp7
e2qY+i7+XngbyQ5gFgcf575oTls2d0QDUdlDYcPTTep1Y1V5cW8Hi2iWyWRbC2TuwB5/nS80FX9x
Tt2QhFqVy0LYibkC9vBQ0RNCUxRXwX5d1O7zzhjhQmu84gUEMVbb+wINGVbGMRQ0aPHeXOLV4awo
C4oE+ZmCuX6InG5ntFuPDCe3LkzIzMMbI0XxlLuOF1hfNt8wuAY1SgbIGRp8aiE4Xerwyc0M4V7b
8FTbTaFl9ZVSAoBlFaXJHHb+5OuUbIZJs18f3qbnt++9R7X5qtDkl0OxT1a5LlIXHyVsgt/E3URB
65HnKpVMwL80+goiinKQKGPO6fFIdHhXDZ2k8ISLRMTosffDYA6EckeBixPM0+/9onmIO9yqnqjd
xD60CRa0eYBw3UZl0Ume1SqikyAmpEcyuLDzOO3XVMwIkKMyIxUO8LYOPXlnmjBLcTQQJVl9rejq
Qm4RME2aPYx/PIRLANT1Q9FLcQ1TrAsslVDBniisBV+MgSGUuSq6uEMMzUEmgkb14jqOMiW+na05
sKyNGbodgjMamlgeYt5pYwaY27oFV5z5VjMSacauAX3B3t330BTI0/C5kZGrXVVmTryVB+OkLk/y
jld39hYchPzXmQOxW2WEQEc/pIaElxu5tjjua5PWJqhGzcNJezThbJ3BhyMMrJVjqWNjOJh8VBVq
dd/6bePuR1JDiWuIT0TMw/k6MawFhyXP3anoVPXIavRVXTOg1/kzCIPlmFfD2WLai5mFzhmzB6wB
7OFedtroF+CyzXk0UbmDD/PSBRCG9u8Zgnm0ORRr3oiZ6X8RVOg9J2k/9q9SLatQDdgj6GKyH3Wf
1xQNBKNFmt0/JT2G646sRCYCZGKOWfrg/9DKOYxfeR03d9qWgNw1l1HOKXvjyMYtPRE0VYTHqxXQ
0w/wWWfCXvphSPwHl/1WWcUrn5WHFgUucxUvyriSQz+8WVRkGqVSHKqj/FztgJlhr5mooVUlQFyj
Bt+UdvxgcFAFocUA8TpZajyHBrDVTS++E7bJJ61Vcqv/Dw7XoAwFk5XHidqNaxOyIFEqA70Keq+z
xHEte5oeV3hdMMNHlYbvLlaIvjNjh6+XmQ79+r0DCsUquVb7lIt76Oa3wAYryrhq9JTXbm55U4BM
fqtq7hTkdXnSBEv+By5F9PR0FtfklAbbkz78DMmpswe63JC9CzWK4q699XNHspi3wRkt3VImkcEj
C1eQfnE552lrPr+OxUA1ceTWv2tU4PgVcJIK2UUGI8Os6B4KwWc7t9bq/GP+VGqaGEcNe/e4Tf4s
ApnjRuiYfg2UyTfn0wn1yKs67QAclz/MUKNlCX/Nq3SaJ3EbbJdc8Mi3ZVBbSahN1b+1ct1cyPA5
D6Wy09AMz39dd7HnsKc3ynXgx8cwwBLM39wchOlLyXYzdNeAY54T+sfybqJTspYm3VKhUeFon32u
vpzpppEPWDkkRMqRpu9p6wzbHJ1hvmdC1UrS5LKPu7zXiN0zjHwsIbEn40TlINOqkReFzZ4UhBxv
5tQWDy70rAlQBi+j69O2i8Rg+YL+06I1CpmmLSGDAHSPrcd8sjctRqI2WifhDRnQHDNPBLuUDzMJ
HenLXNnuLwf0coVC5DEDjOkl/g0oEG1Aqt65qKKeQ/NsxSJlcIR5TDrVW+gV5Cg90FnFPFYGf5Xb
+xFMuQawNpM6Ox85LmxaAabL0sZBrFyagKbGFM3j4RiMkfUHD1Hjhr4U7cezYxRF/viPDIl7o9BG
k9clCbBGlMDBN5YzXUcZw0wgvG44yU5m1Hly55aJfXIyOBn7dd0H/y8RVre09m8LXEojfv4Vt154
eNLwJSnaxLkbIPoQOqHuMxUxuBEyp90NjMVGnhIOUvz8DjTZd8l+hqlQZXfD0kNh3nA7tsfPx3hD
x48vU1TlPjuOVyXi9l/IlvIYRqTdLroaCr+5GLqwKMq9fkRFzdxVP4yV4vzXvQED7ENpxpAGdaEW
5QXViv9PORPJz7unl3lRAcy3vWcTAmAEu4lrVWGbiHn/xb1+BB5QvxgzeizgvkPNlz8TiFLF0jFa
3wKr8N0i28Pwm1YOrLM37p/CuBs1CcUUF5YXM45eCMhlspUVbWKRPdHBAomD5zW0B/BtdGGKHoxK
M5R3yaXP7oCsNzpk3ntOql7c4PcnFR/7oRyC0zF7daK9lPO0rMZmbNIpd7r7ThbVRSKEZkqynZyI
9IWRxhU7b0tmGt7n01c5RfQ/SCeL9k6AXAhf/SXlrQOgR4hVdJgYAf3uxvRD/KxVC0Ysh5VBr+TC
it6Dv2qpnJXD1U1gCraTZiNJwq0lVCfAmvxPd2JlU27qShDE0CNWHWpmtTsoZ+4YF/4xVuVzujOP
i2kSmR5HvklsuwN2WtMbLhsTBAukW5P2Wo0XqqLAuRE4wpcrN8dLc8Iq6058eWcn0Bmqgnhfr64R
vtebliq9EsmhOlRd3cgmB+DD9Rz/65T4ZZAhrhrCXv71RthVMDAWQnLWvXPe1qGOMHt1TgsqNq7V
tK3raIjpwreL71aDhUClQ+UBGdOrHUMNUg7fx8CPcQbVodxobnqpRnmZh8hGtZUnxblOm/jgCj0O
8kegXgOV90AG1qLI3JL2dO4pwRi1JWlw9e6s1K2Uxvz/bNwID7k6f4KUZ9h5OnbQRFro4WCVTZ0F
loUQxjfv8IkE9Yk/fSed66bMxH2Wtja22ayHtlkZPf7Q3Q4R1Bjf0B4Eav7xg7y67ttWY2dSNWFQ
D7MaXDrcbbyT1qJsahn6px95j6KgxqLlVS2vOGcgbPmQcQh17tZ8CGiis2zchVbNSalMXNIf+5Mu
16vtlQvK5OgY9TAUEYtKC+OeJWAVJuXPG+VqoHLzlL0Qouv9J0O3cVVHxrRsAPLDCaIvBav/XVzw
t4HVZh8XXj7ScoS5vYYXscvdgJkLXjH5uwjGvrk8zN2syfWTXijB+VMMf8VqgsUV/YMovGDof41G
vl/ce29m6WCSnVKFisdhGlVVXhIMQnoC/6okY27y+WwcwBmU5l75lgCXIZGM5eq8OPyL0tOBvfxM
2MRfOLOtsEnnNwvfTW0yVEjbk8aQ2qscd+Ex0H1EaOBlncaiqYRXhB/8W1mBdEA9j39M3kkQtR/d
KrmjtFiezNFcVYJhtEaLM8axOPnrkXXSy9zUfUDaJB8tejgHwl9VNf8PK3nZl+pLuZDGrYmlsbEp
NcRAI9iHNfFyc1FT02vpyT1f9uT/mZErWrAyi3O2DNOvaY5BzEutwIotfBYAygiKCmhLsKFaPZIC
/9lW0CQBf4GGIsXVw9t1nluC5EJrkekMkYO/80dGeGlSo961NkREHmjdUJ/tdV9rLGDtw68bOi9k
cl7Z3Pq6l9MTP6nZsqOKJs9A+/GUR8AS/CSaR0HadfREU/WRA+zZt0XiI5ABWY1E8XDe4fTSE8Ib
LcKxPkebqGjzH3mUUnjIx2P52nX6OBV1g5GQl17o9TPXiFdQoU/eTQTKhVARagevlzCn6aXk8rEB
sfatAkxjBV5Y+uDqAUjvfravr37FW1ou1WimtX8RCCq5Y92ewsuUEXCcadwcLDyYa6SWhHxj8hxW
ynoZph7LG7qhoWf+D2Aa3SsK01kkN32rwRyE1xhODqG+Muekfo1Y07CXTcPTZH1Kuzve1V2v8UIR
sjJASKwgv/MWZaJcP6SVLh1tMXkg7OWuj5u8PwOeB+xtwI8p03tLQuN7Vly47TJkj7MNFWJNY6kO
fysQhhSlWcU8MxHhpkr3pwrWRfSOwaKG39C30LLwZkAuMOSXJnbnJFq1S/pdqQoRCyIsOYnH3tYA
vmxxirzPkVU/WHadbQ6DecassYfTVczjEgMbH74pbaH0ESFJ0rp3cwQ2lEq2kuu9oXwSEm2UYYCx
HYRtO66XXDIlkoY14JO3uiphffFQb3Na4fnVeu7X6cChx5PwIhYC0G+22v7PU50vEbqu2lu3a6zh
tU1cmfhnFwlImc+GhwYKqtT+si8ud9JBsCBxiRvH6O3bp+MHNG7EV0lyah2S2mHw367JlBd34aSL
86vB6kEtJ2P/GcgrLV7T9j9Wl72vvc6snAdktxZThGKqN+ftiPN0vWVCkVeBIb9c1l461af9VKNd
4+ekPxgZ8kzC5/sVb9QK+MtvsNdCFjfj0GbO+3keTEU69HPHOjYmkELOzSj4qvQgopbsoj92UK7Z
OHzwhjBTwV9KLdn8DQSkQtxPOQpKtLlfMHxkz+CuLwO5WfnF2DfWvRX/kjXEReRD3YKYLAeiF9x2
LAuwK0LlBNEQkmXYlTWpWqtnhLynwLLsu3F3EP2Y6fI7MJUcJ6enBuOOLyGidsTL6bw+O4BzFUci
327fe5i0a+bjYMISYxUqKATNPcRIjXabxZY3SYIsTVlrzNa5ojH9OpvDEaMpEdgYiNka5SvZrsVY
ntI/x0cRUI5Cv7r9NxlDnG4D0sM8N3ZC+e5G42pL0PozvFx3DkFD09sGbVnjtJmDvgmubsRxhhWg
zHxc8qwMJAa8yPAOJIofy2EfGGgRh75FpTrJbJY7y99kV6tNmhwVtD6CZtLiMJjPgqp+O1LHzvhm
qXCJxgP6s5CB2sXIqfUNAZu3HfI8lOasKxD5Rfg1ZwgSyFIDgDiQZF0YArplotTEJIi8HQsUOmjA
gz5DXUJ84yG5WEaMVu4INVZz5EZPOSDVF9CdAREZzfd3CmGQ65aixwKkGrCXljKYxh1lZ0Kprrpk
ZTfUqNI3xbtg30CE7GF4/D30k0lrW7P0Xm/3m80XIPNQzKBG5Qa6wOQR2cNSk2o5lN6Jua+LNhjM
4WwdMIFsz0OTOrWOC9KEa6hCdrZeVL3P0U5aAL1RNr97s5YO7Uk8wd74V1Ej/gZjaG9cBkAgYXL+
oQGPZ7ikChh98YAFaiYUnU0C6bVOhZbwa8eA+wz9+TnolbV7dBemahZwiiW85wm074d1694YfDkv
MjovUOjzMOkTvupC3TaBjqY7td28MlWnyY+LS37QpQH09YoUpalaou/gOWVoWwDmJv/Xxdn70LHW
rNK/L1FrTLdHCUu4bOp/no2g1ELw3NoFKQjeDnziPI/a3D4kevoAXZY9ToAXpNTQcA+BjNFAiLy9
HJ4YnWzGOSKZp1Hq0quorjqwMJV0mcnkbfzhYWuSg89ULqLDV1EGaY+kx5xZbMvsw2amubYqNPKh
gB/PAME5axCDYdno6l1EqpvA5uiZqOcbX4aQr6ocbn2g7OdXGxMnIoZ2Y0S+PFtncvtsb4vb4kYa
AugNKpp30Fb+EBeMT1/pB41sdMqt6buwdXo6h2gU4h4Zrdexw9Zk/qSfqjiwLrEnJZPdOM6uK9NB
DlfnPDJxAbaTcNnFdvQOEYdrfMN+EdyjcIdwKWi+AYUcLcuGcQYnIzVEqXsnwmTIp2F2OSIWhpeU
HazBNufizS1CcL/dxAvye5WyU7qA8Z1gu1k61JjqMupCMz7X9NNg5dJpXh42jb7Vq4uuQOchYmQT
YLQW1Reg2o/7Y23in0u84Mv8UszzZ+jsfxdkv3zzpCj8KJsvLjlPvumr4T5YhWH0Yq5KVNik/V3m
jSDk7JT1c5LuXmjeXHQwUmqwgxlQB/evvbdJT8UzU3VO9hn+49GnwG/Dzvt/cvAvkCi5gnxUtd13
V4Xhgme241cAwulkQGncE0db0zPUNFm/XGkKE+46MHvyA9YE2DVUoqMc4n+vCu1c6amX23tISGpU
CXDk/Mo3a19pAW+f4zPprvwa3hWFQV1A6t5Oj4YC99uUlfdq5ooPdc5XZJCf4Wz8avPwus6dWrpL
UfLWJCbRuyNRrfnxoCaRShnWOMUQT46O7QV4nxsoOLVbT6qo2O72H6Cf3jmUNM2HH/HqyoqdJ4JT
NGiWe9ycx4CR0O666JrvgV15Q6EA35vvoY1/OMztJbEuqBVa581MPQTluBW0Z4YgunZpH8oYIXJB
hFaWL5eou868DrfIXG8m3A/B2ljJDoCNiN4M/hU9gcx0ApvMrhmSdkLCrYm2BIcRvx7EB+objIWz
sHBix/sxriCBk4hKGolbnyQIgQRFO8+XbIbo0qlBI4J4Z9v/p7HncIMUX3HtFWVgvbWhhRGemoen
VXRvMy14h+QBJx/KkWkk8YnwC5zWuYOiaFwV54JH/ZbEhQd4h1MjGcYe86+DvnLmlgwV6WLvZqZ2
y5vRsg4Mt6N748m7tYskQAXzfhcE0r5OHxAJZnK6NgTpKQukqdmEsF4h1qMFKWLH8xPsNPLgQ0Vv
/izNAM3/tnkJmhr8dMe/VvOohDukoifv7iimMncD/azcuXA/y3AqxVKF59qOGEzYosCaoJWNB+pm
XlLXdTCNe9V/yYHoaDvCnypkbsa3K6P67YUC6La46TJ6B2lOKdWYDimB4q1sf+DSNgCcURGHu6tR
bVMEKYV5aMSbyKdM06nsClCICYW4Ca93hn8BA5XMTCuJ/9AofKADMjjr3WQ6bJ/E7Q1ofmwn1843
Gkp/TdVHnVQQBZcWHXSOasu89cf/2r5K4uf+GTbTDo5SgnY+hxsPClaXSH1LWL4K0UGTnuuPh9Bf
ayKdHY+TkMp15B8snNYeqIwm7g8EAU139kIz9X36p4nzn/WmB51dwCPy3RmTWYdH15jYBWg1/VjF
y52c2SMLK8gAnHCOIDLXBfD+qCGTCo+1jX387JFcCN9C5zpp0CO0Svy3j5SAjY/8B2pTF55qi1LX
iQnTqZci9u8SFlA3upqEcq+Zl2jyA41LQExDc8IRPsglrL7SAZDvUnEfODAJDmVuKqRjskRM0cWR
MCZDmexdxGzls2+34SiPX0G1yuvW2vtvLA7/YmmB1C5F7rraPvFIvQOk+6nugemPloQoO9iit5k7
RdDpAsJcW4wCl97n9dIdARpeJQKwn2tsXctLSrzPzRVql4RFl0cK1cRrSZdGQoXDu0XN89Srhmll
AwNi8hQ13asxXewRriAASJaCKcuWgPaHkQp48tDHXYAECJF+k3WI1RhvMtbB+Sp7Myk6M8SETavR
V57ZcuRgEEcT754dw6ksXgZZ/FGGfeEMJLrRZkrLe1SHvrKNu2akruYKmHE6StpG0dmNsKaCcFNx
LNGnRFvECUmzcs7GnZRcOCN5RVVsyi2diGj54iS6jhV7qep79x7OaSSq0W/zyrXFblyUe4qJklz0
2M1Yrw8bl/GvXpmKDLvIY/mS+RlQhVPqsccGb0jiJ5c8ZMf5LL2vg+jOAZe3ysQzF/z+miV84xM4
54r0bX3K3aPeUC5FRChOHW6UGLEMnB7ZT0T4eQBubjJQj7ND81z/2Mi3u+lL/WGnTCAgSCxNKFBp
+QD1wM2lqZvz651IIPY8du+jLPlaf0bAr4oKzMXjpvGeaTU3WqakyNgy5c06xw+1QfXSOaQHIGGj
jl+vifwPnA98ON6EGVl74vT6ljxU6ak+ecUgzN2LSauvFki4p8rdtfjEx81ZOjkNhBSJXXyqpCpV
x18wDnv7Dkuf9QUaaMP6XSNMncY1lvMwDoqj0hiq6hPZp29bJKHUTg+LYJHGZ29AJDBhvNSabog8
r0TxkGc59ITJwhQtIFPGngjhsOqYxr92yeNEgKAS+F7UAuBqiXDFYXPPHyVS6bwRZFHLQ0R0GB14
NQrFzYrQtQsDTur7P3Qyma3FJeIf9tv3k/UrxIUaMBEVUjRa2msb331+iHb9ZdEaHiHjxSULmTbj
ploQXgnzLdHlHfQptXhgNsV0mXIBAI2NTCcIFLDDQjrkuLMyJZhm5nFvFhMrlYtmgKZJmCpOmbLJ
GAlYqy8eMPcWb5TWzXSsmPhFjIfmuT0p0dIflKUpN56ZPUAKrSNUXpTz+yvbLzcETcqRnVYe9ssY
lMDUN//L9TW/hMM5fDCwtw0a37A1sfX7wpoqvvty+qVDtYbkElCaC5Rjp+1ELuejMOiOlmxAba7q
FqXtmfd7Ta9KpEw68FBj8duZq7wQqqFqeulE2w/277Qg6B3htPKF8TyTTDfb0pLPiaoOVxOcXkU5
8hOiXLSWMfOankcnbryhQAhmJ5Uu2gPVpY1tog9vcUPQgjYTTsjMiqd8dIjwKMlJrYJJWfU1OUUQ
u/tqeTJHCXYsgU9Ev55lYO/gs5j2pkRHKBZNwNSSy8sw+CWXeWrsBfogYUGLZkMZGdU4SjwE+vm8
JNndR7aaSAXur2pXHD1hdfsfnoQ4yx0XkRNAS1r7iYiz/VxV8yO6IIGY7SHi00aBiHvyqVH0TSB8
WzP6F7ZFCdyVGHLyFerCtAwvHtFAiuZeMZ8AE32PUVrmPzfI6WTNR1ANswbnv4y5hNEc4Uiaaa4L
MnHZ+qQYd8jJMiAJmRT1tSmmS2A6eL9GXs1eCi3LKLVJhsr0FAEl0dCa9Cr8ZCo3/GFYB9bxWkrd
1IpIKf4h3KJnyJShPqy4DKz99VBA7ifZI0zS51UqzSnsvbw7wZLqiTJ+kgS/8NC4c32CpKfKjiou
TPLSXwp/a3KvwAgSvsCjiQPerj7gTnDgP4CJIJCEQt2eNEvhZHep9pBGBQH6JHZNGiT7CqRuCqlj
PpFiuw6atD0+uWLW3aqB9qAxdSYB4Si/VqJGsvkh6FuN2Azdtnhxftc3xOTPyaM8rHCvfgjAM+H2
lACUDjb/zrFR7B96gESkQSms/1NlmD9mKmc75H44Dgph1Mwc4fuKpdHGbtviUBP/EPhiYeMr87/w
MJgnPRX3H7/NC38wBgLa3eJtJubJHtEM0tCOLsNY/LjkbN3F21SczX808zjtMXDxJSHyqzpJ3OCd
f94w2Msxx+/wM0R9MkzYGQy36xfDhpqDDHpbZYuIaQ6K4cBcnppFIU/nEyTPE93mTkzGJgYYydfm
Kw/lYKqptdKL1LsZ7xfB7JAonWXb7RM/ngIZA4i+s85NiSVolKF0lbUZW3/LtOKG3IkZjjhYdKhy
gL5POPrZeK5m0LV5S6F10VoOqRNxSymh77U7HU1AxlVvc6pJpSS91i0muirhig+5CDTMYF0m70QN
Xy0o+geCNDeorYqZU6zCYR4yKca3weVO0Pu9jl+Y9hvAu9ESA+qxyIrLH6kHLjTTKF1+gcDW1XGy
sfFyv1Jgy9WMcovyjYTrMHDye05fh9hhTuz+20SpQlFwO3e7YJocKJsLQlL7GAEK21x7Ki/StY0p
jLzMINUm6K5Fz9E4ZmrQbIZZjpwMIdXG+m5vxFZVUR8dg6IHB0RbPSKwA2Qa79NqDL9qYyt+xdaJ
sG556EcIn+eEV0IouBVJhlsABOsUfqOGkawM3z26SeNF/Qi9MW5NsxSGsvRv5l99VN3/LgQT/7KF
zyxH2UsDPR6TYUvPFxPgakcn10HYXY62LRtzr/xNQ8PMlsXQsNo7qLAyApDCLQOU8Mc92MByIYO9
hV71BwKrNmB35iAtZ92oGsLjbzWOIVbzQ3dG+ph+4t4bdUfq2YW9Ff3dDLOnYxXxORcSzDyPuu2U
TzZCQqpbBHFFAgJtVyqt6tniVTspsz//s1EFepirfS8PTSVSJzUrLk+e57tuaCkM3D0LwGTjFxwR
cZa5m2tRYshDIbFYJio1ZlEH0dtdI5VbqQaKrCG9AJwh+0y6FrazWHklt0Nd9yT7AAnhp9eWKtab
RJ/82jdZO3TjMisc29ysfHXBJin/abkHkKYVqWwr9Jb+6enisBaC/btVr+QMiBgozy1YmDQ1y7t6
wE5OA/mhKqkZNWS0+Pmrl/yhC7t3bYW2Njosle7/5UW0prVW1yCKRyjfZoXEYCyu/YvW6bXP4x8T
YlCIkKkUmrWR0QY+Et5+OG8DQ7dCK/SLz1n+riCa/9PIqxhUq2D2SJuc3pBZb7yabNZz1CyQJNlV
nDL1Yl17gzEbO+Acp+mAE7GQ8g5JlxUr8be5HjPlJL4mEZw9Xv5HBHRANzyE8FWO3PKCY/jPrf5k
+oAPsJI4qrkoDaaRJ4Sp4HOL9ep6MZ4gBKq0dPqGFBZN5d0etb238mmEwBCRjt0jCch8lZSiTjG+
eirWy+nSmFU+JSNV1+yNiu8mSLGgEClZMn+PcqiVbK2wluZEQzpCZ3WLw0OQndUS5POJUTw02/gN
u97CAfBrDaJd91j1mD1TV4fK8U9VPVVTrZG4VFUdGp3oBGVinoN7wF8ACk6P6lsLBg2t9OGgz2DQ
TgKgp69lBR9NR9mtcW/5p18A/VG6vhRpkZMWtdFLFYviQCnYAwXkZOnJnGtKBX6ivDMsYUhgM8bf
8YY7oRF9MFZdYSiuecuZj7DfDLFmR//ByMhYw0MlWaI9UgTAmXr31+1WdYud5tSpbySZOjBR1IGI
i/jeD0k8+FY1QIZPj3sWx7Q59cP1EL1I/HxV9wBZ3L+ZUq81uG/7SL5TGhdRpA3MKLezIucwEid6
bZoklDYDqv24l+35tFPtSwONHQysfqsbkZiNLU8y8c7CIFabO6Q8650r+YR1IdgTi/vFIHoRM4GC
rFBEzqUDHHJv+TZq7Vw6ofeCBhfDLSE3Y0gxGd2X0GckX0OdsPHHntqHuTFJFD4edDEE80HrZIP1
dmB8y26bWOzGsHDMuuITiQPCmG222YoFRp4xW+hqww9copXmh7fuXb15m7CQxPwFHB2Nehgr7VaV
2LtIeWMDvRAWo+g3SJZezgYMPATFl6F4wBVTrXcZKohmXDBflRucKyJekLrigJvbCQOdsaQ6Hygk
lLdrVvN6TInysl9mE0+OXVYQrECRJEhF2Y/e5iIIy5kzgsOIPvaeixlHhHJofzE5kiu3AW/9Qr6b
3SEkubbhOBZa2/oorKmVtQqnORDUsGaPaVxlHSb3FqKOkzMZd3UPkAOPiUJYaHQ0Jc0kQe0FaNsX
ez2RicykmQx6ulhUvWs5Bx0GJmKuobyesFua+WSDwlWMQPRKkawldgkhSPN9uBB4UcyDuvvfGu3o
w8T2bS8+Q07D+1EzIib6UJXrz5ypVRJEASXbTVn5HfXnFKspncD/SMXIwmXIznQ65TATwVtRJfcm
cXSKlfAtYrzzWZbrkRvzO3OGRRsFCFzkmyk5a9CMJLuwppBkeLnYO5Sq/QwS9DbqpZZ7uRdIhdQC
MIrwrJlLWIDG8f53owXtht2nf/wEGJNLBXcieBYB5xJ+EP9Osk3leh2YY6OLYgYtYQsoyvyabI7e
w5WpdG3ryoagW36SbplirY+rqkKXiKscbbW6B10H8Q9O0Jkhdm+xakZVWhkMogenlgspIGEksV1c
J/orNG4RhctJJqlWSj/zXmW5c3BktnIiCg4eo/qVBuFGAqzZtDg+ZhTazZeqPPFnySc9RU+SUsS+
MFzRbUhtyIIPhF+vecxolj8Ec4Z4uXHgON+zj4hhUHVZACbt3aH6jAKBvw67VGKCnntCh6kZAdEJ
0hsf/tndXqrsYMqXNi06muaKxxUYHrDFCNRZ3ddkFyyF2xCcizkCLSE12n89pRdcgNLTsgeqz6w0
4bOdolcCTXBDRkKZS2Z/imAegdawUic2Dz87fzo8phqIqOGrcoIlRVkjakWFkZSAIvA2flQMUY2M
SdJTm3uKs8ffxjqkb53CVwPyj2ASHSsiEKISYKXb0qGF0ZU3Oz1vlpQ3rPGLnDHwAzD9FMpwm64N
lmlnU7a8IqRavTQfmFG5CloiRhmmnLO8hvTM01qqgI8IOSz+xdxyYhO68+6GR8WRpKozsXPVrRLf
Ezqq8d4hoveszq0Cqsy0I/5oRBAiJuARk6ZtSquA7/jJQWnBq6lPs+RANr7pmoLX0KGYCMVO7vG+
qi9y16idI2u04hEDBL+GNiYEj57xqP0GbeZt8VyHNFPZbUpw5EHMFHGNpRnEa4ClGCnHFTVU/7LB
42NbhzRYvFalEI5+/u9k1sdK03+Z9HXUZNKPltPV4FIAbiWliB8ykSJSTiMN9Q7er64PFnl/DWsJ
EKh+KBlhhMLeYcUBe52LgRgPt/87vsyYVpy4TavG/pQubpdXKKm5L99UF2niV0sI55bMitX/atXt
3nIkfja1yMDck5eZnKQOMBDIps02dgsEPfCwkMJ7MaqsJv25mdOYw4f6sV6KgiX1bFjx4Fl3FKD9
9ryAqL6Lye4qqj1xe7IfDDsUo6oQyDDWGE8IdT/BbuZzUvUDvXk5qazGxyUoyoD1xUWGAv6Iz5ul
ja4dYQhGandCUr38mlf1dLUMwR6NMG+j2iKmCyhlL7kDLBRTp0sruQ/zWWcPnvEBTq8JMPGkkycL
r6xc/w+iaVgmvyxysltZo6BEfZouKkwGGmWsl0TSm0eUQqlvM1tSVS5PLHI5Vu0235i/s8nGqlQr
Fjv/H5RgARkhxiJPiKl1qd26FqZj5Qi8xLVwQKC7+7/50/A6OKA/ZgeixxTyHy/AxYIDjczWrX9q
fQi5Ds9iQi7QAnRl7HVuLtLctr0CauA5vG4pAd3QQzSJxyOXo9ukwYwFYt51ly97faSSLpujH1FP
8rHsBnzwTrV3cRjXXf9uZKXsBvg6I4DbHXNXqqpqc6IdIhNLux4VQ/qTG6DErYivv0EO960Al56/
Uv1gZ/G8sODHzValxDoqMZ9kiM0sfH57+3v8zoiowpZM6ivcLPQkWH+qWIrvWitdw399KQgsnyLW
MNTEw6SWPV/3ng9YLq3k0zU8qzPF7XEpy9ZkH2uAFywxb/mRYmJk+CEX0zSE5ZDZkJwYbxRb6ETF
1uir4D2ATcH76pg2X5jjcgNb/E8GhqbbDPR/7BiPDInOWD/xztVks5ZSNez27GdYIAjWY5XHeuFS
EO6JBcpTDFtX/uXwlUfUrt2OKdIPpu//84bI7n5luEzoaBwM3kYQXTqdUv5eLZcz3OVcLLaq0o0R
QnR30RNqgoWE1xccNadQgD7jAZQbzasU8FgMa9xAw27zqoWkgIRuUodz4FDqtYjCE6xdvjLzwflq
L5+fSU5xYylFeUK6k9U30z0rsHJm0SzTsBLF2T3XIwSxi5jSYF6rUVL3N9gJekQF8nkWoHf1QbpX
IXYF2jrVQFNNW6CeCozu4BbvWmx2Ut7tT8kO6Ts+8cd8t3Y4kuCrhFC0A+mH3m+RN5FwIdn1lZM5
q/d03TO6oWTbPakFOZB2AoQpR2sOQT5ToNz592XGiMMtkHRpU3Wmq4X7ibH6FyU1jTYEsP9Qdxph
xbI35x4LoAljdurVsuzaApseEFHxEILDZ7M1zcfpG9j6DvU1MkP+Jwzi7j1fANzSgdWfyHUsSR8w
8BOIWUjE54itQnsGAB4PczWV/VL7Ttrygq0rZ6AVXuwRd1fKz2+pYb+KckdYi/WrqWe6gckN1WP2
2GkG4Jo1FFdpKgQ/ZqyLA119YUe1Y4tH9mXW2AEOhNaFz9S82KSwaXFy+dOBuCFztJuLthswDLpW
7DhwsJ4nB4B8xfMEq/wkKI9jcSMxmUMfX0nN2cZIKu7Zmy6rZm+xR5hPslZ8hcNLeva11LKET3Fc
yCSHzyr1dmIn/2nuonA2ZE8Oqc0nKr6yLsAoJuEYDIbKNRir92s88BVHlzrJAmLYvSQaoM7/MpM1
sSTRVXxp9Q5IPY3tJRoavVSWlgQadnW3fgT/b4dBvzGYBdIcyAdhUlGeOKDeNjfhbkHKLqYtRow/
qtrkM3bpdxxjtq/Zloo0BMobL2O9aaAfFCuCE3Rgxzf5y+S+IDDOieBvvM648Y6uRFHEAe9+evDt
9q+nVh6ZMCEUBbHPv04hELa7X8HmNo+rWOazpN273ElkGZdlmwHLpRMrd56XeATsxw5mUe9I4A+8
w5O5viz9oyG2oYcsVn53iIwc+BJMI46frrFknMF9aa9zebyxkdtYFK48fFXKBM5lJ5AIxdkA9am+
gAs4ISeV5wIo0wOtxO/8iueV6M/ui0DHSL0brEvS7fbReg9UySeInliK/AMdqwg1oXAcmUwjTjb2
cc5pVEz6RF8jMhfmQMaQTej3TkXiAtGxlHwYSdq6zSFiKpzMsVkuUpfNt2mT9f2Bj1qMCX7g/ZLH
lMratL6P6nc6yPUOZsdp1BLnBG6h6EKghaqqAKpYJfbcDZQEhIY5Uc05HYBqto2cApa4YpZP6+Ek
5RxzEFIlSFNpQkoFZTPTAaBYOTBA6i9R8n2EuBA+P1wnnAvj0juDhgI+N7+cSDgG5RxsMBDeqq7R
ArBJHkWS4BLolA6bhgYmP/7tM7y8Ujgmem2SwnE3LFvI3dPanGnEWy0Snlx17oYeFxY2UkYHkAr9
w7y4NMkL2CuGh0/x5VpOBlrZ2sFH6KKnujDTlpqKaJ8lV/ZeAv0eZxRAnfmUp2op1niTHTWLd8TB
a7+3vXSHLGBXIynvZ/YrFeM41mO6SHLvlbk5fq4Jvt7GpF/UVWlCs05qJkRbZ6KxiYUAIjO3vtmD
E0QXy8EHus80YsMDxOFnV9149ii1LDKyC8VsMzTjx3FulwCRO6sOtEKV+XKS2q8VJGOOS6x9M17O
e+df0G614U3JJjUqLStF+l+8RS4dG9x8PMKqCB2G3j8o6T8PLCjz4I5zHVbMtU4LKeDFS8G9d/x8
f0BTkT0zY4iYADjnmJtN1SDT4kTP0A8xdCOU4+WNpHBfnlUT21WSenEPr4xHlzqdKoPTLuhcgEA/
CjykLos77zt0GWZ+c7dsQQCePNbhkjWj/C/ZLIGAEWWL8+Qc1ROQvZjSJho5YWde4K5+07NQcuL/
f1f/RWbTaBoTLOhdfjebbpcJdLd8iyO0DLLYfsm6/kTI6a6Ac/s/GWCtgfMON7XOZ4uJKFSeN0fh
Z4bIKuFtWUYe8SGiq2fjsH/atH8y9NeV6Xm/9gBGhjW78lXi4WJDu4CZdGRbmoJgVmgBB7hJgiaX
g+IcaenntVkDAHaRw81gZf/8aV31+Q3LaagYmVMUhGC/ZDON/f0wAR+QVQQjHEuqhOh4mxe2aKTh
nvnQyyox4yKlHzD1r5rnoA6kg2tc4SvoLm4jXbnTXtyeFiPUFfx9eThy82jYs1Iqdtnw6oRADhVo
t/sT7Qi5dp9Leju+DH+L51Lulff6nizm9/3/COtTpYB39O57+RIwCoM9jrp+TxQpqIpEl/9n5DQ2
09U3BbHhOOvBbVA6hf1KTvW0KFv+VNe+yAvUe4x4LeD48DK2oZT7QRlo+1vHNxgJZBGNOUH8e0sj
lDlC2gffBYASH8gIx4E84qgR7p2k+potExF/AYPsQivWAPMOvnzUNeHeVpt52iCymVhdFN5Nki3W
/wIvzrhcgioHrO2Q0TUaqodz/Ph2ug2vMBRPrfbAIHkEiKYszAVZsW4k564sprIfsXFzbsW/1c4m
afmPmDRKuUp/yiWBgn5+fvK7RGP4wl5QSlRJNXYttcZ8Fz6yx2dM64A+yDw4KMZpfsuGIuFwaY48
456fdIXHmfDpu9TF98Od0KV/VMZEY7QoaQIhtzMnpWIEjuX7StYCa3PGrj6Gmir0x8RHhx4asTwu
zL6f/TvB/RROsyGAKc8vhVDd19yz4V4w/z/o0Qym6vvKfxy/2MjMmx6b6plPPiVyquh3+gW/uTCm
1aiPpfi7+7ns3VHgKq5VS8A07mWfcEIC7hNceur2gvwn2RbX2d7C5C1xkhKnz/NebMkHIHDr0FQu
uQu8KTdDyAZ8cCptX1sx4WBQZFpO26LLVkNV5YqU4mXTS+YfzMtNzu7JqZW4nEMhgJTf591XbUxi
IcBxoazsT0jjqo4Z/QGZYblK3O1chnZBa/XybIB+mJV5Q/vUZJpxc8KIaBGfbhnNtEzkZ5xKAFR/
8dlxjqSA2yrWbbQ7h3fcawlptVmGDp9K7wOw1khaErexVCrT1ruT7CJDFQAGX95BT4gOokcrlCtR
6VcMC4DYsXODBOKL635DF0uca0NGEOP3LQcHevILQkr3rFcgfsAQ7ayblw7r+9LtC1k55zq4eTNW
6Tz2+Jl1e4JCg1Zpwd5dFfLT6i32qifR8Y1btl4ND8lVRXis67OGgoGAgW/bMN2N+JQ6DCbr1Yag
Kh8IFWHePU+GpsHh/K0/jA1+pQDl1z2A+6vyPYZR9P5R1PV1FXACFbgeb4F6fEftYDDzY7Du9o9U
RdjrsHL3DgAnmqM8MCodjvfC4fpJ0s8b5DNEovZ7t7mKQHKmVnCOJ17yn5wJ4g6GPQQt6VWxkX9X
jKxrNm5UN7rhaV9HAOEvrl0hXRob8JjNSt2cvQpwt6olNH1ncakWJGmHMQfsRTYVB4YGps86DP9T
XKo5hSl9MtegAy2AqUDT6YZzyN6UBiv9fdLGbd0SV8p9YbxJ/NmrZWMStWQI/c5DYXgWUHOHjuDe
AcCUz4IEgbFtMri+ODAJUj27qiargM1v8lDIhUvpXbXioeTfhsKhdkz7op/VYJucYs2Wc5dbSikR
iXo1Xx6G5ZLgR3/AQuw/ZiFXs/H0jWfmsbTLLvmoXlXQTaw8k/0xTD9uETOQnO/0GOaTcDCUiUgU
79wky2CtnIX70t+/xAgkNBu2HHZ6EZwXMvYDqPsN/ar5p1NlzxLRk/KiGsdon2pJmSHGdnPe9zWi
x97kvUhhA3uIQDzmGVnQnKjACyUmZc79uJq7xEisZVSJ+PgGgeX3BTbm8UTc9QY1eBwaP98Y9XiE
liMIU0hMDHl2bCJg/VG7YpuU64yKuehl3y+MnBVNjxwJ5CZxGofivspb0/cO9wqCmLi6wTMGC6U+
mfocqKcOzzpQptmUpeqaWk+xEKCjLj8N5nTdWreFKFLmPsH1+dvnOLec54K0yCuN/Ez+H0hbm6fN
/v2VKS2dNUiLMndr6+XCwuMS8COtTuVRT1qSCLxLtORPR8w7f2UQeh5kQeW/DrCGaiTiZ+GlRTLX
N++2t+wFzs5szfjFGGXA8bccypStBUK/iM+7WSItC51gJ43VQwbKiTd27LFGzfdG2mVe0HKagI3z
0gqwo528VoSdcy63FtHP7UwKZhxeUobYRbZC8oMr1S5JfcZGQLC0dsDTOPb1OUR9QhZn/0TQC6lB
cTEVg3X5FlhDgTPbaxbPzHyH+v4IMswWk5BGCQLsEgKqrEIm/aIHrr33vrubB0Vs0YYIU1Tl6Wy+
5+OjlUtyReZ654NriCc71WWFaPmauBaTC90k8XUnqgXwKJQklqvrQ83W+OM9J2QPNU8opt6NLZsK
TeCmdKgExS+azlz8eYkvrDZTADxs9ru6h1LIESwQ6bxNnbhvZV0aR9OcqZQtoc6sVhgZQcfOk1RU
HMOn0+6O31ji+kUE4M8uWoH59BAk4JSDvDfgo2bdBTwPQWcEeRIr4pF6hWB5ZDAheCgo7RNaAflq
9BUnjmJdIi0OM/hq9YZW1pqSSOAiVmL+ZC2H8e/Y/WU37PvM5AEixBYT0LSK4MbVQi/L2SQxUBXQ
9haLqG37cO/Cxl0FELvAnvFtCKSjwpYmVts7SanSvUnvD8TzAW06LrtpTJ2VbmK4gISCWuEH3EXQ
WsPk+2XS8Oyq82xSPmbr8FE+3+z4BwcVe8UZzG5+jknEcpam8ZjO1Zw1dKNCi7DVVBDKC3R6HAgj
xogF9h5FX9eeyV7QANafKJ8E/2ik4UnSNcjD0jzXS4N/YKHy7Ov0omqTjveaFD6orBJ3OVvOQrH3
IAN+W7XmEryhjV1PlmDbd84gCQdR/BxtjB3J8rcfn6J5r7HyCcz4Xu9U+WF+VLMU4WMTEMgw17W1
oUWbLWT//q+481XI1ta8MSpzAKuZhrscb/wxjjvVZu3CoV0F4xZPELYntFoL6STyUNlYQbGZ/Xic
5eh+mwKriklvd8WonvhgwQUK44Rr+lU3BXMadrsyOlXmr+HgmMWHQYNH7jM5MghRrDnFgqwbDFV8
CwPWaNziazqEaqdGwvjTFie40y3AzUPvaR1FwvCvs0sZeoxnC8zF4gyQS36X6P6gqvNu22xtXgGa
ZB642XAnvRAVVNAZhp/gf+HwldMy+qpFVDijKNjC8qCBCTbSBk1Bs+H37Ss+CIa3PQAeuJJxkoi0
94tNnMg9bLqCU2GrtOKExrlNoJ73P+zsUUwXJHPHlo+Ra1wYZLpswtzolVwoZjb89Hd2VAhS4lGn
APswcm3cf+mPR/zoNg9qiKN/RX18jF8R5HMofnkvNDudH4VfvJU0xiwQ7WKqHiafNgYfoqZ2+9ls
H8o8FRSDv+2HjpoWgCAcxlgitpb32zeX0SJLRC2EQ42KbF9DuJ9lBo1yyqD3JMJPHYt8zjd22q6P
8i9JtkykTgBM7+n5YkFlvQ5RVm2naI1mQMhYtuTan8nTKGPdYkpnL7b7D+PDatYhwuNZIZF8M59/
UDVMuNyNpy83o0zDRnRcTEc4LkzJYdetvhIVWobg5KFYGkyJT1IvcgaviJ0r+FN+8ERIHYGWefQt
rv/iNR+praS6nMpz6uB1XHEen9M/SYUo6SY0jUyYI6pI/pFhBYNm0RJJzZnxpl1qxKWNPxWE9wPo
V8RBrCBl/l0m/Vx4IADSR4Kzdmzd/GRE2A/EfjQyUtqu9gWa+UdPVn8o6GsshYYbGuVe5kilExV0
q/GqBRi8McEbWoWKDg+lUegd7xrKdXGgWznhsti7duUR3Y388oxbfIrdGy7PZ8VxjKE8lVATEu6c
YM0TMmqcIhceYxF9NDAI3gCeJWJR+J30f+jEVQWPrRlukoHQkEwjMQoOsFDwmHVil4MM3E/JbUp0
HwbB5u8vZDhR9bP7Hh3LjZA3lusNPAj/egEwLSyKYgMEX1ca7lKwtXLFmZxYpFI10qVKa1bFeTrC
Ug395MnJZXKgcW4HhVOSPFl+JzK93rBWkDcSs3IIPO3UuLHkvqcJqCgFecPfvAJjcexPSYKSZ0By
N3QgVs5Mn+ci86xWJ9cBlxDYl6UdUm9K2VLzxK0lwlsrqVSYRVXpZCWTJ4Yx5rmgtGv7pUC/gLpL
SkC2XxCElNPbfYMebqbUJ6Zn8wKVP4u0OekPEZLpJuNhdujtZpRmlYrcgm9DDTXV+xLVPoeA69cX
GVvwBMXQKIM+MDTBJbpSoDaFZZiAesxkRj30tSRMNsA2f3X2TngWH/pFOV6t4fzFpFRh2atUY6t2
6M1gCCCb70rgt+Y5RYDGupxH+3L3/eWOJx1UobEixlgF7RdGiR1SSDOkKX2emhWYdC1DNNirZnpi
fcR6M/ak9ejuHdgCyXnvykUu14qvZzhytlIEVDXrGNwyf21JT9eV8xR27ZHg3xKtKdeEkPtx6MxR
MKpNEIDVAYLSqN+gmaeA4wsY5kkB4qbt2uJHZjK8W3z7sVL/mN3I9NsJKnpFYOFtUwjIPGgOvkO+
NEmT+V6PFftwIlrM1hzvkVRCJGMys7sAbHCKS9OWOnJ26ufFhouL8W1vaeuhoXEAOl4SX2F+uMiQ
9yHwyKk8at2L5jFKyZyWYbB7hMmd4/+EGMni2gW7iGn61RQAD6P39hQwHgk2Ef6EnimQagfhIctJ
OuP11Vv0aCNnCaUtWyZllqCymMJv9rnWMLo789EDwoF4BmXdFyWaiiwW3fPniJdwdEjo2f+vb7au
+KSMzOTqDVZ4Bn1zNzXl9OUQ28qkDHuVG6wnvLJHbvctCXaZ17NkGMsMW81T1BzN7QU5H4lspl08
74UF7bA4DprCtNeZYsPlDSclu8I1RpMtU/wbs5o8dNkv/iotHE/0GnnOEDA6Fv2jrFsu8GHXYOIa
NcLu8nIDXjwkRxiVZk2knb2yI0Qm3MjObfyoGVbQ1YAw6Z8ojrWF7WaXlRwGKo+KHuhusBK25gCV
FImkeGpTanBtsAlbxmVhq8AfT2NOGWC1x5Q/4NY7Jv/sWtUTuX4ES6X4tU6MQoUrQvzhrY/gXsai
ajm5ADXcCrGd+3w2CwTOm+B2hZiasjDM7GsNGKiiGK9eZR2KZ/o3ySnxjwpmf6RvuT8MaDb3UNTL
ukoAOPGS0qNKwkugbNz+q0OH0s47TKSWc8y9LJ+38hwo8bcyqhcHgd5EmqaiUvor+1y4e6ujVUYD
9YoE2uyXP1N0KVupiyJ7M7WF3u9Qj/dn5BqPvftKpy8h08ObWKI6nCfucsC5p+YlZN2rtM+rc9Qz
9ze6kNBuWixq5sCsUCZy1E30Drl7oBrwxaWcdmEM3TNCUClOXgmVQKrOgQwLHCvSzGdmEdgytTSH
ki8wEBUi2wJNNRG8wQQJklxxk+omJvzoCZGE64I6K537GjvYH+syDwExzjRUNuG7rRefrKCSxNlc
57jVmnovZ/heI3QbHVF6Rva8R46jZmbYbNcCbyHj2wS6Ur4qLCGbYJ+waJUdo8Ba8lo3SB8Szp2A
RL8MJ0FbKCjMZaNgu2K3aZ2arSpF7jHPQXCp40P/FdLIMt/fWlizbAYpd3vRkKe7EFT3JnYRItMr
6xPd9mBcJQqwbVh6/SLODWl1zUgs71hfwzghxRAMK2BYc/uPHV/tB/j85l7mGWyFgbXGH2sd5ZQj
MoOCE2FJKXzeRM1dEmuyQ+9E/7tLlLzgHsFivLBnZyHm8fj52pZJq5DM6saMni14IYdNtNiQPIna
BGbaNXNLjni6+KAR8Zyf2CBM3ccd0zEJnQZ5lkPVQpfWHOIEEoIU+zXCJjt1CReQudjPlwvcwTGg
qAezNNsmnArFn7E5l9jYFr4hCgFzJ631WWp/ZLxZNCGMGqul3CeeuDt7IynJhjnc+z3Y324Bjjmd
qyAkUjoGRbf8pEZV9MUD6FbaFFGI8Bz2EX4ND3E/M8kh0c0vfDDKUMl1SstdQvUHHTqbXKoSVgq7
1CuIAdVfUmDktguaTdPrfph3RYPjhXzwj8fFk6r0rSHlapS3mV8a27wx+tmRYXvmziAi3x0VY3Iz
AStsuTwzVNpxVasuaMKaABA9yiHEZNKjUjW43pR7tUDeG65IPhAsIOM/Z20FjpzaqQsXbf1oCf5D
GE+WHUYyZbuJ+BUIu20RedRzcCihVUfd4cb8HZTSwTBV5TIUbxW+eRN0rTzKSn3BTIa0IHKuOWLF
xTxaZ1o9CO7Kkp+bKW3VRNf/dQuraoHvNIYUiz9HrkZ+GI8lneVR2BC/VWLn0D0jF8rsweRuKNMP
/FlkX+AvV35BoINNxf00XnBvT951rY33pKmLWk0bMwi3o6CPfR1w1eV3+cds17q7N+tDycliJwUO
Qm2Hkq9QplXNlDgSjwWG/vkC4eWAZtFc3i5Dk5+GaVAChQNF0c72a7uaTDeJ2R5PremIA8OIiTSD
rGQ2tZJX7mSb+EiPbGpzRi+fHB+UKuRR0bcc5UbPWBvT3VppZ9eiXZarWYjoctieh+CIXbiHxav4
EVEK/ssHRslcOEUt0QTb7poipLUpN19uoA9m4k6T3Uv5Uowny/A3/tTdj8aJVY2ZaUi93c2sadhm
y9zyW80n2UFo2KuqgPQ7vFnZphlyEFB6QMWmedjzxSqL5cayLHPdin2sn+hE1b42w/MjWPsafZMC
USTX5Efx+xj//WdoigzsmtcLcrRN8Sc6JoNTuMHY+hLqkSFLCpiioDGbhArAybvIQD5XqACCyJbx
Fw7RGsUKU3u1MVTwJsHBtoaLh61L9hGkyry2pvyHN4+TR3rAoiqdbfw3++nwshOn+fW0NQwEyS8P
M/i93Pe/5ilFlyroAqUbk4s3B73OVSKLRUD7uTvtT6xLXZFpmm8FHszdsWX/DLS+C/9Y5DBrtMCc
kmOaygGf/41GmVAI/fmXF2gAkzen9cnyi5gIq5KwcFfG7kbIW3hVGRZ+WBLQR0IwFPwPtFYPbpUZ
JlCnoIhXaOzMLO9B9+99WSfH7XrL1kv27cTrs40n/3yR7NyVKoIMsQFVgPuS/fchxB3Oxz/6Z9UC
cyFppIpbzYmAuDOMbbACpziEMmMN2n9Q2K4aAHwdxvnBo38UQm71XMr0hISA4nyK7snXpL7grI3E
go1RW7v6nQ5hPqCM4IihOJhav+GIF3YxN/jsCfJalMmQ+3U7ToTIbOuARLjH2FCNcfXPxVgq6hVF
sg3ve3/J5rrNqyUTOubg+fZDFB6sQjs1uEjWJFNr5X5l/HdigsbyG1wyDtnG5Ddir0hOpSEUkamk
SKemG05uKf1S55Bj2ho6a78AnRoAldnVljXOyl/exbo52Y6azWDhH7Rk+Pz3aIT6Zd8cVQ8lGiuF
+vmDB6NkWI12Uh1dm9+w08jiWPIC0qtFjTFhks4/rcp49ei+gpVgkD4/2Ay+tCCrwacwJcAtUCZN
ut1QsgahIkGQ3j8LsTw3ctXfAJ/ZTDUJFOlocrJf/RHs+mxNBrqjRcfsPqG5pAGhZV/DEGBQEEtQ
gNiB+8nTlXe4v7ZJs7atIFa0KZjT6ZnPa2hwLQD68zvs8mnlVtsg/j2C8rtZqGWLCvcpP70yxDc6
HfBKJtNdbrVDfuKaewjpwgAOnanREolyZWW7eN5vJ2u6Nl37UcmZhhXSEBxaG5ELN/Fh1xdapcer
AFeFm9lKAeTawGQPye7rxXo58Aole0ADbnEtrUIP6Fvd2ubpXE3xYzlDgZYzU5zdspAs0sEWuxHc
fGfMciWqA/qq+qtj0bBGVb1wY7jN+NeYJa+GQfOyqikOjAJt8Nqh7BKQa6f1CVjGiOrHjUiR2L/W
gKMeeVdueUwOs+Uw9h+mgb1d6shkFm3XXjRBrqd5oLHPV1O29kAzY0lZC0cPPKLsb7JpRq39s3BR
bF6Ji8dkyMxy/Z+60l96I4iLl8+k8rSJdqxUYG3lh5SGwun5Aa2egElyUyS+Jst+gIDSxpWZb5B3
/OBQZAl9q8Gh6g5MIw+DlK13neqRzCPpojMpPI1tENNb0nCLRjLxTLCtt8fgq1e0b/fPKCVP6FMH
825EgywrhoJwcuItiUxoPntOzzuWHsi6LqP4pwpGMnwFY7gD5KaQ3tDU5+CbWvG/ikelHpRJvkNA
sarPv8XQj2PqfCy3+D2B+YqWz4cfqhWkOHMWeic9rQ0zIY2rlsGbC0dR1Y0FSMA1vsYeIY64P4UV
faUlm8r3y3KemLb8QO9M8G2hfCzMots4N8ZsbQtxy5xIFEMmDmhf+eNnlCwr7Tvnle8bn7L+sY9s
LTpwc9tnSu+EJCdv6sMD2e0uT57VTOo6Z1wQb9tA9iw0RDQNy/yqSV86cRPZ1MjYgjCy6deqEa+1
1OAgZzAW9HiOvMNjem1oNE32OihFVyD71KY15nO+YjrJK5JZeKkrBDDy6OA2fhD2Ek+QwlIVIGpn
vGtaQmmygp3ur9kBcvU40ITW+ZAZ+2PQ3eZr3mV4qVXVFEyhL2oR/DQRDXypeUtz7p2+ZamP29lF
caFOaNqwDPrlY1DDCuLwg/GdLiyUXBKnZND2lwFNNFHJk0n4usUfIMPrVVUDk5cPr9po9kBFYkcG
fKB6LT7Ksume5ZaSuYwZgFBofifVaChZ+kMNnbp/Emk8FBkl2T++2Tzobt0s5/J2MU5/W3OLcXTn
mxk0prqjG1sxQmCGVZu89gbJkNBlCy4TOUZbNi8swB8ewAs38T6gmkq5K8oOMzyqtlMkhieI+Lci
yVJFZPviVWEEwH7oIIwxeyeEK/b5deQxj/+7833th7zpEj2gRZwvaUNgK2rO2uOOgY2/YtEI164A
VgeU11G0U5uc7dHLNACoVQ7JlueD27CbMOshphYuavduss9AjVntis+PHK9UiTqtrt2xP1qaDuKS
Pb/ZBHI668C07Ng3d/B1TpdEk+zWu+NtIaxi1pNaYzdDlZh3YkmWsd+ukGHo/rDDetcaAsmcQB7V
dNMO/bqP+n8si+fJT9DQg04Fp4be97gUW3c17sh618FzvOvSGYIuzBHGtUyFUI92T8NDZOCRiw95
4v4NMlTFn3pu1u8DhHSqdX6InzOXvMyz6+g9pito2BKNU2PGxeAcmEZnNOoHW6TMqQ4R3JZLCbkk
S7+PF2HQZ8MtBl+KZqCLW0aFYP11R4CLXCmWHYDD90mm+EE3g57NFuLpiQXGaBG5remU38C5oYKX
EzWkTV0IReJet/7CwI20BOUIbSk6B17Ur5hyx478YfyjjkAbEpi/0DjRCy9S6RDmgFOxFRF+Jp45
DiZUg0Pebr2l0r0HtHzlhh9RbLeSc9wcL8Egzg7uczaJYPBaCp/7m6UFKHzgdiEl3GKubezH3dy6
tYxG9Jr/kYonNFIbIf/xUvs2FoOa1z4scoj8XhlUskWx3iroR2FjOvy7QLjcwEMBTT97yCEYfmib
vdxcZ5pklu03IAn7o7FY/UheFVcRdiWVXO863rYN0b4xfzyybe8EAU4d4w6CFJ6Hodw/ODnpjDjr
DN/lp3K4zv2BNauEttxhY8k4PVH6A/tGf/b3hsob6ezejJCUnlFxhomJhN9fmbpPuJzLiBnjx/y2
hilUZ0fT4DuS5m6WJFPts5won+/3/02t6nXln0yJecufGxJ8GLK+upKPPtCCCC/ekU+TnskRBa7Q
I8xA0lzdMMGUwzhqu7Dgn79L2N1EdKMPSt0H9fPFCJLKt2/ySRnNhxj3iU3+n7HpDixmxoGRJLNV
VQoOEBGmENTtLY2bQzPU63DFRUchz4Mj0J3hcZb1ABbLPXlFcId3nLyyTTfO24JAgkjPpD2MhMRL
vADhzT/ndu/vmojE1VprbtH+WzdnfsEHv5ZR4vhgYFxNYehKSTS7dsteXBvtTQ8JnEbVbnXmRDNF
HTDDoXpf/snkuH6kEvIZzRrgaYPgwLy5J9TuAV7h4/d2BKjW01I8FfVhHPL3JldHQWumVWbm+tdm
RYUwqqDvEXNtnF2WchvrNTA5eWpHstPX6CNiCyXl6XEXqPLqS8mkCNL9pZ+nd3JTJbbQLTOaCaIN
T/UjCZfLV6B/kYz+FhVIDiD9zBfA7aRFvMW1DJEQUO7tz38QIKx9OjZLhjXiZ1ni2aNo9yIo32r6
P8si4rcsz4LenNLagNI7Q3rFt6kNS3gxX5HEs/ntXnkLZB+IILx59jbDNnT/h7xTuezrXfrkxAmm
WZD7k8u7dvuvlCukN3ieMvieQ7xtIdWjhB+jcJ1PjY8FuhZpvI7KJKyZRtNmbr+QoEP8wZS2/anR
Req0keTlo8SesDD4bx+OGNQE4rr+aTCv/aybsGFXba0YOBdwGxdg1d41KGaclYyQqJXjPnTN+v8C
H0kMIsHomEyTDG2YJqjJonoGEAS8FszCQpnd7Xuru/nyV5I+D1t0LW/+QYf8S8DAK67czTUGuI+k
Qh3Fu4bo1qRkDeG/FAGBnBhJFoJ3RFyhaukbt/eqfAcP4tOK1g/hIG2xmovw/U7/kPsHax9zKZt5
nXibCKa1ruC0/7qs3lxUFCcCjjJO6NYOmsxtQCK/gk9o/4nL8QZdZe/yPzEHxZqlzsr1nniz9G6X
oOTvsU/RpgR7fvlUGk3cF4B3YdVad7ZIiG8JGvNV/Omo9xQaRrrPtp1ee+3kRMl5BpLwOesb5FUI
ZWmPiNhYayK1mB6dxLa434GRzbKY8XQhkrjkxRzWDeSNCVPg1a1po5nxEB+iQMF2TXs1QC71HPEK
BLvdCJikTse4YMfEzhF2FKPJme2q/yNPMGvyKVBkz0WVj4d21Q/obJiAY/j/XA6j8ytI98hkTjZE
8ytIDziKjlaN8z6GZk9X6mWpYJoxBtbvoNSg0eXjVxMlfkLPfzbKO5tDhxhTXNZXOjuVG3iErYI6
mGHM9amrxJjFlH3Ya3Pfpz4L/Lh/VRyHlK0LUL0lWDYuQoHSFhc+YYday2ubzprzYpANyi74fHwE
ehi+kBDk031RoRiLhbJLx+MnpdX8k+WVMP49AI2r4THEIypXrsAZA7OFf7kyqRoc0xHkung0Ejku
EMqbbp029x6g+2+BxByZFKpldKLlNWKkD/N3e9jQqp0TtbfprN1M5gl48wRpD6w9OMEshzw2cDad
FLf/Kzge0FgzjVrK1is+FqgN4TDL69hH35OGQFDrXhA3w6zOjsdTVvZFs1iZSPCi7RDkbZspQTFb
wLnJRy70w/JFyo5vgIcQGLvPLo6qNK4OrcZedd3VlF07nG7PJzRzNR+IrnvJ++e5zjWFF905BcE9
nBBoQJb5+XjzhQG/2gcp5G8n/x9d/7PJ3v9+UcAe+lHZ9ZXpf0syd3zFCvs7+hzSGuPD0mIis8tS
ws5u+q24MjEXqapS+6rSyTOPYYBW5QLDf3iPILiH4wJuuaGijtev5L3niZiOwy1kR5XiydxAsLFE
Vad2SpzAYll8+RiDZx+5apwhAcE3qVBQQcY3eJEzHRib00krMPOlg+dQ/XcL8/qFehPG0OAqvlRk
x2i4Y7ElWXHIvFqli9q1eF1++Titw6xja/hia+IWY4iNLLFd1J8SL8c1D3BUcl7qd+lGk2yfKCwt
3GuFu0w/VDvXEJeY1KrHsIpIeT3+Z9n8d/p8OZKPEIlVBO8UfAh0ZaPaGV7YzvG9S5JB7LxpjClB
CTUMtT4lRJqrBLndWYMrD6PdGbl1CgrWeq4FhxM4qSIWH2Tpo1HMX1yN57YgdKU3AS8yceSeCjR4
p7VZnuJzsnVRdJgVpuWTcYBrenaIGtojhzNKJNR56DDPlcpcpvlsmepgJ88rh9uz45TuiVmZoSYL
bhUp1Fcci3j91U7V1AK+HLqfjd5s5qVP0bmcv7co0D0oE1dvsCk/gqnInRa3tO6iK5PfJbD5MTJK
3W9B0giW23aHVXias/kP0QxEzl8WajXDNP710/D1DzEw9CbmDaRZni2ygQ5b6QqbHXkmX7PmUqHr
ITAScrHsQO/ykmjSUDUv07t+YsDfDdfBlg0D0fOxvzaZOz0XNWRY3qkH1HooGYHF4fKRq+Q69WI5
5AL9uRV+UssCAexoJrBvPZzgjeYmdkxjg0T4iA3DclOs3gaOGv3G56Anjwd229WkSwR1G0utRV18
VjLFhXvQ3a2gcCyHLY9hLJJPbG5RpsFxS6bKNA6kG/PUNbznYly0R61m60WLNhtD7ON9FLgjC9sN
PnRBEm+fxbsaqpJYvjIhGFF7CC9RSdqTVXC9asGS9L9mf5S1pnzgUQNqeVWRbbsCrfZnSNqXtpYd
k0sQO8w/yUrSCf8YUkAmu7QVuSsY9Ww4i6W+M6LuMRPIwZZ2LkQTAyal0ESbEaniUb89JVpN+xoh
EBBk9DGkkpKa6c+tcspiLmHWtv8YhRJZT44jE/593U7mHTRyMrjoBPT8vPcvTkB9jplLAlb7PyZL
bKi8JFwoWwew4vPdb06FLG6Y7BOp+x+cFM2Z8KqwcgK13o+V2JGTnYzXoZ1aVNkRdCE22gI1JZHG
c3L18/QuFWuPqIO1zeEaDoGTuSPybX/TXkHdKhxC1UMBmTi12jTyn1IlkNvnugzrUa08nmSYf5Lk
YEqfanQqs7nvqudVoTOE3l8cnZtoiE26XQsfQ2lwzVsUU8WJvD78uyFr14UVqF99hpqhxCfVzBSZ
ggLJN/+ZmLNrPXJ5euWAtIPWs6TcLY4/TBlv07V2pCFjlAx6rG5CjnG2zGPqUNNSPKds+sg0bzJr
epC5GdueSeeOGWLSr/RQn9qcTe77esKYRmnGHxaOtSYSqBlQCut6jX/JsuHoxt4UwuTqEpzB9ipO
TRqiwX7U3aLHzC8aKCneI5x+AcP++fTtQ766dOPDJv8t8/EAC66axP3lrG+26su672WVa/hjuke6
JceJpcCuA3c+edSsHfnM03mRGRa/KGoMvd+ztYckur4U9+29kSUQmeb1pk8e4zmU7EfBZ1/xyrTz
ry42JEyE5nlKyGfx27Fo5C65lkYYibG+G5gS46iuuelWaJ1KDR+0qHBgCm845q6e2SLiPHw/XPhS
mo1RIwv6rBL2bnX7HVJe1QamvyUTaWOhBtW5nVvsY495sjjZ/oi6uAnh1Io2hZ4ZXEIGV1HbEcyq
sm5EDuUnnVSX7Wcf2lzmzwYLQzIh/gTRTRgE1xIg0FL1EXfGauh/PXnhUPw/NoSX9qbxrNcFQSRY
XbH28fD2GwnuAYUlTBIkQifurDdLxGdaw35mMQklXH+B21wtc3gldHxEXwac2YQ+hrxshZrVR4Oy
o392ISGrDp1mP+iK4twLgwAifu30t32G1OxE3wfd+HMJNYujRBREkF7nTvnqx/d2nzEPx8KDNQYq
6pg62rtuF0ym4w9pNmRIPyjhM8oqmta8uoTxAWXvOPZchvEvVKhNCHHvG2AIGXXOvDbfk++WiUUK
6Ola7L2qI5iqQMQAG9+v3YMNfkHWeg/6nvca5XxzCV9L0Ee1VRPNNPQPAt8dOGuSguK/43nH/BzF
LWk4DAyGaDPXnAgGGVAtDGsx4mmJRQpF9Cws+piRcH+BHKdrJXvK+Oe6RfpZ0vZY8aK6P0TtNZNV
ePq4p70neKZs2d3U/AifLiGqeU7prOftFi+mwYrAglU6Ad+8SaojHIhw9UDzpHlNHCIPOZmrC+3V
HgLTVE66G9x4pwx1sQzmvYAexMoE3ti4GWWHWbXbfBRMNVgbxxCkUD+NtJykLXDiTdwxSA/J56iA
0u0alOCrjn/d8mZlRejNad76KXOxWdJvoejmn4F0M1E5yuW/F76SgtGOc+xYxSnWK7cqOSpkp3o6
LHA+0ZktcX89GJLn3EEYLmVCHqUqDie6z18QzOW3vebyWlKmTEl2k0kLiGAgoTn5tuHDBaCtopvy
pbWvbCtKBtN6uZaxhvE5Sx3zyUS9MPtt3h/J85xFVavj4tMrQC5Dp5ys/vVRtNoRqQrQBy3LLx7O
Kr6TKKlUCC4Qf4pRZudADpf1Y+RiVjaGKzjOQBUiFibhMadp4hyGdijNEj925VnGKQnvaSdTggVF
YfXqwvgycVjq1wbYR61LL/oBjhamU76LsT+hSt0exoMb8DOwIXVXvJLVqDBPl0xkkZ4xiJpyQSY5
fhjnjT2Dfg0lNUGLD7VLuPtR9WpJGToCgJ9ZbH86sG1rB48IGjU/jAfFW+WMQ3wv7NlQMikIBSdq
h9D5kwdPGssNcAz1hr0LKQiV/403eztzCKcZdEz3DUeZ/vjm92D63FKv23L8HDO3h8sXAtOaN5CX
unVgN1UpINSfCgqnokBjQfafm9g6iIWEQT09Ul5OxWXygzJScJ6AZ8d2+cVsrHoo+RIHGzlpCrlG
w7yrOKp/9nIDHWG3g4QGYo5A/udwUKePA7p2HnmTQ+6ZGYGbWeY0eM5yqQNsuKhFm0wUGM6H34Gi
NBkSJFle7ZCIUufjUjzvVyH5j7W7HRBIVSuX/iACeX+b+X3JvllF4N+2bfUAhVXGHqXGH9ScjRcn
aW4x1H+0v29RidF04sFHrFvgC2wIN1Zi+7oz2rBgS6eB5r8N/UoNRwzNmqBdnTKgBbQFuPaseiGI
+h+BFHr+OQSwOghKj7dr+M6gjVD2v1tpfIPAF/viPwPOLZtvHUaHJ/kCqCPwlx0hmxMzEORDKDiH
bB/OlPq/OSaCZWJYWjt9wUJKSxES5ouVhB860gbBSpsXxv1lG/5uIWSHLX6XRaZVfiszBIPj0M0W
pYdNFGL/YdW/d8P/Ku56HqBJXdy8IlnclSR1ng9znyKnvKI5u2lSCg46MNgYgwr8W3Zo683KhbPA
g/Sm+W81rOdtAShqplbI2sDi4+IkVuucwGilUZIuHBw3vq+EfYsc2DpXDOWBJAHVAfa/1ZfjDoq+
1NOftR74bJKHtb/pqt24XrsuqHImPYqHJnSNH/EZCE/K9d+APAqGUw/VF30rn4x5IFIrBo9TsM7l
laN+HB/jibSXP4OGVfkDi47AEl4k0KZyERhPFCJQ1gNm9JuE06x+Gg8SyEqwXi8k6JSwrmWuTb07
mfRIqCZR0cDkGYSEXW2IP5K1cEbNVwWTpMKe4ZIT0n3y78n3G+VPQkT7RrjOuRVHnV8Iw9QzXA2V
W6CrfNVHN3y+qda4DnRQ4HAvLw38ibQNorAOmY+Fmv1lVzW+9jX3oQIChYMI6hJXQzjmn/NxrD2D
s3129FXfrc8W/Hh4jaJ5I0FBNxzCNlTpbHyLJcswzOOq2q68HQs2EC7P821v4HcQrZUbEKb708YV
wFBiK6fRKk34CFCyHNe01Jg+lfjmEsZds6n1xOzbzmC1peRrLR/mUTUDHpZUzwiQZSxr0PJoucQN
tHkEFqUzUKyVC2zPADTmmsnM2GknSW1EcFFKM4YVygnOTPDsUR9b04xJj9d9IMJ+kQtCr8L91t5f
NCfzvrSDtsoCJ4nf1+VrSOCz8z54N4TLk6AhbkKDOhWyWP9QEHjA755YjX1zghqcdzzqG2NUfZLw
FWBwetwoVXODKlAm2+ZvBYni5jVHGRzyh+spb8cOU7qdbVkflGwFRQD4tT/sGyX76P/yTQQyML2i
LjzAasXuRBseLg1raod5Quzm7mfu0Ub8rbATR1g4WQPG5D1NQVsmcOodac5pibbm48ilHfKUESZ1
G4xmVfgQsYZJLabuZIt3i6nc4dh6+WLigMPznUQMh75W7f4MaLNAyi6r4shz0AFha0WZ4lAne6P2
vvy+WtYQe+P3/5rZ7OjrrxXvVfPElXjGkOt5HqCJs350zjPNSAIVmQENPM3TBVG09XOnj7y3tAKK
WM9+d8Xsv1bWfiJEXex38x7mU753aZc3xkUcKAF8krhGZdeWjD6NtpkTe63bMZ3n4JYkCNDXNFLG
JXEPpXnGW4jT/XvaihB4uIp15Hzq8ozBb8eTuyLHMN7qIegwmIzMT7Xz5uQDXRBRk2eNpBWEUYIu
3n7qPU4LkuHAJGf+wsb6y8ziiVThxBQBgA8PNoMx1VP6yfdWRBqursXzPOfdpjlOmsXmGV8+6/TV
U3Ttg9X1HlCMZqJfM/zC1SKnuK0Qm/uN5HOsZ2UPIu83nIBOFgm4ETbvJFZu8mbWm9NpoqLL0I7m
Hu4Jt9PvzN3FhR5dzR+VCjTQUCZ2doIZmCakh/ZJ7NrCiKuUBHZ5PEo3YHLhNrzP+soKO+6vOl4V
kMaAdw5i+08lOP++8koEdjgT9PkW2LaWg+a+bSQbXieAQ7UsuPfnz1dcLCAiODgZHVFuWPkxVyhQ
oRXyTSZTZJ0UZVmY5w+25ObqCmGft2ZwxVG68oVMj/b7Ysh2sJSNYtb+X+NUuJl4aNc3sAcCdkHY
fnoAcRo3miC1099OxWxwb0y7F24Kwy3+DORxBgbqK0YhrujVMCLBn3wuvLp9parjbweskpJQ9HA9
qUSLwvvCWtlN+DDTPO6lEuYTDjfrdi83hbNfTJD1Nf+SO5PpdSCF6dwJqR+4K7qdJqnBdd6S4bp/
jI6yY/cTZRgX8FNTZIJkIunJcnyIS1roEPdB4hHiiV2mkkHqfdhj10epZYTAGi3tSxT/U5fqYsSp
Aw83tOJy3/PMfNyDC4ZbiIiYrbR61MMaODfXBNBeOG/Gkc/852zXNp8OXChxiZY+ExjOqkTRojBZ
djS/NkDFWakZ8eK1Q99prbJtUiWeuNVuUt1LUh+JM1qeLd3lgb9ySlSX4yhpTapH7zngmQB1wTxs
EMLqB/BVgx9Y6ZVwmPsTekMiFLcYk9jrASqcw3PL8cjs82byz2C9FGndVKT1yEe2k200mSofYVxH
fz3yY/svwxpHYZsVZGAy8W7g0dAOllD/hoiiYEaeJZSjVUJms30OaR83OejmcvnhJFyNIeMlkn9g
8bY9l212yy4ReDG6y2gc0IHolobdzzExWX712MIOrnSWjSfR9dX4LrQx9t4CulO/VHqpBR5rVcTD
bp38anhC5Teptvb8kXvZ6lLfnjs2tYSf8MNYeB+tODz8zxgT7bOM6GzhL3ap++zg7hTnsUbW2Wmu
DcFum4JHzOnZIJyVx5f6QbTvk8CHYC8HMrD3y+5Sk2dn106T5cv0yNVq1AFUIocnSYbSrUJSrw4Y
LNziChwnThoia2FjlKQMrv2/EhISmN/fzDEttqeSIvmN1nmTtCmMYCDHo/psUZAvtdXWGTNI4Vc3
GAucLXBuQZbb7bZQldzEjQSk9RAMoa0MtDLfvOPcJlv8tQx4F4a+j/U1AF9GHbOXryn2UQXM+gnh
duyy71gVJ3DsHpdkkTlHz9rEed5HSMr80f7QNG8VGNjTv6JjAc0tAq33oVjPNsdw9CZBjnkbaKFC
g8XiiacVhtWEOHLuZZ0sK3HynLNVBEx4nPZgiGF42awg7YhKHdsnqxb6mCeHSNZspMMLF0iLCPVc
2uHUvdeQoMMRZ1xH/5QIQjC+3BnNFjvcQO3aRjbH6zPdknHrSp4YMFFerXnl/IUTghUi2vFT3r0Z
fpKPQGIgEwK/ph0YejUZxKa87r6mOxAYIFxjMm0kssbabqEhxRlIOFlz3SJH7xE74AI07betVIr7
UigVbupbz4OhcpIT6dxRllOD3dManEn8+C4/kFPWsyOyEUv/+WWhz/ObxkDyGQQ1NU+QixaFQP8c
3/IVw5R9vSolX29TV/GG1OTC4Ug7I0GWCFsla2ruga09Xkc3Olydxa6zZXT9vJG/XTDsD6HjpZ37
PVJsgLXW2Ax/3w2rFcWNuYJYTaW1Rw0JqYzA424y440n2oywvk5JL5CHXsqAYxw1tfXnRpcASH+J
Kn+sjpN8O26/0iZlCNjcWhJSd/wwh4ehnbCaHzJJO1UlJFXkUlvUh8ihXx54FHWYPHWeH2QZTprc
AJmf5ySJy5PYzPRa3m0Y50YrxLBqh2Y2WEEqRtPgKHYj7jwW9LltTH08nSeKm+D3g42Ulx/5eitY
EvWhnINCuB82PYC1HWhbHZMb7V/xI0a7gDFuHszoXNZpEa5nHxm86ay9iGFEKX1te0Ms14lQKpsa
I+WKEeUp44RbLC8I5r8m4d8k7Yils4JFYfcEfbbwRGk5WCzpNRQdxzF6FN0YDS+NyIPUJhfZJUrG
9vpXrlWhAQ/rATY/iSh6/2uVqrp6BFj6lswGZWpWwWl2XmP56Q1WXdo6clzifSvkzt1RtUO8uQei
FBsXuFgUmIcMDjegaZMtZuI+PnNR15v0DE0qQLDOH43OIckOV/R+OSwL1DT6q9G2gwnrXSO0nR1t
zDXvlrXezRo/3dH6EBQdRwPz30IIMjZubhXp4bAfwwy3w1IpXW7muSB8u/21db2GN4UPhtAu8ZAZ
bZFfdIrw58PZoVz6qhoOuw/TpMEfOAkPV2XlcHjYMTrEH4FZ+CKxLdBuo9Yz5eC75CJIuYAQ3hNK
ilHixtA1bryq+iNtqIjevIbpCvSaESEc6vGAayc0gYsWQu6OFYdpk4SSYyon9EdEN3gEDTiy1Vnu
0espnpvf7/TiPTr714IvTQjr/m9Tyu7OCB/PmwAliXtxlckXu46cKElC2/As9VG5kvvyI2aU/cOo
HERlMZvffS3255ALVBrXjLr1wg/aN0QX9xC/YIcZAdE9nCtcSENgtjIQtxZMH3N+Llt0J6JkKCdJ
/fKWIIZPd20LCkuFW9Cj61M4XOrHfIeM9S1WTfbZd/S2bb37k3XlMUn2yUlRn46frJkLLgdvn9XZ
YLgrOvka4abw4lwgJEmpbNSLJs8R2QOvlwzBpB6RatfuqCAWIt2r0OXiwae8C6GigmipH3Tn6/Xf
V9H4UfiVed2joUinKGVqsR6AzvwF3bWefNpWIyHWvWz1labEHMHcckpqeAyHhlLqx+Iif8gh3Z19
4VywLoDXTTcX4W0h6tBnwgdj7K+c72KxWJy95HRs7siEh/vao1It+qxuC6QxjtwO8q+87qVdfQoc
F2X/24V1Af9GdcVdhjNpc7zs2uNXshoENm+muzVh3xj9Y74RzbxlxEl+SgF3oLq3IwC8CCYn0fXS
5X39C6v8hPBuEz1yxqnHLy7kNwXdHTEToug3k9gvGUJYpRE8HM+pcR6SoddzfHp+u0Tg3TLsxjqm
mGVZprjebssmrwx/iYnkY7z1wu5taHZM9MxZmQW4a6irIpJrbK5OBnWibQWFa/xb1ZC9x3jNLyyr
CYw1xZ2x4wKW5SFPsR+mizu+MYVT2+C6reUbIB86y2L0FW5xOjQWIZ2rUoz7ql+EKZ1tU8cUuowc
W9QqTQ0gG21Fu+GvWiASTp/7gbtHagnW5uJK8s28TQjS3O9aNn27LVcczLiYtTTUqUu9uQKFC4Ef
ttPYHroQjQQ4xoJ0tVe/PlBfzNZ+rs3Chze0bfK8HpwTf3sE3lWUb36LcZEqQPUf59X2wCfpZNO9
Xx4nJ87WVvl5f/lYe9/H+C3t/XzRRdwd9a6P9rRHw4e6zzoUU6kH3Ak1+YOmoWas895sqKirjqf4
swKv+uiuF+gBotIlCwzguR+bxD1/4/tWOFG1GD32Ld4f5qA9D4/x6FR8t7H80iMkaO/CMFRkEFrj
J/M5NLoBruXIEzYNhT0rDGv5QlXNIAxNhEMYg3Ov9OmWT0RMaZoN6HHPjfeLzvFjiugXCYtssDum
Fmc7gt9yiF3ktXaxFn0vhONrfnzKt5q2PUEho/fMdFXKjuILHQTVTo4WMj3hP99+VGz7Jto6eEp0
q9wPvJ99/jNR70BS1qNY1lqDXPBjw26woSlaAbJDFQ5zsMjbK367vk8a7nVHhxdIjKhCM2PQ6M30
jWuKA8WZ1uCJiRIN/BsIKyZcK/wBdIsNJakOSOrYG/yDZwxc8ZMx8bPHsOewK4+OA8JKRghoP/WR
JzLTnk+tzYJt67AJvIokLAfNC2bXv3L8uV+gFZu8hBGxOByYnfiYWif5p0gFmvP0T/by5MFJuDdd
kqFI2ZSluMuLFsHot8hf4cJpoDxD2Nrz7Ntu5Of7zubtR5kI249P/cF8znIMQbEN/sfDtqKPObI3
uJJbc47MdsUskP1Ow2stOmMvrfRbDkEcmEOjsFbdxsPnmcNJ5rjWTraOhhrWje+pzXOnTQHLbXaA
sOc8z9n5qYWMfwEq0+7Gow3IRae+7fbTkHrjyi3U7JMfZ6NQX0hHK6PMSK4VmEa1aaF3OJN2Ymmm
83S2HI8ESfhFSPq9KHee/vdxJS7BswG4yrnTqMtT4gChJFBp0rtj9CAQS2hClqEqpXTCFxfIMmxe
iM9l6YZkPYxOq/6PCtLRUadjgbTG90ZG7yAqQB0pnxOlCNgyAHwBCDF6xltmo+XcdvjCZEBWF2zI
MWDiSXxI43H1nwlWCOYy3iawuGBO1HKz3uZhzc9mScNknQPrUlZ6Zz+eFeomHzQ5emK+DNiiTo+9
C09uRnoLseBnWOC1MMHAfdWGTyBcHRNI8y84EKXea0Fw9qTzdNnuIAFkQpdiVq/Ur1hKf4v5VKFY
huqGn6Ob8lpZb04aemH7YWKVsLiHZDjxiQHVUaej6rvmN2DA0pYm6KDtqL/eX4v/adAt7gc4iUrr
mCfOakCoR65LldK/PiZ6Sa0DXEVjbzd+F5k8PPf5jLrZDxzf9KHRWBLRfNtfNz7dRFkigB7Pt3hJ
FAZcmpWKm9RPClu070w9mnQVgTb8NGohnuvUeM6m9w+qdES5b3wYIVLJSVfQkeuqfxXy5VMMt6A3
ln3fTlAqEaNTaF/Fp19elxQbjAsHkJTS/pZI6ileH08vn4Mloa/O2HFU/tpK0uHiNn7Z1IFp0rya
nMtW80xAz8Y5nhfQqbt2+dEeDMvS5Jh2Ys5jH1dEFIjjTnTW3oRRJx+dHEkejmkUBiRUxDYBNJN6
2cKhtbzmYRcT1lrr29FmiCZlYfLVV/Bi3naIPEPvY6sTrq5MkjI22DJdhlYeQyYxDggMFaPiNk8M
X2mDMPTgR0M4YwLz1zNHnh7oBZfDStfx6w2TGTIWv6G9l3U2bJ+zt2fvTCF/s+ylnAZev/LcK4pS
hFg7Y41aWqXyBUqlmprCkU/Msvq8emUBW3AA8zRyHWhPmCB2FshvcSYujSbJmW7L60jviUF7zuhB
6g3YR0iVE9HE9CTfJqaNoG9kCJs75uA42PpQZPhtKPrhVx7rYLWKEx0BzLOSHfDPyNZZEwCEPGJG
i162RG8JPS0RmkgKS7prJRBKTyWa8hk5/lNAm5Tj0LVDR4bjBIKTjhhCZD8zU7nVIfzoA/TKj2bE
7CTwwLYEMsxptYBSgKaxLsUYKRqH7MvmwPOjR/Hg2qSG5KepCA/WdIMU0vYOWL56nXaRSHCRKZGF
zJsT2fb2+YrXIKBpRQJeGtsX6Gi/zS5lm3Fv3OF/JO0/iZnKwMNbf7jr04X8cEqgS2q2j5bIVu07
7jAKwPMlgjVuSidHCLXpW+vPONjqvQhDzMVbsCyDu3SmWIilbT+bYo4JoGxZtoT9BlKsKKjjvUEN
kB9X/MjuLriJU66maiVsZUzN/zVE/TQSIUt14XasWcPzj3MtB0aNPWa0HDkH4IzD5ng/u/KxgjuV
MpmHgpfrkSbvF7vU32BXQ25oJhlyX8+Cs+t1O5NcuuUBmIc4hzazQpuS9b5H9NN/sLh38xaBmLzC
8Tc2iKEho5Lz8AhjpUH6+7foM9AWBVhL+AEB3JoW01D6FYH7Tfj4cqrK1B/K906DK3xZd7KIUEPv
Szck0bQbimCFM0C6BMkfN6CiNYsXl/+27QaGAUqJfXY74kHU6XxINpJw30PwzQ5SD544HP2IfbFE
vIBD/sy4XTmJNAyyG7BwuzN1XY12ReZkXX02V9KzulqoGGt75Jfi2kW7TusHJOSopt6z4/dvs2PS
FwPT3l3phd0B5iLpzcbVvPhOWDuLB/jZFdHZVNpzwiiysnzMaN3OuuVsjcCA3xdSBWPlzhyditaB
iIxsqE1gxT73L5i8MoHcPMbFFTm0MiQFkC3ZJt8A6RlAyUR4rJ740j8+czbxCIcimO1caa9G3DpR
grdzHFBey9lgqj2UmOToHB6ToDKTqc8XkCxLvci4LAtXZ4R8OeMLROqvEnT8rSH7iS3WQGz+WgEg
CEsoRieWivDRAmQ37HtrY96t2Rfa2WijgyJHzDpLQ6/gYNyQ4Wv7llrO4Gu9WeuO6/KN9A5UNbFd
+V4rb70tPUHS4wq+WqIuxV+fpWpp/loHnPUgZkxHAXp0iYps+7WHfjMChLe7l73SAzKKFIXDO5sZ
vOKzX8IC7nqD6YmyLFQnAvbdwEezVKDRBYD0aTGGpLZq5Ac1BT98eXJcwzB8A/ra7DC2A0S6CoFh
mgSomQAv9XBudr2GXsV5tLkrSk8OMyoMpVqFbGlarD6L7qIY1XlEgd8MdsKjvIi6hA+F6c/tXiqC
xV/9C9TPNGF10vui5VxvDGFLI6b+s0kngHY89C5TO1vschN5TItP7dTObXTPWIOmYRoejjO1wr6b
8cunBOk3HQ/oAGJOCUKkbq2Z0Jv7A7swcTs9bw/qutuW28KNfC56erCxZy8Nrx1VOfrjxR2vZFlb
pUGm/i/x28DDzo57JhrSTwe6+9b6oqx0ZjatfQxJp0gVyWfywaOXQda4qiQDMTqxFhXnEGfOyb6/
WewB8mewhAf1SwgHDs87FjDwZU008zZkJyh/7v9rMTY+CFLm1xkj4LwjQjrAM2ifALplucNPDBua
NfPlE1RbTvSkw1yoauBZzu6zVAs6fGRRkrlH/drGjoY0/SK3thUOvHBFbQjfirzEIRH+I+ZQTD0T
5MBrjQOxMoWKS0l90gdXIS87FtYV3R/pUcU4CjupKy4XjJQgnrqJ7Od1i8ELeNrK6ldTEM7jXx/e
lNAblMZatNO13o76GajOIE/3Lb63RRrNxyi0ABEejAA23GUxZk11pQobXcfwWG1MrpcbZ1X/ctPD
kDcPVdSiDWRGpqTyXTFV5BsVQ9n84OWu8feXySQNaI29T7uEm+qUQYzc0MJPnpI9WzMTTQ82rBCi
m59GlSS8PktKNFEqMHJM9MnQeipca6UfkzpozwtCo/sMX0zkGrrntXmBsh3PM4lvXqoOKy2ofSGe
tATEnvbZOSkmE1ykWmaFP1M9KUa3plAzwEBzn1UFC3KtqpxMMjMHKJHs/ACb0EAiXBq91XEa3Y0C
HC0PMZlVkhWk7lR0KHpzweJFtGzJ1KXfAz8t6f1fCWyKsZSXMKB8/dbRyElpmFFxNFEy5Epli3E5
qbG4OMD8czy3DOVSyNtr9WZBTAqeHYUPU/d6r0I2nmHvYhbh0d5ZwKcWb4LsTVPY65hPADo7AyKm
tL9QRZzhSQZi40sGVnQcwOyW7XNkEkA+XsVi6flH+g2p/XUjGA+mcQAHvifyN2juHIjRyJFvq0AB
tVnRHbxQE7mV06PYRBQ3LAz65tCRoGXxTvzvkrHv/UnlAEe9Bc9AseTgkQCTk7+12kfztxIlWZVH
YWZoY6jNg7ZoFx+/CKe1KTRR9FFMmvn25MnZQk+j1O8PYulV8pwXmPGZG22h4cBOCJi/NSchzV/i
hEkPUOcRaAKvuHbaeFS0Z2+9d4ZTWXIp8I7VWftudpwAp5utkEuP5HxS+tVASVpktjtaM7DEDUQc
E6JndeehzUhLyBcrNeFAF6gDOi+EZtKEM56fpCbhJqTPUfsPW+1VEAzUem1SDWZ9HcwPkkmo95uo
GvxbO4JNmSGtU112SR+j1ZgAAD376Z9WQZvDd3O9Tu67ZyDwwXGHvc5i6upijWtoKt9gR0w24QB4
quIqXV+JiVqCjbSBxJcg1lCDSRPhvY8VidMIuH07pyJ0dyZTbXhneJCjpOkAp1CerUoiyNNremem
wUS+NwZRM9buo29x4/yf2Fpnct1TsBvcQFKZK5QZl0PSdcSomuq6TcJtzcssYq2ecF2/fDucyALl
eH3bi5CAYtLJSEb/rWhSGbIrpCOTwCFV/Yq0zBMtk6v+2emRX+I+y1h/MlhB20jpJbnLt14Mvt91
+8JWy2lXROnAxRhqMmFpIGvkQDydpTIOVtu2KFJ2TPe1kpjLfZcCt1s8wsW6GwYzT/gi0DLOdO3x
j1ErioEb431qa5dZh5m5vzbMt49U8OJJRwiLJUMvsJ9bvNY1i1Ikz6jVb7IOinImNnCi5pnJSFuh
LWZbTFyWVGZb1gv8pfspABwhjn3qom2hsJIj8VygPBF1AB3X2OeU6EAEwauFGnViQKtsC/9FDjKd
uHi05k1zBjcYU5bYteHC5peZ4zaKx6dsVqNpyvM/Hr5ZX7xsS2SGsDWXvccxT7LWlEpjDxHpZy1r
1z0NcCDt4ojE42UYknRe9NmqZqVBwjCJ5RPejK/WLbAFGy2gLwwlMLY0cPzQzEvHyppM1xUzd2Iz
zgSXO2ZvVZmML61BUwpkygeU5QTHPheH2+Sh9OyBWhoXtjtiBpOn+FPhuyAlgRF4N0ioX6LLoq3K
xBlvxLQr8812adWK+YJ0kw4lcha5kVKLXz6LDE+Uf8W+CC7B3TOMPqsIoinSV9LZJRyvXsEM0FYI
PXLYXZB13amJom/tvF3zS/TF4EvWdzcghzUsXckmQu3wDRqQRxNBY0WqBDqieMpyQU2c1gtopTvV
rt4Srm9IV76mdkjqyP1cPgbn1ZIXutiFSwi8MyWWg7douNnmdgiKT4nkyEBXkEnZghtElNoKo3i5
0COzqjldg6HifP4ashSYykCR1eZjM5ixRJa9COHCOHTJJk/vebBH3MFRkj5jbKvLvYCRQ6zGXbdv
Z9gKUgj9KS0eiIs7cuHzmdAtredpBwNKx3bGwehZ16jeeXQJYCXq71YpqZycDc+PyNgIAX2KGxIq
N7o6poZcNlJE80lpHnWBMP/vaFsB24nFZC+kdqU7AZ9jxAD6Tidl2yf/2n0S55M5j3T4SH8Scxv2
CzAIdW/6WKvmxUf/28tO8pRM5gbG8jpvVVJSoe1IOjDs4hPLlUV3Coc8+pJ9lodCm7wjHRRYiJJ+
IJfwd8p5hSReRcCN6QcB2P1/IHHiVZZUBwIzq1DIdC9rvL9dn9xwAJBvTUARfK0QLCeTN64YiTVD
TaSwOBZJgzKIZ9jWHYOOf22qNj3cb50UJflIs+YWoKEKWpqI6a/yvXuUuxWsyebYdwFsD/ZYud/d
rwLLaywUrnhQ7cd+aQDUUdrHedZ6dFay72V6YAUv5sOATQMhJ9quo6irQlhlfHRlZ1DnOamXYOPz
O1ohN9CTLR4EQqCwgcXTb72Yhjs9vj++UYEQKQsypEiUl1FjFuQO3O3iIROQhJhvZcrKz14g7160
jKi9aUmfyWjAlk8JhxQMqqSNIW7wtLqOLHclcLBOT4S3Q0+H0dnkcUAqaH+7VvmhP1chhN6D3x97
7U1ety1LjamhOedP7/dUyrrIz0Zpwj2O+juqeWR4mbJ4NNaR1QIMLkbcSVgZxLJNhNPndwyNjTp8
SxSzccDdn4ngKvSjbC+xpFwkwN73E1Zc2Nxb4xaow7gcxw2ZAGHW7nXi2lJiju7b4NM9vfa0KLBQ
ZNObXM6imG0hQHL3yWLhFX9OTmloA75ZCDaMQ1YSSisqdYwbv0gQS62MUBdbTw+BrY0AQPndqkf1
gIngJGHHke/eQwfwRCMvPpN9pGqHrkYqQeca8RvycN1Kbm9fwsF01864RaQnO4pwv5acx4lnMMNQ
RvQsFPHVAL1Nhfsn+jEeiPaAZ9JxsarYkdBwWfNn64Mqyv2V45yUXWGleB4UFqUOUmyT/L14v4Yl
E/X0TffWpSm3m8hAy7wpi0mDlIAQzv9LQOCd50ouneJSjB6Z4jmgobFLm6+qNXIvXvNUybl/wPt7
QmqeupLQVJZR6aLDIdIVGaJCgf2fzyjHMbKm4swqLStp6G+c/Rkn/P2YLXBNs/WUADTl6OGMVCuF
eKMa1zlx5+38pzGuMX1fyRheDGQuLHmQSpVo5yhtvw5SYJfZ4q+p1jcK/iq7jFYqB2H62AL2s2OQ
ER2g+cf36oeMRK1XsSt+nVQzJl99OOksq/St4h11LbXh5SFRHJ/oKMHRDEzcbnqEn0mJlAnRhsDA
QXm7C6LycZlNTIb0l/tHcz/3/e1mO9Hgt4nVnEOcZyylHT5qIH+KYXawVFBwNYOyffqoe5CyuVhr
m4HrO4Kb/HNRuJV5KC1KByX/F/YWozMnw9NWHYJT0NMs1xdvPuu1Mu5wt0g0e8KliY1O7mg8lFQI
yJePkp6tbn5QXkOb3P8GBpgVsMSAvb8aUaijWyL4a7X+mgypgoml/qCST9VRMVfPfIDzqYnUBp/u
ZOychGU20FkgXg1C+PNgnUygtF6Kxu17IfgbOYdTx6lmO8H2K3D0oeh5CxX4sfwFLaekN9ouQqmT
6UToY+4Lx4Y+WrZNg8zE2rtoVqRD2FQtlmDB/OZs2klCc4SU4eD5FTTNlxJnLIEqrcx5czuKryS7
XegDzdvYpMNf+rk3cgEDt5OJKWsFEQOQXWfgn97UYwPPdiTMpnbcMyH2ngWGxTuGSFcbWQMQ799g
HxNx+CFZE+YWLjprCKNGXrJuDZWCKs/1zrsBcLzsc4KEh3U0UG6+9RzGVBMnoKHgCfLn+gwQdxK2
Pgzho297XXdLetjdcFDJy/xXufVEiqOBclKtnwEeGRQk65k8UnRw+fBYa4P8p7yVWstDJiF/N2yh
kEJux9qPISpcNtlz2ubBBOcQPErcliaogb+CjQDQpzgfOms1ybBIgmYypPTMQSKvSxggPQwfk8bv
6UuWaXh1i1alv98uk7t7t1flj6JZepUn0f4QFFH1+OAhpQjxNX6HENpwNmY8TcoHIqTSS0Bl9KXY
HKguEjhJOneHok6QH546UgMbvnoSCOz0x/5hpWCuZqTdl1wZPEvXOxLFySGdeCmJPUGG0WEckdLL
uarx5hTJsAjSOUtp8b0184/3OOJJVr0FKu1HqEQFf+q+eBAXUrDf3VddM2ASm+b3gCiUvoikvBa7
n31qIZjDbtsRWw5VEJB1FI6CcfhGpiWSIODonpacy+STHLw3zm/45e0VQ7m0B3CRfgXF3mPaXxHo
pGsX9X2ylsw5Ku5IofgZjvN+5OGIxhtmP/IEASlPCrQO65c7z+aoV0kAJXTuCVYWFG49UFFO4aLb
u/01x68IgqbjpUyJqeUKoXQEA3e4cQtU/ndLVFle2MZI9aeoZHSqOn3ztrfVtegYqhZj4XVK4FeL
H2pEMFQJLQO5iZftkIyMWqn3mze3R5sImXpkafP/IRoyZ0xQCj16gmFM6jedyFp7vxLErf8kjG84
KzzNBZFwP4BTmkQ0o1jMkbO8PIH/fLkh7yccgK7Hob/Hj0sdv3CuTJ+GkPD8xIrz3kZTU54wEL0P
Byc0/YLadidu/HDiSMtgNtnrqZ82+IoChabZXYM9jH7m+UIe/DTEjBt4lhCwigHMDrFdBEhfdK8/
teqWZkRS4hNqlWeoDVXskXWWuU+Nddhh3OVRmW9xt1pc3hDeoTlbd2xyovTPzcNSgSnkAe2FOB8R
+30+lp23LopT1SelFCYA3/ItkqbUELoxc8LcPUsET/TQWO8AGZCCyIu+UCiTv5LCfCfBa4TLPB7+
Bj0SWxXG4VPac4N6Yuxe/K6ySpz4Kkro0uWpcpky5p9yVObJp9GPAPtUUFsJd5KYCX/HD6HuQ99B
HHiT/y01oB/2azB6WjpCpz3hDwquFU9wYo/GOA1/4ETo0O9awBpQt2Oy+h7bW8Tu9CpQ24E0aXv0
hfwtglz/hwtBsDe7lThRXUskDM2t0VEPnG0TeZss2NGg8SfzcZY7p5weAcDBlBAG+ZXYCJix6TnX
z2tLDoJXALyDRWPZXGCzIbDcWs4oxmencYA1hk3TzZb5+ato0WMXn9ofE0lSwgb8jBNlUp4S7zUJ
xUc+VqqUt/drL3HCqSBWxzro0D70sq9g+GoBKCySywceEJm0LFZ5zxbpnAxD83PG0XcLIM7QLXlv
nggcm8XkEK5bsF8GDwZGgavCIknc2kbR3x9qRdE3sLrJ80ht5DUrpKx6oKYFKffxBdKaakQOaWVw
RI0WluThY8rC2LudLBEkSe/7qZkKRXRfxOdKslXo4BFaLzpcveqXuBQXbKXqX5nKc1tfc13rWdi2
mt7h4XMS49G/gwdXEDYGzSsvRa5GJ4rO4EV/e/dXng33qdr5gnSf6DePPMtod+9gp72cDsqwWqnC
LruP6moDiuI1BjwfkZJl4vbQ3+pFOWcV4PqD1RaVH8R6PZl9LXTw3E4CZMAR9+gxGFQ/XOjydFFi
kwlOEdzNaOgmmMDX2nhTgXPTqsmnOkTqFZcA69ds07yqmy0B+V2MVSelK7zoMThP0tmTy4nXPQMu
KaC7E3I+l+6XPVkQKw4hSkmAu69HanN7p/a6YMDuLgjIAHAetWXPHft45w4/q2npv0VT6qyLuIYW
1WElV+Qpr5resJTns43ExEMqq6Luv8w1j32vCAZ2LcOfraao1c19WmH1kA1+LDpWTLfBQ6FIQ1Sy
VxEHGlHa3bekBYLvXr3Yv3SmnXP3Cs9QPKtP9N0sc3Q6n9xTcqo7RNVHNAf046H1G+73BYJhWLUk
AHECdVb3Z4/fRr+KLEPAlCNN+5HTUwu8XxhZgpa2fBBMiOcKya3dvnXexgttc45IuKyxHNFTY9r5
F/O9Sxtyf4IzE2l23C0WVPmdNWhHVptYwqPwyz/ZY8zL6/56EG7CAQsoaXwzBecR5J/wKPmWGxbN
FTGXruyZVpttM1XFhIh+E+UjuNj0gKcuvAZD0uU0HoAVcuVNM8rTHHyUpVPGtYJI6mrOg07vRguh
0QqewruioyPH8GNw3zorY/fA8QFT5xohYO3rLsjChq3ZNMmCx9aepGFl2NvFMgXeqxIngdEmyjVE
1nwwsp+d28mdNEWf7NjpsvvnlrAGxkU7xC3abdrYrwYqHQj0lmwC7jbMsJ4WX5UCd27sv7fiBhta
CKMaAG1lhbEr+DAMXHslaseU6nXmJvswhL0UjCRSAsmygodXAWVf+8nsoGlhpdi+0ZECqlb8ewIu
3vAkV0QGe9YPWjmZP3wzxSjzlJIDPq50xJA9jZ2neVem30hj3Uy7YkC25xu7yhtVvxhJGxrg7AWo
umV60Mf2elhMBRfd3qWk1+dpI1z5FMMk3xw4aon2hTcFvyW9wbdz8ljr4dvnfdwZ5BXhUtGObUmq
Lt6w0LVFz/E4C07EHdTPUhSzv/7GF0ks8dQdAu9DSk186Mmfy0c5+F3CGkObCqbhmeooUBQdWQ/+
39RbgcGTxg7s5s68WoU8KEapsEeHImtPqeBkMbXfKz4k+6ThiSnM2IGZd/didzVtqX/tocbgBEuV
ZJItKjsrXMPSHmO03H3TeZP5pr5N/KVq723nn7uL0gJWnhFrRga7GQQFpK/Cm3oGJGAx80xWIpG9
8MQOqYkLO64SbUDpfnmLShIu+vUEnK4Yxwsyhu4J9n3E4NfRpv8xQNgurM2kS7uYC88jwbCM9mLE
7v9tDuPIq8JK/j4i9Jhc8SYC6YFTcxMRxZRbeKUiNT39jVJpySQf/+J0/mhsDfBayEwD5w+Qm0MU
2Dp7utTVplGOn2yD+3Udgelk0OLhHJHZtHBc3oexK3RtIWcbuU8w3xly2Qi+iKskB+qfEA4/MUUg
tVoQt9PviVeVd8N58IwgEu49q7wxRlSR8RaRdGsh5bUy7TrfLeYWZyvNgguLw8W6aZuOPE7xD0BR
63EiubRxcXp/bpuu7VXeyK/6jIU5abRZX88S1oQcI8dVB9Y1xYK1+aCbb2B0RRJoNBZ9Ifq27au2
/SbGFbGGsEesGy+gFoJYSHqjOIelRm9eUhtCByp7F1XSiRySemUhcJH4Z2CUP2Imz6jdeekjP2y3
wXoWSHN8oGjSf72CMW/Akc9KUfoanGNuOL+CPOyOOLYCdoHDOY1xQHw+QYsolmiepZlsNr2HNyZ8
EaK4HFIVc0vddle8w6Zq0nK4iu0mDiUsQA/py6M9zXfCGDAFzOTOLlW2NG7/TL6yTboXcUl/G+DF
VQpMccjCB+8p/k7Sw6NsFAdPX5SdlFWWF/Ek15u+b3zTJJa4OvqFr+p1GtZeLmnM2nQ710SCir6a
nIVcXEEY/44OQjDclbkh7qRsKHi0nW1Ih05qGJ6y/uUZjjYxHJbVaquas9SaBJPb6UxjeqKU8nr2
BYF6Ssw3tkGTMoz15iBk7aRSG0Y3aji+GEZHAfxRxNcB+GN3SV+8IWDWmyP8S+6KDYFCZPURQNA0
2XYoOG6qxZTGXNmMi1zKjLKf7tvZKjUG6K+8N0r3LJMf+pPsF81sHOtDbvLSsbLZ9vtrVtHszm+3
/1oxBK7PvrFI6h5QwpM3GOft1S4f74TrCqLz9cc5J9uSHi6K9QEFFM5LD18Du1CtIh0LgarW9LMC
ag9ToPpSJomHf0F2JLqBJUGGs22M4uSh9LHUWE3gQsKgbtcMURZ3w4v+kZUcK1l2BDK5/UAsFlMp
ka/bF18NSeQSRmqEgyUYio77/l9uDP+cpJ60zEF+JDK7SnkLLFCU6tpVrbPH20hAj/qoW7RgnzSG
CyKHslIXauaTh2t3+mz9jUdxAYD2UmCwGMR8KnORED+l44H0ARivopNrxKz+Xq1YzNnWMUCey963
ffKHEkPmseKx0yq8/zpX/SJv+gb/LPDzzaja6uTXVED9qRHjP7wMLxQomGw74DWS9mjJydqwgN6O
M7ox21i4B03XEKg3eTgD970upqHc00RHGHsfFTy0bJwSYl9jjAZLNPZeYtSDjyEaVKtHh5pEvZR2
gZHB0GmIVva0y74U3jdoCwmwp1IW20s0hgaVo4RNC8hlYcd//qDW3cN+e4p6RJUJqiL/n0+EiF3d
WHI6jYEz+gPte1C+gYCAPfD+OF8GAp9vnIMOp9oPBjCC6iUuGbrumW/jLc3ZjLPdnor43hffZjZd
eoQToXsd4uKHqtfQz7vQtp95cSaJDzGt3et5bqN622SVDsvxb/+aDsxqHOqBKPSL7ArKSC2Ahyro
dwg1deoPPlexMaZI2DiMcLd9BATDp1n3KsIzan+jTc+Yn+ESsabSs56X2puxWXyOT1drHPe1EQcU
p05cdjpQ/85ofxrJJkhGrxDqbbO2k3tjbjkdIHzyf81VVZ2g1imkrS9JeDC/+8xuplzJ2PzJzfvI
azUnh9LoVAnzW0pGF5vvd4iCvDuZgeKfTlIbwu5cQV8np+P1RLioVvMKlxYIrRxn4AEepQ5O7TgT
cdTfC+qvtiiSns/7RNJMs6jpYmCGNteqwlMvt0AmoQ42HcxL5QfBvFDnkHOqic1R255g2dm226qf
uedy1AzbihG5rrMEfPO3No2pJcupYMqJhzUMNrV54wuz955CRarZPiwzA6e5tflajbbZ43nSOmd6
BvOiyz5gekRJBVCSG+uqIzbjWU1O+0cNNU6Cvx68vLod6obClpCYKrrCKm4ey4JfibGSBIg4QPBS
WoJH+UGHhziVGhger+j/XljGKXNm1LhvPBxk3f9kgG/zxSx7+9UYcVpE7Ema8YdBXD450aNCbEVn
4sIL5HfPmHEFRJcVHX/2U3rggC7L28DIrtW0LXe79S5oXvNBop8IvrvnA5xj9szZSqiLM7tQfe5v
5ZvWASOUV3hdYug7NjC4tbziTtP6dgse6j/Rq9Vl/Z4wj+/etuRZeNWsSR5csVHhX8X5f6uw/Ru5
pVkDpqItOHF8kxiuhNi7tAiENr3IXxBMBBN0CIDHIN3S6M5o1Oa4PoAgNrMyn1LPUD+A0UuteMxv
dvBFNBpchgz+5rqcTkvcu1DgKZ8ZquhM4lAAjJS6xvyUSGM25ipsGTlKXm8jf9U//H5NjYQC7cwQ
nlVWAl0UMTc0UEA21zJD1TZo2O75Bi6/1E//zUhe7OwgPgEWqZBAtVhSagtqNhgj8rCUm/vjuA5e
40eGJ/tr4BZINeoUzK/KqWCpe2aAkitTJlvFzk3w2jBZDInVjWUzAr5S/w0cJTHImrMU3Vo9X9+A
ByFkJudyAQlxAIvNxbRAzLqN4AAGE3buJleBNj/646l9CmHNuWDtazxXpiylrgoOeV0pQOZBrbXn
iVU3AzcgJ/DUDOpiNgqkt/XiHD2iBceiEdayCSgCJYGdrHrcWCKCZnZMCzaUcJ/iuAtFSI4a/FKy
2UZsDRWjAYqazbSsMXBAZLfnOYvIq6yRtHeCz724KYa9oq7oH0EAJF8LTkddCIRwASJcoq4WIrWc
SoXArZLygGKqWiUzwneMqVamO2uulCTEOFLnvc45BMqnVO5FPpVbY5daYLap4UAdmH6EHF6YP22y
kt5JjLOnBjc1tCXEf1urRIPYpwEni6cdISu1N0E8AFPPDmHd9j+Wg6XAIStdBfuiixjXEPuLRp8a
pLx3Emgp6bwQp6NxyCTSnH6XhwwQk+oq7q9tfd0k7qZqv6O3Trzmwa7bRxfDaho7wGCkGB+OhhBc
C6MN32BPI3hsrcfpGYrGxNmDFRW4MAVWwbFUFoyhQVflW8e7AUtGlpOUzC2ql5V0w+F2PByaKzFE
rdUSR6eWBVBlZZUkAZuSWmSJt2ycDygU97D59r9U61G/+7biAjnMyhOgbsoKVxYjNPNAmgvfkIu7
nne4lLwwJIX0JEukbBWwrMngvaT1hDcCoKVSKh6uoZWFPavJWrM5H3wAUcrx83WnbBEjuRSGNnsa
PQ7lPmCFogi4k7cvjP5R0VjuX0aqSLCU6Y5Enx7CePgynCSkLP+nGw/8nkLNkaFSWEMTJynS944v
1/xtJ8p97XNotGMUKZ90yPPT5ewO1RzZ9kU3gBKrHsShVl4GGXYbvvEc7wGaPKNi607zNN2pJ4Uo
K1huZTgztP+j4MJcpPtSnIE2BahwO4ght2O8pgW/NdLVDDChbVeXn0jmJzzaTgRvLzy0FI7V14YC
sb+YYPei6CCXVHGCBIfeKrMt2jPlBV1Rk1aRzJl7lcAkdhdsAqp2y6NRy3aEm4rGGNeTIhQo4g0Z
XPkBP8k88wO8sh3TJ2cDB04OX/DLO/N92uQYaQwssA3pjuZwY8VFV2AKCUWZ2vQHxqdrTXlXPT7c
45AwBl35g+JmhNR+QwcZUKdgGdn1o3dZorO+zy3asxKsqE7AbjGsjEjXDceUtgdcX/6sXYiRtqOt
y/vX+2IPqS0p3wfYBUj0syEE5ir6XSdjKDjsS/WN4gYaG9253lcLgahP9xWxOmJJQ0jObxFxkCeH
A7eiS/GiSXa2WWHUZ+jCOS0k2ydlYC42dzEPesgtghpi8QYmtsfZb6gPZIcl1iJzzh7LggJR7COc
d3aDjkKox1LFCmTT5sEYVPeJFCKqfcGFGSZf40K271OIXZRbtyMYvUs9jfhp0475eVvKviSF6ZYv
sjRVbMWr70csAF83XBkMG2Jl+e4cFVTN7GMlyjt3NJtYOAaMcgbYBmk9Rs0uBSK3hhNG+NwINlWT
eE2vZ8kPfSmZ7MWVop7VLEM3+PPquP7MWrqUrpnRBsp+XZ8k2EQ0C+P3xt0oQrTKs0kQuPFGhWGC
tv68Lm/VG6om0DoFGPwpqjDx94yfFCnU5DyeRwoZ4w06scXwwf6nYD7SFokiVUSjIfX6+UmyqsNT
Ouk/DD4vsJW2TMJZ8AHnbIjzbbQeoYFLdM2X51B7KaI8TdGfRHJBlsbcB8axRZ7PszhW7SYzHW8R
Ie33jGaXozGFbU4nPxWtPu0cVv3uM1zezp310DrOk0etubDfQlXCFvk56WYnKoWMo7bIrf51giiB
+xVGiDlPOU2EYeYIbIYPtYvU0GQ+SD9UoMvqPqlNmH/G2cfUpw9ED5C3j6bJwwL93fGVI6uFiVpI
gvcLwv0AG3bikI2rsS9s+rmY/hO6T1bTLBIPVi1bMHFSxY8FaKYXOyPt86cKin7vriMkqZvJ03RW
Rmuq/4kICVXPtZWSKbCxeJ4BdJKfke5XrxhgZ9i+tTNI5JVufmm+yNTfx81DY+YHxU+yTwkRTJL+
jsuUP8uKkoHr68BozXrxc8DF6cggjP5pM6CuwOtUi5rLk23mQ+3SG4AISYwjFc7kkWIrVK6AE5+e
xyGyAiIba85xoHynoAMK1a4DZN4moxPIJr0037zvWKg5jjwRC4g4vmkxjhZjss2/zfNlCc5ZPP7+
35/IIIqlOQuIpgqGT0aFCnNEfH4WEb6rD95L7XxWG/ok9mI74RbyVj8fvdjC7yLmPwgsf+xXnZAm
eeHltMYfNRTL5WLYakKUoCBcbSlUs10D7gOKEFc2q4imWg7gYyjtCBZ1k5wszxiVZHaFyx7p7ssH
wn08PrprxPJTZlx3FWK+K0nm+uk6v1H2DNSo+wrFbPuXuAV7KRk/mijq4IiRnEuh9sgpLr+gcBCp
2xyYDTzmXbm4XB0Zrv7f4idhQF0rPxYy6wJubnj7HiXWhg0eiKAMeMl6Ev+zBnC3DNsuC7ThdwLy
CUXtEl355+zC0HtC+r8Kcdv391L+AXmsHumWrC5MF87BKK6CIfckSTpyOyDtl+CYRwJroAqxvVmE
3LsAWLvjQZ0Cn66cmgkCRO55RqMdIrbSV9JA66PTNkb5EvaJ4yuoEm11HUyuzTyFXecfwFFpJpGU
1NmxfoTNvCSzlweCiQx4UyJC0xayz/8AtFbLGfsSLCsyWN+j86w/uOCsse8XoOrY2L8/k7sO9dZx
V5iAzrpv6vdEr3QIAsr5OVyLeRqrWQ7kVFGgdwuD9hyVNhqCeyM/kY9Y2gYCjEeUW1xlBjfkeWHp
py1j7xHcmc+5K0snoZFMSw33L0yTYWOoegsNc2sYQ+PsB/PbtCuiXzWZ0abGxe0bgxr7qUnuViHr
ms3W0lwJZlb3XUo7mO22TVbN9m1RgT5XPDOvfEGM+atsrBxEvds9J2BIo2Qc30VrU6NlcCaC0z8E
VHefr0jnnnzTSYyPgoZcx/vSPJj4ak1xwydofXuyHZYWoJubNcK+G7ejj0oYzT97FwOO17P1UHgz
AfJId5ZNSLKTHmJFPuWuZ1b+AS4dUBA3f7awOha7TI5ns1+Nh/aTIeWWzMr2otwaYgo4bUuB7z5w
Wn7KZuPqOFzJQSWJGlDQLus43uUnHN+/gytHPnULvcFpDj48UUgCDmMw2hIR9cS5o60LrSdFpyFu
MA9R+94cYhJ1iQM44p3uqVuF9SmnBh92k/lndTfvzl+IDSIVrUnT6x7BjkwAN5z51B7ay54FR08m
yttBRv5bkZkoYVnHMRqVkZa+L04n/RBtA3AjU4vivnBrcZRpvX1Bn7jDTrePmIMIqnCniOadHc+w
HgqTVZC1Ed7j7J4OrzB3KLmM+TS+nWRvA0xee86mO30qbFAAaWn45MZggxlCNc+lEtdcg5aA5vpp
Ct++LgYycLBpqDUat8Zxcg7b4p6c/o065pCY4md7ghwSYiQzQ4jbyx1l/lSywaBDdC9hLszesUPZ
eTvVh7QnajWLqgC8HiRXTRRx3PfT8C5xTJa1hygApJ9MBW1vvxpCOZptJBiNQ/6faDFKxgqw0P3X
I19NEzU54bSiG1ToqXwdk8bFPnsm3N1A6/CN0o9Nh0F4C/fV2Fu+ib86vRaZf0DRmEk5307tCZjb
HiglfKO7N5C+6gb2YdAYUgIjSUeGr8Yx1w9zz4r8Eqp6bzA0TZA8Fvui8mFv7w7vFBTkQL/EKoWd
dt9fsjHZgRVpJmyiWXZ2O6pDwrR3VtBGzqTnwW2HTsfL6Mdy8ZxF8+BpeIn4OYcY1jVFtsTpH51m
eEG3gaCsfoZWptnkNZxq1ua9lmjsLF1v06+wTXodQ8T3fNM1drybDdwq3RvUhzklnlrdMHAr6fO7
EI5TQegz8R5IWIjOqbuwgd1ySnDQpD+DFcOBw4Js0ql5H+yWDuV5QMhK892Lc6izNJxuhneb9yGm
OmShHG3nZPqO+xpyOHu/HskcQnDpoxepafUfHLRFVQde+oVB1UVX0qUmFCZ0sdfvSB8usNP2zicQ
r3IQixD8g+v1PF9bJkqCQ7D2Z5I/AHrWsvefxAfIkMay5AngqIiyHtLTqq1zXlrqSy7IG56OCyWS
elAb4NQVL9ozAOnY/94DhqatRdBermoDHOXdMPD13MoVMwR5FtUk/RPlKEamURNP7PpQsBVwnj10
rpxaXgiq71k4LWmDWHPHcr8Siza3RED+rV5OGIRAV2n4DHe2JkZ2ZrYKA00aipCVTElBS5t03cLk
7LoZDOmx2uMOx8ve+5kb9F78Hi78q+zPy4wFAgmErQClXV0fd6ZofNgZfXM8gZ/50UA+Tpcfqr//
l7GHgNkN9kH0XyeAiovopa+2bjXaTSXg+QYVCpxjRRh8EUeeJlPTpDtUpNUttESq+dfiWvVnB8Wk
E9EAznQZ4/iJcOCINk96NUQlVePAkpiKxNj/699qodyP9sobc43lfph2um1sYiwGYVfThqsqwhk0
jKAWLKCGJeF1ixjjwkxcskynOh8JLLXVzDP0z8qG3qaXi6O5LZeWancnv261ASJO3OPPP9vTGNrv
eJ1RoAw+1k7RMfXHrlsakTInszizdvEmtGaHD4PaOhhmAjfbqIGKCKKPOkFgoWHWCO3GW4XJXmcq
XAQcKHV76fdm2muDh/2421ISnRf7kTZ+y2EwoNiTqgNdoYDWbjp9U3ZNGb2Uh4V1ozMk9ZYg/Ak2
lUP03DnWICDnYkJbPnBccHd/u3LLjwupJkBUD+vVaEpJrXeR3u+aels5DNFbrkae2FhHFBOMXYN1
NYc7kZkmS6AQfK23BSbQ/iBpbKcSMtFb5wX3Yo2bcn4/dwRWADChDv0x2rC3vx02vmnp3WjwupAr
5LpewMlcvc8RYzF9ls8lOuX8AsvLMJzLdOKGXlrigGmmISv5cw2XOAs0lC8xixfEQ4jsJkFfNfRI
IfCy1g76kKCuVaWXWPfvDSrG3Wzn19dBU4BauK4dNCovYfnBai2eqshVdXJfkTwqBBYuFX26/ipv
NhVcl2k8YCwwaIdVzWb7IYNGxERru+kvpgHFK+Zzz/ojbM6JGEPGc7HCZunaPQxMkN5l7eoDQg7v
M4xyorLzPUrEsUiwHYn3jET2WWW047+7kSBixvtnSgqQwaAAN2+KhnFcvAQ/vX16fYFVIVsyg1pX
+4o9FuKA4Sq8JbJw2R56ixgexNZDs2IHOjcIyr7r6DegyuPIqj1Tvc2WHO1NlIyo+0QWDyLr0T25
Hh+D7DENY0fX3rpCW86szhskX1vpCr+Lvq3R+mYty8jKnLCvppQl3HqBgo88YaWh4DAxUxfurfxl
wnv2b+qCCgVSxMfwPGQnOwNdrv/dSngYMNxN2H3PtYjRAR2QTmh9UfP7KXE1aQlmDKjpfATWZQr4
uwdLPQH+MoPbAwalE9K/YgyfEYnENS595IJXId8emslcMXW7ik3jsjo66eukpN43EvWVrsApeImi
prluzCvIU+GrB5L4EOCNE66TAUjtGHD4zDYvmtSrFM50J1H3F7WfgQi0nWqzKqUKBS/8IVBMMeUx
cerqPUvK4KGfY4iy1XeeXcEZlGfndKoqox4kxYbkwMm6s8MurIsBtG4Vh29wWoJbCraVPHSKdeCy
Mv1QkbgDpJYdCBY3MqndmmU93edX7QfFRZJ5dbrGK9LnIxjLYMk2HQh6wWiB28vGz8HOIrjObH1i
TUA1MsQog4vQhV2lp950ZEaTU2OmUpYuzm1Wle5cXx8S9xOYLxZRw7Y9rFlnRIO/ozOfFV7LwlFv
Jc58XDcQ17MBwFaJ8E8cmETKHymx5u3gmuN3afxSaeQqoL7+Mzr1VJ2po5XKU/D6CfWcEje78Lw2
iHiN7Hpl5sMqTT+SHXBwa1X+VJpF6pmkY6VaV8LpFngWZZLWNledZZkond7Ip/izWhokM8jCqb+H
x8z5fJN5NAKQtcEU8VxA+i3DLj+1B+w1XOTFkh8CcsFvJKW3ZaCTzsF8Vv52m++x1lRjpd6lNBnK
AGxCVEVgb+LTxHFaJwFmrpX+OuzF4Cil2q0/LchhY35t14NUMIzqE528bc9NIt7ju7Nv59NLriQO
eUgJHQ38gfVKkve/P2fOOF6jdvLyfItz6dDgufgeFHJDERi59FKnujn/w0XEchMeN1fVdGQ4PpbO
qdS9IkqaSZQNOyagfWBIoVAVL6k+u9OPWIdT8rmDoOtdl74DgM7aWDpyMJNbQUp4QgClgUE1GZva
HKQN1XXYTeEJB73dWm1BN907Oxt5ttNe2p54WfVEZ6JRGLTR5BONhRUzVMVl+90c7dFvaS+qjV4i
W7JmAGa6Worh5kygQ8chrXaQYIupv75JWwTMWEdT8l6BOJemwVRs+mGXnGiFYFDbhpmIb3TAz9Py
9GWHvwXNJMUJypWSo8sH0qob9EY87ywRnH7vxZkMT8tBiS/A5Rd6Uq2x0zgp/trU+XsR2U374v+I
np31ffpA+mvWSp9TNsCTkNef+rgWZ+o4e85Xs8V0t3lm7GJRTxpLqrwSu6QipZkRHIYbrcqHgRCz
ZbAaWJPkXVnCWYhj+wTz6YZ4ihUkeAzdVPE3D6Wzm8EzLVqrB1XMS4JCBfpftOhA7q86iBWjmP0Y
uj8JEbWrVaN/uxna4KetfDlAF219qpsb3nDCW08WEnXb93UfOXKfBIAHATPnSVVW3r54Wr0aqLqK
xWm/ngu8oVYnFCBZsvDJF6EbakIYSE9usDjW6NA6ciayDXSyOjoPaJdF9CwFuOFYQuoiPAHgkkue
6d4zoc8RqWoL/3QOxPDczYqGfQYNH6K8UujPpykLSAbn23wWTWPFz34x6rcKHO4A1qvZvf7LZcG6
3DmYq4I9LKvJUvoy700SpSAKHo2VcfD2kv4UtZSCO6UQXDuMTfRfXIN/NfD9OUJrTBXuR/0DLcX8
M1bgTK4ozsYFQAoGhyi18ocKUaCgWKYQUNRJBsy6hYxCAn2raffo8gXh22iiK7licFfOLiz/fgvh
9t1tZPsycSx9RHUDeLqAvLlOp2HKi87IGCDAM2UTEcPpgNIkwhW7r2wqDKSNtlKVsAkt8B461XHO
TtoTAvqdC3lIWTK05oC9hIRa48hJfry4pMItLn+e24wanL9FNUOetJFNA/LBy57VbCJZpLjSnLiJ
yUrfYGShLH2OaPj04OW2+PjiIqe+6g36Iw7Q+D+2/9i9jBe/8OhHBD4C3CPs4sDjf3Ebjkf6QdGI
5eUjEW7PPpre7tX1mK5/7aTOL/MVxmsZCFKtDjM8hMqGSuc53RrrnFdcFY5kJMeuHuo0ma62Xijh
8E7HPIzTUcLcJbN7qrlPrqyCqnM2ftC2yuHKYYcERoA1NLeL0ErbpzX9yVXsrUCA5+RvZVKNmdq/
g6XuVkaSNlOWmihPU/ho85BHppJrdGwJyHDlSWfFCW9BqlBtrNyvDT02X7+ZIAmJF991zykznO/H
p3dbM6qRP3kaYZs1QmsB5nP0zFHF39npV/L0jSHlQMBQWH6CQBSBw/iT9kg70G0+eILVdE/J7TsU
q4bGORX9ehWdK5SomQcMk0VMPW2c3pqnDYpp5eT37uNRL5u6bV2ehK0UJI6l20tQuzuR0jUnTLSh
p2xucxh+gf/AIih61L3U5i3h63qSYUc6gwMs/HolQLeIb++vrI+ql+ytDaTLfqqwHMeWxOLrvwrt
584bV2ZPIXEmoVLmKgfQcHkt9+juliq426UGH1Op1dTMmmTPpntQI5M8adYr74r3AR8JnXkSZDi4
E9UQoxd25EiIieS2RJDUIczxZ4KCqKmtLVwHn8y7/uSFfPrKvwPbmW57mbsvRjLDxkQ8C3Xoprve
svLOgjAWLCg++lvsBwCcDe0gObip4j6G0mgMbGtrNSNhhYLzLw0VgUSDjKWQfbajtyIkche+Di9v
RZpf49MTWYIVnCyWgSrdhas7g/RbmnYT/cP/vfuSqyI4WU2Gn/X2p4VoI9OZHCRRMT4JLtjO4g+x
BElO4wgn+tDS1McjTgF76YHw8gpHuaDhPjrGqZZkhFm8w60e6plLknj2etX/wcU0GBQG+j35y3qA
LGTf8D8AS8gM/m8Pst9tZxhJPEKPMU4aVLlWxuEgTAd+pLR/p5+xwryopmmsz7RpaNXPNmcz3RSq
Cr0FoQ36dhuTdDRVv/GQvlR5gcJzGNyPFvimZrv68cmLYqKHXWQwVVZNfaJlo5rtB5OKgNeF64R+
pFWLInBzJPLQ+yB7HdM9N6NmgrYxVx6n2ZiVC4Vyg/QxODh2yMszzBmec/kFD0qelGg0jegAFagd
psr2mCcHfer+Xae2dX0ExC8KEBThYuCsWicf/Ome4ny9f0DOGetEhu+Z6Kj9zy6TyUnbi4GSIrYq
Rxk0r0MaYUaFG7bhGUn4ksDAQnC9K6mn4AnnEOlrx6FOyT03YYvb3Yk24kSocntThBn7qn5i36mZ
NFVfwAaHqiF+1pmRUetGwgtw5YkBrdtT3bf7hQXu9bHj09w7EC7MW/6bX7hUnCwRpXmF0Le34BjA
TvzBGFsYclz9ct+1nGb1EXrrhjZGmxXQpu2aPMQB+BPFeta1sXPcf990WUX13PYc8ua/qHAqTCbH
sAWgAj7JVdXSes0yhnYUJYlS0bmiIgbNcRVICxWdiuJO+/y71Zahff2sXwMlqQASc8NX85kNJ1RP
VtLq7/RG4eqkVsGd3AxDQ85w8bG/VGgA0LyL9Ypt2TXnVu+vwkelGxnOdWKLqRGn0jbLnUiMArkN
b8WbAjNxfZkWBLMfCp/KkvQbUchGF3Ogb2/LFbdDsGYWpJ3UCBZX2YuLTTJLlLUYUU3vaHaSJJ4Q
3xdyYEWlW1WXLUYU2924TLo58OXG9DkhR6uDSk+RTxP7mKrYGv9Y/v8jBSkieAxwcN5F0Z79MEdv
328Uvh6recAIwmxiJgDakHkFoHjrEHmV39QPlFq+z2ikoQldG5ZgrBj2rKPBTVeDYrK6RsVgom5c
Gfy1ZNEVT+sZwH5QIqOB61nYyhGYuj/Q+N9EiKTvMwSOt4Rape7k8jgU4LLCfUjeyqmlj4c+Yvkr
Y4LFs50C54Pgcax9ZlIJj4fv5/Moxc1nhVx03zMMdxmqmyrGfGLZKgvSes0pMB5qtpplGAx7bbsI
LB2zkB7KsSDYZ6QgV5VfxwhEp2O0fVYmE0YGhcePZFhUKtXavRRkUXxRrfIL81HvEWrStzTHhAPm
RlMRh1ACANAVNoFSmc4Z++1IZOg7MR9qhHNqAOSXJm6e34mk11U3rZcVvnkfJjDbtzCv4dhxPV3y
pq1kB7y6rkqg7kbWpiTKZq+V1oQYBRKwp7RLJaa3R5agtn3sRAtqwcpOdRQIlvJlnhnGWiAfSaNY
ThOKEqQX8Vg+/hvcF/DgL7k90y77dWwEYLjdujJjEo2VIe3p1qmE0PZGehmc5bCI7vIBKHKZuKvq
/+tBHy9DNoVIb6MmC7kXs5B3OQMBnYKAqR/UXlEHlD4eQpkKTyirlXmhg5uRIFQ4xurPP0p/qMXq
dFrGQ0R/vLSbP6/fmj0nkq22Zh82HNdjKIbLD3ZkvMkHGSDLYP8FMgm/MNYLlpz2A0Fy/sALwc6h
fklKtuXn/lSrinS3ZG0tMTMIV5i6wGXmRQ2rtXZ90leUCCit+7Ill2FDdhbPyMzPRLTmuGLwu5e0
XvByh94ecF/Orrs/CF41wXAIT1eCneAfEY4rnKschx4MfcS5ZkRfhrsr66zRMBxbwro7CnEs+l7F
hloDceCtO41zUHE9reYkCeUqL7uDp3sedZFEYaGtd1gsRrRD4wnxhyZTLsFoR68+ghhGZxVOq7dh
RfuBDY2I3Zk9AW3J9zxM4CQ8J8wUBjMg5cUTAI1eTIfrRwTtliQwgk9Jh0c87kW0Kszpbo6RQXFQ
6hoGDUEZtpjjyquS1oViNyKp/QgX5bIqCYhyhdGGlABZ2kFSXhKZAlWzpN67H7xE4vIZW4GaWMFv
lhwBnXlvBeHi+pTcQEZuJcCoXEjTq4aQSHyj53+aEH/haJZfRDlatVII7DHP8cbycejyZ8UQcJoD
G540U4y4U0urJST0cqAuYbZYg5x1k/BcPGa/ce5sdloqQVeVBo5gn8YjvUiepAcoAd5dqOgDOGCQ
+7ZoITY0/o7RVAZX3NtJf20At8/G50EJQL4oSRi12ntU6WRGFSMgLftYFWe/N8IW9G8J9WFMiFSa
v925U6vFdh5TbyRi+zJ4ugUD74hVaOdnw/bXZNC2Cxs4JbjrcdXurbrygj13rrnxxeCfPJF1/oyC
mJQ+DaP0jbqQy8hkvYCdI68Gd9bHBpdmFSRNIyXxfujyIJ4+TLKYlkgySNhgqUqdG3173qB5mAB8
BKF1I9AlYIwG/IqylrKy9LwKjph9O/ds1YhoHcBjCiOHk9I40fMP/xBXHwJQbGsin1uxC6eVApiO
45/NqBRuq066VDBi2NTTzN7YOcvKiwV9XYU4QbEk+TbKf1LQsQJm9SMsN9RJ3coetzVMlsLbXM0J
Hg+UF5g06YUnY6s7lFrC7kYAB1bRAmB63Hy+te7j4N3v/mA94h3pVLCuKoZAuOqkU32T2lgFRFy7
xiowFkFlzQbZbW+1m8UBui5vFV2NOea9Lnh7B/onLv2wqFpxa6sqPvPvoEXpIVbZ29BXFBWaKDib
nTW0ozga1Q2usjavlUdZpWKI/W1riPd/IuSOA8ATAoq6Bf3kpEZrTVS5+6VO92dmxHRzHx2NwW9l
Kwi+mmNi03LZurD4j2ObMufTfkCn/dm0XisUg0IiPvBEPqe3QU5MTnREeLAlZ1B/2SpruRnukCaQ
BixGoDDtbomZpwRpT3Tyv2nv1mskwZ04ZStjhmg5O87WCWyRYiA/MtgSPFXFN+MMgRlOz3D0WfzJ
0iLi/BEWgJJi9W6Xkh9dgFMzewEetHyEycSQtjHwesPO6h9sg4edOO9KlsJSKtujh80w1i49Kd0J
IaagEQOpUismk6u8AcPkj7/TZXO6zmCAmtgufzuUOTzUFRJbBBjUGu8HnhziCJtRDeNJPJehrzAP
C0k13i+iSbZ85Z1Bh355ivjWn2Jdt+yIAsjVBv2UeGRnTKi0zc2MEVREO7XfXaLy0AZTU5lhejcF
2ZehXlecHfqIgBEIW3ihtMd9A0TNABOu7td/zNv11nUDKQ9/Pzd7hpgOIM0RBVqr1yrSiNkvsMFn
inq1YMcgaIBOJuseYk0lkr1+pFljKaw0mtcqITsu/0YekLsnbmZV7Lg82NpAL2TJdSuBm/ZHkzj9
JBmjLz2KD3QKTb3MvQl1yDsH1eltxQYWqlsC272y0ZF57erg/9Bbb/uvL8dUbYVA/UMsOSM9B6Am
plSR6HXA95GUfPOW0naRrmfegGt03SAZZy9Vrz5JEfNqLiuZkvyAq6NU7hRLOKWHEt2NNCRfOFcY
yGxaDd8V8kG0CglKIWutpT7wdqVV2lPOXnq+Fr39hCuJrpqHdipxyD4ug2sKS3dH/I9kmEtEPbQA
BHRF6SEEXfkSQKspQfiX718Y+RB5qD/weOa+6wfhCsdMt0SMTbMxeFeFZpHdHKEKjLv2qhai7qQQ
XOu1xWUYBtkn8+ZViekjv6KSHcUtY4sMxM/0nOQI6eWhwo7kEL2WhBmHchcL9GWNqK1pW1Rhy1sQ
bd2NOBiD/d+PWwXma2oo/H8gY28dB/EcdVu7B7cxnPIRnzM+y5/Z6dlBira0ejoYFWV59xP4NcLk
ucWr2fcmQOrBD2IiXHW/ou8sTIjs0P3noaIasl8DT+uP61GKMdndM6pLtSxnhzVprG4qfxTOguXQ
zFHnefQUGzOi2QxprSesDmpkIF5zL02oU9dkC5G/DP0rxlYjlz6RjhfWl2pevoNtna/ApWpcmsc6
sPsSgRTxXV4ZJ4myNK6w6DBzXR9XUjgQWyAQhiqct+CK60nT0/LqJnS5Zfowi1FBuE65RN2gbjpV
gBXY0yYd3mAZ84rdM2LGt9MNLW6GVHoACK5LJB1hpiia8Cb9vKhMfXGBHNgYeMrm4O0af1Exm4r2
aGeo+0LQnASsa9q+xaJFh81I/ZBbIQir3EldhrQ5spvOI5xcAQAJEHm7eARuy9g24tvaJ/Ks7wux
7+/ABXK0BshUNImXX5Een6jpQHDcKJwI0FZ1dwnmArIHr7Xn/p0jo9qQ7KTgAabHvl+7puxQqgFu
zJtCVTVoM3+IwkC2Ghw0wSnbFY8157HBRi4kU3L61s2ju1bc9SEMMC6cWK6NpsRTaL1QO5QItBDR
5qlwo6KtLt6v5z61rOYmkUu9c0QoAiHNzvooc+cHnfgwKlxiJxodV8blur0rmDJhS+gt/ggPzAhq
cS1l/07rGuS6BZ1wbG2yHIUbgdDRRc7QNNRk9FPA/9UUkJrjAJ60118hzNMs3gWsq5LF3HR1ij1j
4HX3z11RR0mW7IbIF7T3BGSbMHghcs/YojDcVfWJU9EIPWGP4V/hZEx8/6T815PyjjFKpV/DStzb
sABcODa+A9HneAwme6i9X7hZhCn/+OUAn6Wdi1k0ewdw84MufAVIDRryF41Z66plKfaM3wYCfMPn
eEhdiOyzU8YUDuJTBi9HiJQ35K1bjE21crzfSEK5RGJ5q1jjxQgDfXpfyzgxg0AXhmcodUJptCFE
Lti21AucP0tB+y5zvLTSxHvQvZxm6IH24jM5SxAT/UKYS+mlW6pDqMY+3eTNMLlG8nfkSarTou/e
1vBCRXF0WVfv0WnYr8oNSHYPqzRMkT/hVdybJOvsb5n+zl2w4MbdbHLVvf9opxAcOUYwlSkYmQSM
r4qGCr97pOzwY9APJTsS73XWR/ftda5Qy7YGKB2dDcOVMCgSSrJqn0tLd+jP0JLfFlJkvKuo0Yis
ES/lvLEDE82bVLkFZ8bB/evUacSWgZlRBUhzUhn4aZTjwzX36tOaRT+8HJjI8kxqdnKasmnoW2uW
FVqKXLRlIHMMlJg1lL/CSGwR/OHrIdk/7V64XWqK78h8DYBmchTHbGrR4xwNyQ/zy4EWBnA1HwYf
0ePK27cxlanC5pTAXvDcQ3tXwdyd2i4AQFM5rsTSrDB7Ht88hbmnf+P+hPzh88tMr3xnRG3uN5Vk
/O5/9yDrtLnkgda2qT9FGM96c6maSZSBEYUvhwF1hMdimzg7jJqDL4J3vbqlDAnpOhF2fngbNxQI
Q0m2lNgpVWj+2z07pxMIe8HaUwIwB2pQGeJKOC8ZTclUX7gufuQdd6WBN+XWMFwRbC45S9NxrAfS
iAo7X4kE99NBuPd2+8PojCs6HjwHCC12eNQun4urByrhLPYqnXsRIQ1WhBCyK+si3YR69R8rPcJh
TaNSSdCXnUO11bpbVTG/Bpjitmo/hURCJ/miUYLaAWhh7O8JsXGSaboUlFUaebsKWMsMeMLDnJ/E
rssNnknILxU88Lz6yyanhzIP2h5dkGI/z9WUmF/kZh+YNBvM1NU7LHqslwv0lggjT3Kr40G87Pv/
xLM/yAAyqF9aFlXwXkkORNhLTHqaZZzaJsaPfCyVrXl5FJkjoprPr5iCIcc8yM+lu/3/82MMG7VH
gGLos6l4aC48qKmMGRenSACTBqe456St2z2bnDHwC5mfj7AAurttlX3Hbgvw1XpG41Ti7WCEaWkh
GAhuSwP1F/yI4d8H0eqpe84Dt70XkBJZ7h8WHFGKJbR5v4p0+AvzpzZezKqYcdwx6t38VKQWJSxp
fLVyhyHrR2YloEyjBPjjavRf7ezc067nXvynfCUFfRwRW1OcZhWCmgizknknl1fLYrLhjNz4q15W
0+RqzxyMDe47TONuknlPmYeq9pfdW/AJfu4wAaYjHmuPROPXtbR+Tjv4L4KAxhs1kHAQqbFHklCZ
E6S1mRyAwg6/q46Nz7opwJ2lCAfv3oYTWdkk2lPsBzJLAZU0RAAKVzlDUKj2SO56g9dmiS+GWvA9
XOQ3zx6KygK0bMY8Wd2UQK5D0nnKrZOxLZa4c0Xvl7RMQvoEZU1KYZZzG92AU6lXBtc3rtbQGAfQ
0vzT+svSuwqVBv+LW4UTeCF5GH0ku67spSHEKSv7lB8iJ2oyuZIW5Q4D2iP/wsHw4ODldNd+q048
M1j5uj3THOIT/0rvPSngYipoqU560Jf45tvLUJ8jaufTzQnCgsJXHE2fcx3nRrt9B+jBxTLadHYH
UQCQ9aqhOJMhUpY31dEW+n0qo2g6sJ9uTmXcrrUezSs7JnHcqco4xliK2l1KwKMtv5Y1D9GNpMk/
Vwkl8/i8gXbmh6StWTNkiGkpTvzsNeuCtc/63jZhmi0HEiMLtn9U9+Y+4wrgHAmU7Am71NXcFW1U
/r+GS26wLnsfmwAEr5YDfXbqtiEWWfVnnVPCUQwWw6IhxOmvdX7ARtXQk0paFaTEG2QcXSYwWVFo
dz67DaIrmEJSzegNgBerBDCPXVElVUVe/Ft4kGsrrMU2GHCe94xpu/lidyWoVlrnAcKBD9JFm3X1
BJgd5Ze0aL7anU3DfJ+o5lpbnlvv613R8AX3LjqO0/s+oOtslZur3RtyCfuo/iDFHilWMglmAXsS
QOEZ/J6c3oITVZYTA7DhyXfgIFeiua663SgjMWBWcepPCZBShyl6iq/swvjB/tZH1qg+IvmdtPnJ
qB+Ek9D01gf0ZYmfwbbSqnWioF7ldXngRvooKQkWAoJ5qSD6N6M5PDj+BDadEdRADH25p6KZBj+R
+g8ShxNj3FTuor0Y8EYatACsmI+TzMiOe8cAr9Y+fLhNRP9jMVAc001AqQZGRbwxOOfQ4Zj5vFzq
DvfgBXi0VxCaK66JjuPP/ZW6OeI0e+mct1FK+ySYCMBO1PdElqdGzigRrzc1e8/tN1x3zhOEov2f
LR/5YyNhFeumnn1hgkjKSZzPRnWcoCn1WgJuxLVfelmZputjXTqcpz4mV0rLayRX82f8pTWWRxmw
96UWze+ZydWJXV0onVQRBr3axxlohqCQvjsRsgjchu0d5zs5WIjnfz2lgzhzNAzujmhj/VOZ5Gg5
bQ8ysCrQHonOWqwYpB1kbxodhP/IJUciTwcjNzw/qz687+/k162waR7D+JXUUVCZ2DUHMM4fylBx
jmPqFnsVK1U91XiG3ItMGMdVeYbhod6RY4kIZppxwISICAdVrBXJLlBoJRumkVqmCNCaCxAWwJgU
z0KVQwGTsTjqEbsVNdcl7+dEe0zRGA17ff7fbB6nx1ZVFX03642GvH67I07qkRWd2bAMdlnpAchX
YtCXTqY2VILer9dzGeYu3AaSWw7m8RMav39/2IednGJIy2B8bZZE4TyHMVzoty9SDMniTnls940s
u6rxvuvtQ3fybm045PzgfsRdrsmWcI4Xquy87MWQb67u+M75S4yT5pIZIqfPPXKqwcmjZAwrCpNp
h1IYBprlC99ZB0e6MuvqR6ng36U3NOy0NyBlvsoup1j2m2eYdubctIkuIa5xpVLCghcUxQeG/Muq
BC2d7NXyaxC7PyRsjROqVgr/E/c1A6FsJ/Bo0QcUuqEIBIDUQ9eyxclXCv+Y86Apu4jQ7Q2cGirP
mRC/UofJc/+UTp6jU/qope6KIjiBRJ5rQjLaSMkFodfRFu5r8htYEQSHtrbcbJqaHaCvnVIN0DDd
T9fD6NeAO0N/XVrW9PmfSeUZdS9Z3PnV6Y6CEzQeyeY7UoX8NdlGnd/DGb7hvvD3QlXILWiXjBsL
qJLVjTarzzaskznE9hUmGQPG//FhZlZ4HU1JyBfq04K8xByxQfDgEiYa5+88KvQUofU8m/IAkrF6
rY15RfCHzvdUfCUcwQubuLqgZj0gXnqfianoqUvdfqOellupxDbQ6EnbxWNDNIrCygmWqj7M+HpR
N3LKKYpSkNOQo43aJE5Y3p0oPQIMdI4ZO/F8OSfWLS6dXcrhuRWCbO4vdeDNyWnFhtYEArtePNjO
bLd8AubMzurGgZacsWirHaUiDKg8dVbuvbkoMY5hqJ7N3Hlag5uKXNds4eVWF//uqnrQegS+d/Fk
LMivrJ3Mwgs5vZ8eO+K5UzBG/353Ya/OEZOt1NJ3Ytb2dyJiJiOwGAPhFYo526Dq6hp5N6EX6iJn
iqArVY+ltYBvGrMuEUfbzoBNcqS7MuluKGdNLjCijj3BZIlzZq9QPoui27CHjpzD8br1vKYOn+22
oi5NslAVwwxFWLxzizDnwRniTlubnXwnl8miUEULQ7HZJJIfqWd72kXKnyEXPR7P5JSUxrNos/Ko
lrzl6YgACDDXbvOKQEF8Dx0ze623iqI5QKNqqa5sbS4z3uThRlfjP8yelB5rADQuSAo0FMBTbJvf
s912sEALqj9Defbd3f9FOpe2UgfK1PSA8QWeiSvaW7cTfeEMKPg+LBvjqGDKLaVnjTUAeJV6GHCO
pzQdpHpRlIcudHHiqEGJAunBJtLJmBk0cIDUzuvkwHWg/mNoFf0tE2gz/BqCw3APWS5B3Qtd0oy7
3DUz5RAQVtn+OeGBQ62C8124KUiV5r67dlH8gn2vc3CV9rc1iq+iHl4F9t/XE/VP1ReMVEDQ6eUu
39EewzF8N6K/yvyXJzISO6McGuPfxXUuQYYtZRCKhJBlQFXPCFB2Vd7Tu2WlUR0NAhi55Fpm1k+D
WP/MZmpxPjYDtP5QyjIUZHN9b5WlMyrAlmfU/Knv7TG2zPbaouU4P9YTGvH3Y+z3DahdF9+UYHNI
nY3jDai61z+BXRBOV5XXVOeoRXKgfAuPOfZsbOlNXh2tESAiuqGs60HpFPWE4KA0bAe/+ozsrmrg
bt5lHqjURzNVBvartOPv1e7Lj1sR14nKU0axBQu/FjorWmoAmlxcWMcra2RZo8R4ILucrm635UdC
6Ydl6boWMPEVFa+62IpG4wJoj4OjtimucmVninikh4NdlxyAA2dElmJJJYh5pNiemC9GOxNMxiDJ
obTZSWLfOrh+sDWE2DW6eArpk51q3cGzb7ZdXjg5YWGVhlocEMmCYSUC+zHXrq1xei6hMjBtDKKp
m428U5LCR8DxaF6x3MXUAURnH82ZicT9/emhJa4QYooYy7lF2ytkmK3R/NyHr8ysTiCpAwwJd4Mx
PyiVKW/QH58fpWOuUdRIxUTnVl0Sm87bxTB62ubuWlF9MNy3Q6AOxD3FUyYqjpC/YMJqTrMPtts5
EYdhGgRUXtn2DgBp8x6K8nAQkzUM/1pKK5P4+AsiNPlaIJorBB5QRkU7jyaVuBwKOp5laKp8Cfxz
Ze5u/4H87byQWu0AfSHHTUwRUJeM60oobUBLDHfzz9+UB8EAa5HEw14ckalU/lT99BhhOKQbbUOZ
29SicEbHGEjxYjdhHW05WY+Kq1/Z3tlfS9CGcHzPePuW1bY+3KRj/JJXN/BtK9nq7iWa4QZQWSBB
uax8n0ah7f2cfwNIPsngGfCyczSLY1AB2GJ0EoCr5oz6RbLqpMZUehppmKxnt112RLgYMQUe2z3e
Dzim9V8H7wUE0fvS3EreV46MEdcgLixScg5y9Sw6jGMGc4nyinTdOgOZIDD6mA6C/yVf0mgEXo+B
g9hPPVSurNTCbbA5GR5QTJ/61FohzwzI+9H0fvTFDbft5ZtFvE0vZt8l7/g7oSewua40ffNTTW3S
UMbJXFxvU3J383YFECam9dNDv3iBRfmzbANY5k9BfDUDy/5t3NvAVGGuo5xADbwlT7zqva8/rO/F
cTddYbaTGhfG3JpYnUldngnWrWLBwXORbIrFUFgq1zBC9GDg2LNjGDQKiqo4BD71Uj9raq0mRBQ0
Fl+Y5wi1qHaZQAdZIRQPMM48X2IEUMek7Xl96a80mSlLb0xIJY2xqiYr4cNIfxXHM2bYho81X22O
u9SJ/VOPtrzoP9/IbWSq8v+GXKoBavdW9chCqAusRtgE8TCM3Q+AYK0eW/SnZcdyINiAR9sa7s70
ezm8dIQk8Cv1ULd4kADhna5IN+sf/zdPgobUWlzyHAshNWs9amxh53n8mPF46YyUt9I2uVzUXrnv
3W2WuJdjKqBuoa7h0JRLZUR/wucbrQG+5jrFOx6kZEewbrIjTVc4Sx4Fk8hJE0Xs8XflLoakE/r2
tjKPv60eAtOKoTj+4y7Qy8tTX5fP+BZX3m4GcDE1mZoIo48ILSs7bkCjpLsGqsun3TDLityI8W/A
JYTuR/7/vg83/qHA5HAMDHuX8faEkHEXVeOpE/HB7IOWhCPaDgmF5+9ZjYjoy5Z6YHRmPjLykMC9
KWcfYvQwI7zDuLAVsncaWq0MZJaJnkHrUOf6MRdpQwsk4CIvzYybrIIjniNZLaHLfpcCnnHhV/Cw
AHrpXmlF/rZV8xwvadMcUY7O7gB1loH3QcuMjtZMaqQbl+Z9yIE4z2TvCUnqLlHeGo+N9hvsUcO4
X+Wd6r4HEmUC2rxh3wdmcQht86JIYCkxKLvaoyLUQBZbpEP+D6fFr54ljBzr7XBiph6ltTZ/LXLc
3hUf2xRHw4oxLA5TYg+DmqiqqBPgMBGItLasTs+3HEQyaPsUqAMiByslTmu+l7cTrHl6200oAav3
XVqL3bhWsy7M4EnVHidb5tOvNbNc81HOdirG2nlimHLPzNkmjJo+AyHKgBCE4uWXFVTUMDW0GrG7
Eyhg2rmiyRDkgFC252TBkfDqmqMrMZJkbXqTCKMSoaaiG5100TMcUahkTW4FZV96Ijeb3f96tVBz
LaayGsx4xydSWGkLIaokz5oMTGwpBoICaFenNem9lcCfUieP3/BL7oM1frJ2ibFuDpFWP2tPLIST
8Af9nU85x5r3KEp5VZDbdYV3PjfGfN34AGXQWn6rrsqXuJXuGtu1cU6KYp7d1/iwIOPSVeD+f3Dg
aicBMx8hqXGFhww8M4nvO03iIAqcw8CV6Y4H7hptOk/YF+34pZLHUlurUufFgVdU7zi9EHTqPVrf
Gm7cKB+iQoZZUHxowv4CjnZBPeIm1KnipT5MreB/dn3+Erg+rRJg6QVQbi3m8Z0uVITeq4HRwMNY
wUIuM+Y/e1xA0s/udRf2KORylJtYCXgHHF1h91f/k5xpMBdqWONFBDoGJJ02a0fa1DbxhX0H4vTv
B5fuX8XwmEjHMOwqfkEBwAbnxSh30ne1tm3mbTpmGJhvjwEDTInp9Bb0zMaBA/rJt+p7TNio5RKI
dsP/nzN34+wcbnwpX3Psv+7LAqIXw/P3ebS+TSxVzgdHZ9TmUe//eochsC7hpp47OyBpCoSGYKIV
eqdvlbpSodHzHvY5lPBOkhdQyft5Yi7cly82F/OBA6ka46/aGp8/Kw4Pj1XCsExDfQBXEzT/lrqn
3fkHWcayAf30lAa6EYIynnuTjxgc7uCAFsBJ7q45FKV8sT7sjjejKdykzBOTEbwl8mBA3JWNKZ3W
ZUzChBGzkDQNHSWG5BSBYMeRJutO2i/gg2p3p1oQjiaVYYZEk5oYkCPvTg2bxVUBwc3XLzGZ9D75
qlBS1c6pBi0liNVLmwK9O/79BPMlqhN9/g/9sPINsjiFfh89ocHbMMbzpK7rQ+tuBZ/FZoW8KfRH
kgGtXm2kMzrZVJA7RXCzX4zYRqhjzgAa0ExsTeDD6NeAsgbcbKkxKzzXgDsITwlYR7eCvLApk9/c
ChYqJXZV+4clTuSmXOYls9qIdjXJTcdW826fRx5wXxxsqPLkRBX72MNyxbD+BONzi686opyk7O34
8muf1qSeyDX+ya2O+25gkKY/R2WFRkNSAHq3sv8U1wgLUjkmhnKGmo6kwTFxHZy9nslLVwmwr02g
D0Qbkq1HjcRYtmH5RI1ErcLFjBwcjxWUP/QoQxj7wtSli+cjVteSz9jpb02Zhz1Zo0TnJ507OJRE
g+1jfvmOpPmKC86E7KMxZxm8xPUqBSK+dGpzw1gbX95WQ5YkVSdaF4UEH6P3RAQPL+542B4oLbDF
gJL7aS2Ioy93NFvpk3hTFdOmLBWke423sjlOs02ZzfW231TKJogvqjpRYakCtuWqu4K02nQUwDFy
7mhvd5Bg7LDwN1Ay4LJt+cn7YLMxoVWqaw8JINaojEMSWXwsls6lMD7LsuKG8xklSiEhQx/If9qF
FWP4h/tflBUZGgor/HpKYvhhf0OftyP4xvhUmIX4hQFVF7PW3QRzZZYI9ej98TmXOdHdczRbVyQe
imX+YF1H5zou5ylFjDmbjUPkY+RMWuVoYyAiD8dOdS7Nol2g0P8aM1IbYsIT2jXWIZG1+wqfMcCa
0/5D2ue7lpPdzr4NyrT+WExAxYfBvJG/Q92ALPbUAQaeZZBPkmAndGWQR/vQfDN5Q38oDLKLmzRq
g/MFhsAjJCasgFosvbLu1ImPNuURQoeSc5IDuefr6C4eguriQ7OaoabUQmhSoVhYsModJB0oq+mV
yp70rK7KA3lM0NDQivq8OsAiF2MSZB38QIfPSAeh5shp4fIFjyoE62+rhMygZKtsw8MAgtl6DL2E
7cVTBnfwCgqi6zM0GbRN1KDurBZWS+izstBf9Gut8zrAiFGLcIVykJz3kjxZ77RYh6+YlCgvG/Vh
MK6ZvMDBtFtjq5qrs4ImhZJUxK65QWgzHkIyC+j96ePWHASr8gbc5bm/rzspWm/x8znsv3gdYrOS
AqAxI6W4rSWLjY5V3NPtCmM3zJMAiPiW5tdujtHzyZSU2VpJOeCX8TUTsK+5k2S4u01mKVhbVa62
VR1u9fFsTG4/PnXXnL78CMfWfPk6oE4odvaIIKgzw3VCqh+k49z7JVsTeU28gSWPk3r6jv1KfQrW
vBES56DQTZtsDVNe2lKkR+cqgiDQH+Uu/Sk30AgxfuYJR+WXJVRz5pnzveU9FF2lQfwrQYsm8IbT
qdelwVo/thQYSBQAGFRBcma0SMkypa9N7uVU8lvj1rHu872THS9YNX7E3DaUSIijomctXt+Sho3J
+6M0UYlhZ3k6a7t60Z/fn8TJjaqnWMF0b9qxnB70Q6KBf2dQuIB9dW61i6Gsf5PONB988qX0rM24
QPjWUaIkqE1kukjfU+7lOH0UVUT59GrS8IL5isbnaThueJE1AiEowNG/3StVoLnvNqNr+dbITHYg
YQXB6g3gTYQaAVyYUEij16BlxELp9nAF+L4qa6LVGmm8u9LGj2ogoGB0DfmNQTMtDEtP4n6IlZK5
a/P9RLT1q7Qr9TxdlhGb5pz1QvpppjrUba0L/s7Ae5fVP9d0437g0Hog193l7KLyOOmpK5xlTtTo
Qo+kBYOkDCErQ6yS/drCkT9Y3TbqIUnyspvMt3EwSwlI9pnPJFR0j5nwiBV7L98jws51CsSSycPc
6BUve4ljhZ+T8gWSQQCjUSogmc9lyHmViOXDwio0qdW1iUiAfSFL6RF+RuyGnq2c/N8v4Zp0di1N
1mpYMb1hkZqiIhzVqCdk3+b+SY/8NyLfukfGdC3i9iyaX3hiKSd2TPx7KOwl5FiTU2K58ea8fMWd
mF1sJw0d9E9DVzu9JyrDJcf69hQbuuZDIfcllno2dWPavxsbUNCrioQYDsLcJWVvuzu9tPmRGiG8
AyrWm/dx4tjSoz4KrO3KGP2ty7zSr/RiSOC1E5EQLAYV/s1tSkWd2CedBZUk1VIkXQNilZryDWBD
UqciW0xMrSmulm81zICRZi56EipAViv1woW9QqzpRT1CrbtaJA6CIazcH2VTUKMgaXoyDIkBiUWf
BkFUuZsZbvUGgoPpgedV98MhWiwW+4EYXOgdApb+Z1mbACedMcj3lw0OCGL2u1Jme9TVglk8askX
Z9J7qa8Dk1QvJNDFCezPWKtetcc8QVWtTLUpHq1RtQUntBGHBz57SEBLZiQQvb4+oVKSBk5wB77W
jpG77PaexXTSHLmwBA8IBStKvATFSSnJvOQq1xWCbp7kmsZ2oCpH7j3mWdxnlRNKMlZi4M8DOGit
qreCJhOPzczcassaaKIhUI3Z2eBPapLK7FqyuuT4wd19a3xcTzNGn5Bp0vICayVBuHUfDS4DVuGg
VacOYZp1z0QJnP1SrvVWd1hxIGMIDwE6hy7g5TLu6Xrp1ok4OZ2mMdc2y+ei26SYMbM6BHvEyZ87
+9I6Cwb/Tl6PT3ako+Q4McpFBuQAmdfX9Fym5xBWGYewGZsyqCXozomsgOi3fbhLxLc2j7Ey1juS
UVhC0GPEQMI1My28gN+ny6EoBgcbhYG72fnoEqb29ENBELdK7E23rih4cjnnxqBl8lkD6noSAU0L
0t7ugN+H+FjeTL3MI0bpj5Tj/cgff32014NQV+LvLZCdlNDeLkCHXry3UpB/dQHAEkF8uT/koA7L
T+vaKtRKc8Xp9M8+GIbyndPY4C53TFHyQxB3j4Yd2IT1C82r3s3odNbLxCxa3ANL6WPgN6ujXyCw
XiVF26FayHR4eUeVGY2V/asTRcN2I9PUSUUScufhfO9dffTbiJAnVLdvczyKHPqU4mKB+SfkYNVi
MQIU/zmRRMy+4atMxtt+BNv3ITPkiueBgLYtwYgG/jjpUfwHn2RqvQ/y8zTA2ys/HLoF+j/daTsn
3r4Nu7+Yuqw2JHibT9dmooaonwEDaaNqTIa6O6u/kNHahqdzhuQEAYYv1F6aQanq4T9aZjPwDts8
LQviMAY9pQRBSW3S+GrF9Qp0x0KMDo1eLLqndU9pb2rWvir7E93X34qlR+ZdbU0oiaC8RTUIcCwF
qOX1LywNd++RsipfwVtv+WmVWoomRstFMHkY0csDDNJTe/BDl+FARLPDTAwMOTpDmilu1ujNho3d
iRBrt8v7t6UeO+HBnz6zyWIYHUJX3Lli81UpUVP4I8fZbe43nB0jDOX5Muw2bC4HmPqlZJ5g6qF7
t4sC/6EpUnPXh+hhfoRM0sP1lZfRrFBWrgMeQhb1+VMxuMQ92+EPDcBfC/McNzw1IqKnEEybS2hW
plKBI0TVtpZ5RG5ijhtZg25OLN5lo/CtFckxa0WdX8OUL+f/6TFC7scmDlPL05M+OclXbueXQ2MB
5b3dTTYho2wyVs8PSl66wpAHfHrXHSDQBmVycsxK3953bl6MC4UxRDljYC2GfvLocngWGoZ7xvLu
KuSezadLTVDJZrGlxc4bw6aP41WXqbRImkmYiM/qzUpMGnlvqxYP14LE3520ypfrBxWtcZAppHMr
4agaAYRjgMPCJq97ZIdXIf4gBsYvE3bZ60/WWenrPNhDsWyuFn2noiIZdY2CUaDwp/6cbGN4dSbn
Si1O0jS5KPl+3e7nt8lNhWqUfwXnOnwceB+tziLaFY0fTR4qjjrkJwy6A/F7e6e8UvaXuk2nNXM1
1f0N/xqdGR8dQ2SEBPsdHrCtyCxlWRsIulJa8fUji9mm+gFl+s5UkmCAooWElwZCerM5Xc0GG8wR
HJmPxE6FH/A1C3f/zLY3ioAFXLs3T2X7vilwaOMfAkeTOSqpfZJCXT8B0yAd/NAK8InVXYpqJrxp
BWtm/+6nLm4YCJzXCbO9E4pRHP35M1Qk4gFCQw1O+e/UmXA5Lckk00qpeDv5tSaiUNY0grrcqkFI
7BfcLn9cEOcI+UO0E2o1/+f7YihvAEdz0nSUC8Fl/x2vf9hDTisSbZk53YbKzYnv9Jcw8oF6lP/b
tT9q4sSo5P007EYjt5kmSm4oZ/YQXFK1rwPPF835YgwLMI1OV5yEPQoN2ojIa5Goy7zaiiecF18+
umBIUn7NI0EwLrnB2gzyDJwMjCnk6EZcTyy7hTaUYRxa4kk/QUgkLSkCZp0pIJA3p20IBxMQXAk8
7SOHWonhoO/Dwkn4fVF1l5JOgg70gVnZXSjkwHTL6THL6NCJNVT40DHNqrcus/NdqT+CQHUtjzvk
Zk8e6X3jhR4t51YwajcN4lbr+NFK0IvRHvyEqZTBcTyXMDQBe4bWkkDkBlQH+hMK6rn3d+AIRFiD
g0eSQKRuUtdt9C/fWk+5gN9KaVpaonMPXFvObDdvdjLJVpShynmkFJSCDo8/GihRsPTaMZ9UjzsY
wzaWnWoZAp2wf2Lj/PEK8nlTgMfzVFUo0mD33EP8kPiGAssrTnBp+Uk0BeTXeouarEO8TWJaqjJn
2rE5zN5xrdT54g0Urk23NwGv1qcHhf4rkvI/apCILYtj0ACbUenqwq3wbY1OzdgA5GlJgkYxq2gM
YBbAHel9UCzJFyqQJ/R1ESWugFsi3D9Iyzb2MgDJIJNUjcZtzERhsfZLLu1Cf8STS4NcIWzYPoaO
cyRwWVF+1WZF//TbJLTiNg6M+88UI5fheR6cOBHkFfHJltyP0linRg1Vqlm8QCl7zb1MTlmF5tlA
JKT+B5U9u+Fhroi96RwCbpxx9ZDYtJAnlVv2/YcMiRZp9v8yUi0Kc+HdpoDB8XXPrKB+vXvXmkcV
KOHA1QZTAOpU+eStmEn9ZAlRhD1fppo6f4+elYAt0GY0iZHitM9QC/3uBl4a6exXDTc8cYMyNpCW
M7HMlqrJcdlZvKT4fb1n5bcTnb278D7R6wZsoVRL9OPP2eC0sToB+CEwfetP9efaNOk45ZPZLHZA
v69Rhf/IOAMomA/RPollxMmLi2ZtJ3hOQX5zgg4Yuu7rpcjwLDT9u1Xz1M5MvbZvywQ7xYL5o2tI
bfcCq0vHYG5XaZ1XJS+qTIBdKXXLw1tQwPmUWO0WCl4lwgK3+NGsUZDqjkex3S4czYnB52SdQBwe
bsLU0yZoHVFTN5pCht59VI7GJqMi+j3ulFX0OQOysPu0GCMYSrzYNy0XEH2OIsf9+AuqYtHTsBwr
rB57lgdmH/mJZ9gXd2NT6ZgpP7CHExrlcRVuR1g4mplcazv/9i9WZdYZjzpI2RIs/7aVGvxXys7w
Pc7PZouXFBnqh2yc4TlO3IG/Myt5t0lQE64lZCGiZPZcdIP9M0sEeRo/DpW0ZlF5taQmnsTvMw2y
qKVsP/SMhVrs76OIo0MWfb0blI5asO50jH38VY4Sa2kb/orgAABkiyoBweUXBhrN5rXTFzsFo9/j
q3lb93TW8tpITE2+rFzOxnjcPfDFmQ4R01DJJkJzp29S4rCLWUArcquY4XJhV/t9w4OJVgRVxvyg
oipC3hjI5OEQAzHPj1BAXv+N/wWL/NnKgelqQe579riWbotVYXVOUiAmAtxcGXE69kKeOaPP8wJ2
2qvNuhW4Jj2gaVtuSvLkMWV+TN9x6QrmdoSJotITaQi1R6P177qCP464GcwMrAaYNzSFgiVIFwvG
5SKq5aKCxJy+nFF/0HTfsHGz6eJYGduVjaRMtUH8pzbwcXzI45e6niXmmusZ8OlGp4s6LWep9sCO
ImfEMA+8mjhI7bXAH3iNGNn9NNfXH49zTocFOUzEpd21RCC8STP81EeKLlhmSJd/Om9NSqQm4wVf
In2jK5LTGYWJPfwyiN8eEaG59KZ35XA+LL/GdYz6ztagopckkJ1y7Ai5HJl5sF02ezvfg7+v858i
aKIIOHGt4CWDwTMtGw5OYnopFj7x8mBmVGKNrD/ZxHhyo0vgbmcUpqyESQQXRhD9rqbe8nfiMOsl
3IwZszChXvgp8+JYjSUzCBz3S/SORGe3MMUJdVm8T2DQYumcvsMVYsuDz9umEFsWg6LxJzwqEr5T
xqMsjL7uJKgq+fDwQJOKy1LRvOACMS12wFzxLdvKY63rK9jynHZcwavTgllejNh2EdK0QlSGWac8
bytnN2IjxdPeXD0GS7pmOGUk6dHO3awSXdq+O7uT4oOIgFhiN27RX/5Oq9PInjgZJlwNJbdbabGZ
jXQwrqyK5jFZlWFpNG0u1A5EmW8eQOsqIhy+sBjH1OFUSHNfPtTWt8+HfXaS/mq3VQPEG3z2WeHw
EyBJZHrnCzRDc+N3GPuOX6/SuGYx4M+VNGOL0UTEdyAqNeNspTswbqZ+caxyoQ23SVQA709Z6nYO
z6Dpzt2j75bEtKrlxIyS6LeVfjlXhWKr0YMqj2y6MyiXUQw+ZjASjo3/a01k5xd24zzjhQJZLZCo
3mYrdKe8v9djkoXMo3Jha1Epg5fTnlPgKPf28OP3LDdbvaeBBk+0o1f7m+QfTOEcTIDq/xZujaTE
pj83p/M/MOSPyO8uThafT7AzLNTGWZEXZ341mFMl3kEUVnL/pnu5Xgr8OqP8tuftRdP7gP3L0d7r
hddwbOTf4oqJC0tcrtpFGw4s0JvgVjRnUlU1NgDSSZtn1NdRop3sFd3pefNU/rinE+wQmYoajSvq
9+N3FG7cJJ7SrpEZxe1+Mo/D+Tl5VPgrA9sH2G7pNhESI4M9lJj+f/pbrHiX9GsQ+0DT481lLeag
DxyQNE5tc+xEy8dHeF33nPegOi7RrzHD+RlsHHWDbLSAfeztRB6XBHHvI0275O2MJCGZH0SAj2At
M9phXh4wwNBalzsQ/233w6IJdx4h3XdJS2/HAMHYXhfopTx02JpQnuAT2/JBF1DHzqumEq0nu8sM
PGA/39jrGA0L8h30096zveKHGPCmpVYIEFSl4M6kmOJFnVzNU68QhW+tFg4gUDeD8HOBxM0Du8Tv
3ejPjp2TO1D0qO8g+o23t7XjzOQw38DiuEUydvxdiBAvcJbIOxEuhBZx/fEm4o6A6IPvoA37yVgE
2Nu37p3JNL09AE9+3XtVyKTir5vpTYJS0eNITpo2yor/OU6QsKh7q3ZiSgp6V/G7En5B+7IHqAnO
BBst7LoQFxEZjKqrpD9yuKEsWdrWcz+edXEaX0J/63pAXAOfVgg8ctSugRDaiSzSGaCkFbe2d1JN
pe84axR1IEevbzyqBlMHFH+Mt2PRNQJT954I8cW4Erer7jrvc4B7tYJ243gIhWXli3saPAqxxvtW
v26ExS0Wiko8doO0+y69AonsMniNPM1uMinI0QZ1bDHDQiRsZ03DiK3dwQg9UP09QVYSMcX0rtYN
hAmITR03tYRetcPeoI8SLZYbjMPfTjvlnakI23TwQi+/0mDGBTK+7NF4+XLcE/vVbI0JEX49r9i7
9vStMeVbRuMSg/cWyc81sk4dtEchQucKOaCMWj2/IIcct+dBBxHqbPrPeFjZW39xpkMHu1tQQ28X
oLIIvnYHSxPi5qpAi3Ht2JXwymozYVyDnL74Qn2AUdn5fPOBd1T/P7yv9DMBYYYmU9NcyUIrQaxW
Dg2LEoL6lsAuABDU/EfpBN3wWAjSSTyDV16BykvvhwZGYDXwagdNjRtTdLw7aipeB6FUr0eTxnTY
uHyc0ao3WjWnjFtnd5mVQkafcXKpfOWZOm0TmyvvKeuBVdMdWrDynBu5opUzwsP3hadn1qVXwD0j
JmlSVOPHauc5cq/q6JS/U36x0MNN+JtPCdf8kACB1mMCF7Y9GtS73h431R2QrwmikImrBeD52wHG
bi/TX7TVHtn9MDsG+wgbjpnzT10D7m7PtLO+QThbvxt+QKkQeFcS3aDp1Z/wa3LcM1wIPG3bAZ7f
Q0sh0xJroOCjR8SqNSWj0jt9r2VUXCuM62MqieUF0hcOfDBBhNgWDXQPNnsV9qXl5AdTual0t0xr
LjrugHVtNJiEAEJoaNfADtM+bsp8+AXqtBZkHXW3/7UgB6s3wkBlzrGKv2SVketrUT/H/0ZhZlLO
RT0bYTl7jz0wnw75F0422PYx0NGl+vOdjwT0MJgyNzwpuRYCQz2lBOq+2pRe0/ylakE4MCAuxBBR
QgB16OgGIbSwGlIyan30ZYGMMPD4lgtiOZ4Fmd0BCcmL2mFcnz8BJ/wSUhw9LsqzyH5yQJzx2V3k
yHIyoH/ZnqkNZGEypUggZ9jr7816nSbZf0UL3CqvEHmF7Wvc+KbL1hbvKJrkkIl2ZxQ3O2hZ8wN1
UvU3VmZGX/pfIL3rVC7lht++GTXOBHLxomOIGBckcIslACArOFKEfAJ0rCbTBV3o4h6fyMPohn7N
K6jqBgAHBCQuni5L0/ZJtDoQ17uXOhCJTt2LSJZYJQ9AohfNNWhJDKy418gNdDNYqXQhLfN54zez
o52c4qPcDAgwdBSWvKnoSL+Pt55fIKo65iy/xxm1MZEGVU9vIOVCErXMO0DqkBqCqW7OyFoPkkC4
7DCJiBhuZjL2M8NaJSfTjORizZ8AgUyYxHxKQkY/i1lnrFR3qIYPXINXYi2+pkiEvnvvSEUq/I8i
pnnomBsS0KjEO7IxfJnmTBjGNr9nQ5v/cPC2IOi2YFxzOFvo5iYqBNXfdJ2RSpUj6oA+ouWSvoNd
g8JA/RSLE7deqbTIAWdnFN1i36r+JD3alfxpIl0F0sYVnkNhYVrjmdTenif15yyAviB7k7LVB7OC
F4Hcd6vhyjy8NEZmqCKs1rrDuYjpULif8BQrQSbWr8aBu3DNPbZFVVkB/jrOwSv/95XxGUipqOpl
keNuiZXURYwWr+wMZM52+l1Qbrhodpip6N+miV7fEwPplfOxOX+EQzygvSrFuvEP2gACcoyhpcgJ
6T83Zqf10jAtnaAXIvij+eMzu5yw42UmwgxTZ84ClZw/L5SjbDJTGIrYqTu/K37ocOp2qfWxBQhn
tBakkNMEDsUPQrydVYHcYeaysFYi3GvDxQrcUKP4kD43YLKhDOu9l5on1kd3tuBl4+EipPdE5xXe
5xCbO4hoh70bREhpMO7c6fz2Ihj3GT+MxbeiCMHl4rKxKGqV1Sq0Os0alzI9cciwGDLuuReqyGSQ
7Q3u/tQECfwuACn6VFVzC8tWdKHch8Corra3VZ/D1FlbDJhPhUg9H3rT7Rsm2R4/Yra0weyJxEbG
9TwUt/QuTZYx1MeSvJHkaMNOwfVYiloDxpCPvKQYS3+lmbOPXxvLLTiR3n6pEmVpL2VKYv2Iq+cL
Qe5kR3SzR1cZvIhTiH8gzk9YmPmBzqiGMsacLFUnWkLUeAnDFwWvvcMJcfHb35f8w1Bz7L59cjEm
44XIfcrKu7MaLIzQGUBHOG7vsVSv6E5Zlph3zzRPQgDL1iG68EywCILxAW8BmjuNT4T71wP72RCd
YrFN6eCz9gTaFjkSmw4P/My4Q7smTA+6fK4ctNSZjadM1xRrxkccnLNoqQZeAoN7DGVol3RxitFy
B0MvMe5+ZrRkq2j1BpOpis3SxDnW9peaZHwGUOx7oVHuI4UT9xhbSJHCsFbGzgC7ryIcyXL74upr
4AxZwpzy7ctQxB70t23mEhNwCjfTiHfQXujWWSkhivwv/q9RsXCsfgpHXGKEnNzlFX/jesYcb3v7
Z4f0sivXZsWUiMj9XMj7oMdYXy33VLUGpiGNIaZDlwFWSBAtM979NJaEhpVY2pmsTYx2P8WCulpY
nrCn9nrpjU7C2Sw60IlovBt/1/OxANtjMPs/bOfVmXIcQKf1eWWm5w0Bq7ISUL2DCau9Ks3UWqVp
mqQP5kLa3BXbQOMyXfU01q5RIgD0iVMFDTysDYkfIr6uojk3Hupedl7M4OtRbLki5MGs1q2q69k5
XqgqJn7xj5VORs9g9AI0NiogJxswtKeuOOuvqWZNz0cKRVFZtPXrrWM4HTRTdcKi56liu8gipLNH
Qoa6SoqZE+CU50G7zuKGRLUjVOPW1anYH1NkqYUIDP61ErPNaMPw9LDj7rEC+1NnOH7/gHlKAbL3
Cv9XMuN2ldzWSJw75IAJrNj91HtX7F0ZJ7DyGofJlrRFDYWJrNQ32QBlRBGSKiQUIlGQU+Usv5Q9
tXKtDfG6Jbh4rFIcj9QFEPWAuJXX8iX4DuoDxDA2oR6ZucxGK5uB7mqE1Iot4OtSRgEBL2tqqQJ3
XQO4rG66upzbbGsmN04HAq5zBY9Te9UCw15xLUIOkLAXymtCBWl3PTcGIj3U4D/Xu/wqzoy1pk/W
Le9l4wO7CLOQOM3IEoJrYezAILJJWcL0vzptXU/+mQxXMnhk2PZhukW7Rb8o7HTn/FbGujKZFtKG
NBPr1/kZ9uXSRu3Q656R8qp/HrIStTTfnX0ctgo3JnUghWlN6zsPPTduzl17Pzbyxcx7Sg4JCtLv
Y0vebFw5qq9FGT8R1vhTKXkNUbCEKN1Zti8rMreEqRY9qwg1C19ZM2Cl89eX+4UlCsGILs2U2veS
8I+RMj2c8iaGdL+Owbm5N50ztnTMgY7FsLxiRju3JPj8zy8ZEmt+RROm+Q0YUSgPqXXb1yj4ctp6
NNkdtX5QKgYuGLUSpWcyGPYjAy2CO1NXXYbwrPvvGZhQYjr0yZ83BXOfk3zAcECF5WDRYFvuFLvl
K+0R2cxkNZBd8urs34ZIs/6Abpo7GZzfRNV6AP2ENazkr0gqd92+tiGjwyMLvpQN6GI0QIzv3iuH
2MGPQG1HgahYZaDRpQj4Jx5HCl+4SmBEiOLecn7IxXV8mhH6genUmdaEdLU/4VfSLX9Z3duGUgnB
E7aisQ8PtQEKVcKQEtibTcBaAZVrqIliOHuZoTuGYBiFNCeVUHWTM8pfS88r8ixNxPLV3v6rpIWG
1PSYTdUF6XVLeAzgU4fUsGMvixX+6jmPrW2A/oWAv2riUp5JdyMWMqsSnR4pHA/z2HzIpMM9be6o
11CcVxFALjcD58zssbobG2FkYAySQXeA/3YFCMXPF/Rn7qJW2raHkfBqy9M2hvpZgRH+etCIu77r
CVAoWOTdO6jKtPU7G5yToxc5tIjUmWD/BdLt9BUF+MsNWU5rAenm4Du1485QPyZ/7aXNEsPsDOrT
4U2/Dk6TOij2uOTUYa3Ow++ory7mgphnN9suturxnA2Nh3BglQbPE9T+XH6lQ2uV4Phwq+PaHB/H
DUvf6/mNYU9wGCo4wH+evZXzqeUu9rBAMly75umZmNptEixc49VU0UW+lxsn+j5jHioT3eWkgVVs
jrv4VfsIK/AgPd3zZYa6vuc56AcJUqwuVER8jV+ZbsaYLXn5n13nZkAMk0lh4F4FFK1GJ9//tmCt
Cs3P4APaMbXeK8ZgImESY4HMGBhGNlMW2QTqanTuhiNp3GcNfyytkD98+Hte6El421PKshwh8gau
2V8DcjbE+ZlXxJuVcgrD0EcPgTXBv6I73FE/CpAP+rb4oDk3UzvTkDnO+5IjoDVOeTYHvTKYzNuD
2saE9BrTQTMSGS+OwW3WYQXXk/ZIlf8slumYjtf/YERd11HqjUS5aa1q+Ffrx81PJpxS1qeZ0g4C
7C0KpHFzb87glZr1TU6uN5ZoN/3fEM0upEOAmeUB1j/ZN2kUk69Yt5XbYe2Wt73P4bUD5wqskGZP
ZBeo9PS0dwARsPUX+MiVemJ7d1Y+ufOja86eXIL1isZayVl1sYc7iDmj/byu73TxLolc9ZE1jYp6
pAWBfxkeqavNUmjPvhxq8gupsMBJiIGRbARwH+iytf+9uZ+ZujHDAVdommP6+pNDjxg7DSbEiWwd
o4yjqUswKTyMCMkHGHRFOQuqIpWvbn4V7ow30sgzHD/BhShCjR5maxDz/nP/pp0J+nGv7zkHPVl0
f0t2JPgN/X348aALTNQ20JuDt4WpPrtqfobrjdn2MFDnopyRIXZdcLelLLI+t1QKxT9mslDSY7w1
2bXX4nEneG1kX5j6CdLHqTisi4Vvc8UVy1XTstgHqA9x+Yx2Y04/C9ft5c5oGAa3Az5wvyL+HNdI
SV9jZa7PybOduhT4Cm/GOo0/xIBWByT5GRCrot5ViGSlRI6dz4jRTzjMEXVcv3pB59a7m89wIo6C
kuZaJQuFLHdAvxtBoHUTr0Cqi52ZHvUO3WA0y4kVoo9O+gsjJ0eKuvc1xyPI6OASx16waPbtjvqo
QLi+bBR2e+aP48roGqyVHWtFyNMmkZExH3sPi0roC6y30/yPIjwJmRAaMksyR/PTVflx16WY2KR7
JB5PY3E85FM1rkkmj38qp7YxfIFoOR9W8ZBFku79dD1vsJmhw/nvlWXrqHNUSHv4v5A1akymH8L1
rNewLTevjlglCAMlZJI5BH3/SkoCmTnxmaUtChoz6N7TtCjKIUiVScS6lMkLNismqS+IgslVTZDn
WDScZ68aRxKkqbIaVY/cDaiHCz8e91Ww+YIQkeIWG9lh+gXohzt4pcKfJix9u9n50SmkK8dH6HTu
QKmkfaHNh/jxsQzXnpoHDsr43zZhFozlrXtxN4diuabnIeM2HKVqsxlKPGsNRmGwWbeMl/vSn3OE
QMrCIpr4CE0UkOz9tAXStP4Lv2sXcAQ3sX9WVyddu7ge9JI1Hg7duN0QRibzf4akAS9CR9TV19xJ
b/0RDPjIOcu3mHrXY8+mns0xsYDpKn3j5iwFBVVpmOaoB6hAnfZ6szcsmAGwaXiS5cKLXN8qUgIT
HFgO7GMYunkv0+rwVWJhH1UbYuHl9nG04r8e/OfkiiG1QYEdMPQMBvT3VcCPrEf29J4eM8bHlkih
AzdaGHzltK8iddr36OM3grerFXo1vPG5FMQRVLVqIYqM5dr1v1MBjyD5qzSq1glGndsQ8tGK5oXT
CFxrXV4dUncfE4QdGkYgh2uCE8nvOpnbn3UQWPShDsS+ACNvGOaSfzihJ2dO38HWqtcyTURuDamc
o+XQtPwT9g8Slzi47rhwzQ7i7lfT5WIQfJPqxiMUzl3XBjHPINufmvZZk315rJuO2oD5yooW9nb+
mWkySamLGg9uTUHDjj0tHzz2FZtvZoYtNLhzffh8Ryou9AnWge0xPkMiN4L55MEE33fYILPlz2ex
SSGiGuE44Tbb3F8MGdFGlycP8fZTHq7N77HliZJGYNUcTrAd6KoFluqabmf0bNu3fPGzmeOFVR6a
HvKeaRXpSDK7mGDnE6U/SX75Si/nklvNKecADK940YSZW/1JI5BnUpKbEOp6x4ux5jqVsW8L239m
uvG99b5e3wOKdV5XZTRI5dnSwAl0jyk3bQVJXjovFj1EHXOCljjR+nfGePXV2jplaTnAoa2K0+Wa
ZylJ+JwRQ2SX5sMzCt8KdqSLydK6TKCd7uGx6xuuCOLy3sG/52GISby7M4VLuwtHbLQD6m4jtm8w
rtb9REe/QIBwTL/fUhnNxo2nxFa2iRwL8/FAr9fDgJe7ZDAkNUzPjQWojhLD8JYN22ZjzWedvvac
ITs/K4K/Ec3NYj5i6I0R3S7hEbFe8QHjK1zIzTbj7cf0YPeV958Zg4r5LgVAiVTelFfZkchWyJu+
FlxJMUk/DqGgd7zRYJk7oZf4Q+qyhq+/wlJARi/KTPJ+QV31DSR+irmw9UPpxCJ8U1sDExeBJIIG
qfLNp5S2eU+Uy3IB9BA7Gjuuu9Vp08mxfAr0ai1vah1GqqrmTbjzSsHzwGCbVO25AQ6j9e8ZPmrz
djbkAssmxiZ1AYbQAaL2Evz/Zt0rtm+6wp/5GHPiG1680VGqqB+IBeUcI8OzUV9qZCW3qyIzkel6
L1IjfqnIDhjFQI/SjF3JsGU4KHiGfCcJAkPBmdwtwwYdkXevnD/1BKBCAbuEq727HWoNeL1hkLBe
m1eC2QN0HxCgKfbDk0ns/TX08R5L7lUAslT1z/2ZEc0zP1Owi58+8KHsgc1DoBKBBdt/xw1gMUwR
olFvDA4qiQv67sDcOuM/65IifrUgf2RcdhOyOQ+tLtSrZgnCWYjxl3MIW4Mg2RIJsJRu37sAusGw
VNYrj1jKcPnqQh2bUBB2bajmx2eyXTcBymbaJ3iISCmT1ZTnCW62HTPLC9/LifQBG3mMXslFLTqo
jf9zrSmKSunDywEvE5635LDKKXLkWZPUERbTzwgogJVDWzzy7ZbQ12Du0gPzVmx35qZ9AY6tArc1
Sqs/ednRzehYABxAlGbYTs3U9BdHQkwDyCZWFJahsvwhzsp89SJ1mKi4P8DZ3HqORzLieYpUqjUM
aOpJYiv5VxY3s99ytduhwYBqNhu/LJryz7lD1ilG2FN9DOpo4dlneB1FbWiqF8NhhcpjDv3VVQLA
+6d3frIxgP2NRcdO2/y7H0mYHIfDa+TQrnPuNCtBjGyJHbWaZg1CtkefWCSdVXa+zJuUkMp8kCb7
1eYPtFtO54b7K2ms6c9/actD3eQJgmdOoJa8qm1v4XmNY8uomwk6b2qr+kcYuIVFALMKDT1N5GMq
RFSN2TXGj6BlSqVnIaG5PxkUWR7ICt8Edb5fPV67oTTZ9Wlk9ReGR22s9PlrNhlrM6l4n8BJ4JVM
R2zCaeeEeLB+/x7xK7/5GjgohNcTDsovKYrpY2+p1OGgauAUil0cqTMiG57jBa3OulpnlYAhBCfw
5kiC5hiMHeoLJo8wkSYT/xjz2D1HddJU/4o3P9yaDLePfIqmUMZV61HFE3s64LrqUxXtJ8Ngge5U
DNVQfdaSKojohW0dVCAKFYJWss3UEhkNJDF5bJUzjKe23tP7jClBLqDgQzhsBcXael3LiL4sORfY
N2X4+D1Ogb7YW9+zXru3UuTwdEKEqHAefMs3nSFeriEloKW0NCH2Gd9Jm4H6HBgFfXvMqW/4odGB
tGsE58+pDaxwy3QVI7efiBuRtjyPmSl4dExSwXv4F1vWOlvB6FB77UP0MFLgydKXrH8jVPX4z6GV
152FK4BCR8D1ixJ9MBulL1anCcB+uTRN2x3w+UEJ9XGIvmYGdoMIX3BSeyKUhppMHATX9HiBE3HA
k+vCP6LOfFvjoncOkFT3MwLoP4E9tUGfHeqh4rlUHkwKuhIon9e7S3XiZE0YE6gEsZn5YRd+JoEb
7mN2dBddknhyqSe2U0hkizPSxaTx3UeqEBdCx/qvTXyZ+NAKkkZybM4Ri2h1xPbbzK72DEjMY6yv
5P3/uRzFlFRrCigS5aDj/73IA/JHpZIPUxsgepb4lPPw3WmZ93XeDTgVCyO5nB15xpPitSEtXJnu
7qecNgqM1YZrF31ejnVvXWToSMiacC9wl7cuftfXj/ooPj0RAmmYeMtLUreL1HH+/FC7kIuHO2e3
oKbehvYsxQphGqIKIA2v++lLDUx2wJu7kCvXqFiL3Lz/b6rIuiRJNvgCwYeoEGEDczqiMq8XWmLw
rA+VxBQvqWF/WDqVSQrG5sanQXjyZ1uVn7Oa6MTwHV1glYGFHbZlYJz7+QNF/b9/RjF4I1OCXWSe
z4TTIreJfRsy0X6a9VQ9GELc3KlclLb2q8XOkM1iCMw6J82LAwIdGKUJ73LvL/GCwTT7Qp2/krZr
RhaQNzHg9m3kxv5x1W6lcN4K/Re69szDIqWI2F2halLtX1Ehk/1zhlkO0N7rZP+rMvIWAGEEf12F
0crM7sNGnVHpiAUTbbUtV25bKxDlTkZVEXKDlUZZvE1tZ5bzrI3sqNXxBFo6xkswPaISc9eMlusn
i4uJwjIu8dH0HMNZbhfRJZ5sHtMiZW3aw9VFQcDRNk16k6cNzrTRXE8Tdlzpqmmf0U2xqyjmH3I9
YXPsy5r359wsPphxbW4mYQ+C35oWSTauOubwnSjNhtbX71typ7T2Dk+0MrrXRpj+5jbe2aqsY+fb
y75M45qCmAqZCEUKSWyGjAhfz7NY2GTGBMkeju0MO0IyQnF1v0cRPksM9qPS3PMbWNFbpENabsNT
FJcwZW5YzXWfP8hjbllD2/0dtl+mTE7ZzeWVDOCvKur6Rmpr4BYiySeIvBXeOpZwIt2U1akrc5sh
baPagu7AZyRuNxBuhCSpiDSCSKRUOk1KLcoubehsU/DG6ZKs+cZ62uMPuiPtew9e0u36O3/KwtOV
5y/Zb7YhWnYvQZLBsk0JNVWiesiPeDmZ5DxggCoYtGSWtzzVjF9q/U8t9oa+cYmxFTiGsnW9Mbs2
q2LMiwlYJ4B7jqm0lQ9koyZ1+EcHWNUUt8ubz+ryOv5uRbVH0eDCqZIk7gPKFlHMciwF0pYOvAfa
bC9TfpmThvdw1lf8O+1Hk4B0TEY5sYG7MMxbkOn8S8HL1g3z24pDt1aJxKvcn75Ff1sAu33VrVTB
zofXkStRmqmxvkU6BGW6mYNIQ3T0oK3oZfLcSPrxUieCe7Q6ZoA4hDNsSsY5s6WYq552HTS/bVZZ
5ltYSJJh2hCxnnTn4Vkf4+u02nn7L4f3Lia8gGf1WNWwCi0tWT8JdUU9Poc10Pv6W+3qprGy9SPE
pcbnaIB/h9jEJyVXxy6pAc5mtM9X2ju3Hpwx5GbBb+J5mpCc8MGTBb5ujaVCo3a4f3XDdZ83prjb
R1nGKGo0TgZk0lKzJ2e6IjjmT0g8qktwpuLuj3XOzlOOU2QKkDOPkWw5Dk70Lbd5braihEWphcJs
UNarpdIqNJQ/loXk7FImR8BFSbwf9EXslQstrgZr/aZmByRCFnHy/XHjZB+qRqJMT5H16tpDD3vk
EYOegU3Jm3GjzUl7iKYxK81wkXNxu1vE2xCiWRnWFVq+yAc+cYRCO1TTsyzFtKktnodHpbX2Gs/F
U4QKPLsHkO4L/SpqpnG10hwfsJvW/pSOU1wUqEi+/HC86l7VONOvj/YT+23dDo6bZnZE6vZfNRrD
gITIzyOqhYcxsNSIIcj9AoKHVYrtou4bJuIj00z0+pBHqnnPMzBBG4RS2FEAxtmVHlZef9iGgnNB
0HK2JHm06WF/DXX1f+n4ll/dTx/3qgpBMcXvt1/ELygiDGqjW+uetofkrw3W6cOQW4yoJdDVM/lA
tXMDNas8nLwVQl8gyfJMLyLVA6qU0JPOvvREQPCkJMeDbC8B7XzzFsTxDrZeScHzjCQwEioYo365
t/7CEnN9XVRBjpCPj5CWbK/zYQGMzkJDor6Fuhr/qqD/P6xSmK9L4voOV4d+ervG4Z0yas7gv/n9
TShCuv3hiy+qyaNR2Iz/oqMHdLWEsVx26ZYCNnSHHFirJmrQg6mRVlnWAXF7HunDPAtA8E/JNrtY
LmzAnODEu8+5YfzBVtpSsVpGCTHmu8NXSFqVjdBh+TND9+QKt1z3lNc8IETUvnp3lJxEFT1toULm
G6aeCBDWpNXXEg9bpPowxyYA1qMzowvGVxMBmQYF/2Y/jFkNo+AxKB/vq8Eg8UW5/WzOdWgZvFg9
A1IoIDnqJ3kpYqKF8PwqsvSvIzpcWsKh7AQcBu5Zko5/G0c9p9KP+lRLKm2+qJLvUAVszyYpJWj6
kLsELqtfJrMiiQ6KhDLvpJ9OQr1LmQ9RHSTcOMoilIWReEufrZVlMEARtVainhGQjk3xfgIW63xy
M86RsiqFjp2W28VdBmEtxvhhNpM5YC5THH61CYH8C+kZ1kUN4SIkM3tue9ut2H2TPv8dWfV2mpdZ
3qIMEAuWZiCYgdhfpYaPICawotbrP8PqqZSyby61y+jQjnwy7dcV9BlSryhqqM0zlK7nkRRua5/c
ZsbfHTYNBFMRSTyl6wTfafw9fejpW++I4yf4VNNVf3krsKNv79xqNWbGyhlkQh20BRDt+QfY3xFP
Gzm/r+Qc9eG7WpnFFMh/uI+jgqqYHLZJDsgmahPZox+Kgw4ntpgNQ4JiVpjXUhl9FYDkBBkbSjhh
kQ2DF96U94QKXmxutPN8IxfHU1ZA6dtFBw4ZweBhrTnKDKaycPOOoYkMRYFJxDv5kkiiF0zCTvIk
gZwoHxRboNc3/79/tr/EBg9Ys9kIUe7zwp6llpPBwLtvOJtAj1Tmo/m5+Ugnvbdp5mYqyjm/yE41
liOoQ6MRYj7TwXKZfn2uEGguwqhOE/y41rre18EMzcdvFpZ8vy4OTXB+K6DWY4XaOtQBQruWJef+
KpsY+RV5N+m6LJ9cJJL8pDq9ohlLk7/6o275u+DLmIbNty33RViL1vwUCz9wjBJwFRqgTby9eYvr
RLc0R8EKwsijHTIhVQ5Dd4OC/gMxJFeI0HYjDhS3ZI2WxdMWnUUhN46o+H3qPwmMlg9wBN3i6isd
rP1U48ZeRLHtQbRJpOIQNthriT9oBWaDaRUHzhhrPKQpBiJGV1yOxyiHVNp0z30t6lYf9aATxXyX
XZKDw1g4X72mKtLFf2NR/wpGK9HlgOyi53+ZigFVfyqlPnNHcVPO3GK152oZsnTe/bhRk0+henjo
O/9j6dr6eivXG10OmhWL/Cs6KHJ0/cFMoaxJyqyicLPMvPR7j4ddE7bA0QyamWAuU++4EhRakvW+
t4kU6XP1kjlJ4PvcRjoL767pHbzamD78xgwRGAhiDUnLuBaYgqGRDCDJhoGMGoN5vmdfl7RElI9v
dHoZCgMGSmFUkZM2L6yBSKflR9wZp18BarN1WragF3+E3hqnHmARhEBj+a8FuRI2d1t9lNrebrW3
CX37QeNuFqsWTgIVf5td5afvgkhfw1V+L4xc55m4loHwFu0O8Uj4fw9ewIcdsPiQc7K+jbE4c377
eOG8Z48sVsUrwHisAJ10MQ23YqR0cdVcX6ABikKxd1M/4P1cldPz/Fmqi952AGWGPUFr8kJAD0jl
7korfFnCG8mwaF+R4ZcepMOXlUYuM+7lSo+FUZJVddRBEjvgCo3WNXdyK9pmAHM11DRvEdR1yr9p
cdJQJPZ3E4T7FIKMMhLKDVfMZ9rYRVxN/cRlN6N2bhncglYd6TVBFDMvyAQuwCSv0YUpHL4+d9mW
j7JLHmMOC+ekrjeoZKF37X4uhVgM9LkNHBAk6aVTZt76J1RHimYtKfIzf0BtKhCMYqAW/VAMjw0x
2jv0BXt+CvYyt8VG6mZicDnm3XseyUp3duqkFz69VA2P1BymQ9gCr8gNYBo8Z5DlftVk0ccpIEXR
8smzofAeFFwh+evCmh36mVWw/QNRvb4R6fKmF28E4lEc0t2V6wTdxc9fLYoE9XLkJTewoc37hkPJ
JwymZkYAq2bPoEKmuM3skHRDSDHh6FSBpHhgVMGP5uvb27sTvO1JuDlQOEH+n4pzGwu887l+Eg1f
DtF7feCnx9W426aGaAyWxbuvlpFIVy8lm9/pGZBtPJ4vy/FvZmdbBLAoSlU+JtzFAIoV3AJyj8qU
OMYu18JkDjxscvijGUvE9s/MYnW1izsEKbQjByy927WP7ovze2bSt6YTWmi0OU8ZK4MjmC5hqzcE
OoyU9HlF8N/a+M/5eLQCQFCYAfVTHVVNQYLqsxgs6O32BjLDDrGQ4/A7OF2SZfWMjqwQjNHW8RaX
kx0pI2NusicFDJX9mo60euvVdoFeQlqbiBUv+SM6F6QYn28RkoJPiAMfUEQc7gzrFZl7Is8h7lAV
8Kh22WIyctQ1nxM5OCTZz4kMgim0LnCNDtNJertqx8fTzW8zaLRUrC4nILvYJGIea+sgKIgb/gH8
XoR/HNV+7u3fH051CJ0l1IsQBNYXQ/KFxhnQwS4iJKyLQzvJ639RmSYkXJkZtF+n9f23b7HP3r6b
pbIv016XIWQu+wPbY44zLiRQfCiaBufWcaB8Tbbo+/L2eJX2xDCFAGAibpji8CJYAs2QV6SdnQSl
Jpqlitn9hmGdQez+GYGKy3iLw8Y5aZIpZ2zDlS/vGjRb1SQNEUk4Pc9+kqIBcanEPtBD3qvJkkfw
1bVOLXGmw0bXTxfLpQxpFWeVmTYMxoSlxlKeRW2VoG+R6DamsYcykUJ833Ev0PFa25GGw8TC5MQt
ESFhJfY6KefQ9iGb5Ua0i0QXZu5ac58L6eYkh3j4Vrp69s9CYoM8vyG8yKLYYgN4UCM5Wn8CCA9X
d0owBbp7OCk7wadlMielLBcR93LWqyQF3O5GF+ZPYh8DH8SaOojXryw9q1YizPN/jhmDPMWWnr3i
wv2m9cCAGNQt/Lkv83i1/eGQPViPLyw2uGkZSn3Ce5m35Corp5i50oagsmZHPq74ecpbuzdwEZWF
bWkj8LL3i11bWPZK1b/uddM+/jtMeBxmxzbUAGiwvSKQ+pCmmuZnGsq3xuUeIUHlpfY0AXnTh2yC
G+EEnR8mYXsdYkDMpXvsd2dQJGO20DN2/gvuLoRJy+OH6kehcVr302iLcniBjBSeCVMgnkebNwQc
+d8jTLT9WtS1McWj7uSF6pY+qww+5MuFEfa3Foo9/XQsiiP7bRzFYXT+sOMno7SXezqeIDFfX6QG
uL8a/RRDsQp8fctGmki0Ev2LmysLte+InsAMOPuoDqqlHp+aHpXQBwVmtxOAzQqtxBpo8o+2xoiA
BRhv+OoON2r5xqAkSja7DuBTrmPBQV0sqBRNtazvIrIIFrLld9OMYmVXccnpg6QXTqKXVPV3Y38u
whdoUUISRNAn4CH1IdyIKM88bYWb5yUcDS/sh9FaEBKjvb60kpbxqqsSBs0iyEmtGDpL6QyVEVZN
/+CD3HsrC7nBMkKj5gXaIdf+8GboWDs9nrkBGY2DIiXacIz+77cenZdh8nit8vK2uBhGMRPQwT8w
7gfZntqWD8wlwybXsPDVc1hilsSsNnp0Li/7HtlC/M1yE36b5u2WM7lnJRIlj/NgFxyHt4NLNIgZ
rG7mI+UdYPAs9fyXRDToZV2067PzjFNUa5hI8eaYcUPo5nXtCbUgh1aS946x4wqRi7lSuafGTswG
l/r2c4affcu2ZNrJoxwXQ6TGo79s9rW35u6IP28YTa4ul2NKkrUcBMcQ7jcVhEYqi3f8Un5ScVHj
YrjPwoNR5Gt2bAJucG3f4r8J/vLe2j++rw9cqQI8anjYU6y9MlDzWg2VbAsQ2LTHh+2EiONN1gaY
rWzugfHNpNchVPKqq1Oz/OqtJDGVQCXXBN8lYBgYq0+4wlcn1mTS4V7jE8fYqLpqbJQ9vtMCEd7R
+vvNsAu0u7dCLvmQNNKlnanQDczgQxInsQgF0HuEP2cfQZBZp1jA44q7/PyllzLydk47i3Wd2Kf8
aPiPyHP8nUl4tQrOJcqXuqKLzHxdGMV8AS3HX/iZ/9fq9nCGEYAp12TTme4PqWFbmVq9ZgdFEMqL
ZC4SbIxJN/5DQPbku3vso93Cryklk0PNLagt+mjCgtXgDjMDPc40EC+eDMfS3e3eS4U7a/DZXOCS
ywWGJitKbUhhL7cvTvtaByKu5FuhnC4RkYPIESwIb6xO8OCoqWpvEQjTONIEKpfXnoEuzsNe1yzG
VbR6RlfQ90TwHLGhoYKfi4gc2wDGoI+I5jCTGJd6R+BNIqIuSnwyhGoFqcDp+8oe3B2BOgMUiZmx
9QXC4KnxyBTnAahMd6MNr5LmKSB21zGVfvdc8fLyx52P4OLW/2FHHuwNNAhelOggOQvSzxR348+v
FC+LwGh0Z4HgGRrmm9V2S7HaKIdBStC9U+ChkuLP4ZzV5QnuGhLx4zDhHfbrlBL0vSTrt/C+dUp8
h4fuFvEp23zdb/5PFgJEf48BKqN1VtUmljlLUzY8bRU3kvFNtG4CEHoiVRE6nKkvot9a9+HeOpsF
Qk9rSO+mJxMQZVdfoQCtgtPGz/WbjURo1eaC345mLHZkpQ6Khe7oW9bfkbgMhnZQnUMHcr/es32U
r7xj/6wiwoiXY+jiFkojD5rQmPHO/Y9/+vW15oiz0pjsTYr7/CgRARhjA7rIqe72akD92lTCwGCF
08hlo7g5EB+eQV3nfEU+/pc5vcNCyhoP4h3/B2CQJ8E4UJvymXHO3LrKQsoLKVbBctSGj69e5pg/
PUu1goYvjCs2OGFuyZY5e0ezyMfn5VIAjab0JXkY/L8wS/8yseEgfz/KXiQMw5Iz5pM7qQ5xXate
VsVvMkEzE876qyD4JLuqNW/AJvyic4J+1XhNBoFSEmZsG4qf4wCVyVSZEqRY5ZIMz3vVPXHrNuys
FTPqMbIO4kSVTZW2a3WZhzXKsltav84mcNeFaqT964kx4G8ecTun0NhVUcN302hbAWSYsqk8+iU2
OUSwsVlr8NrsUtxXjcMMvBd/QUnd2q6rSvaOKgh0VPMsjeRMAxu8XqjEfLDYq0KTQO0njCiPugv0
KjYZ4WVFuqwDi0vYmSQVaOkdS8zhs/JIuJEniWenB/dR3Jbj/mOzJ/X3hmjMeIqSWtCU7T0fyJ3i
nQn6qsqGC6BS0Yg446RJBswEZs1YyVjM3opU/AbgWaoiwzJIvSQEQbc9b/vBHTHR1CoiWKunM/iD
3fRGg2waUqtNkHsHtc1jVKG8K6hlT5KRpxDII9mQVaBM7tX56VdHxPe4tUyD2o/8McuoPEbUpWdb
4nz/xk4ezqY83dg+V76P0tVpWQe386Gxxp+ub6Rh6ZM3hQCuPxN955dwWt8+go8zpFF9ta5DCcBc
16mCmnYHHMl3DskBfCTRhOK4iP+f2M/m6CGIntC6R98JcoJTVfx9lrcmbJ+k0JXmRor8rhKQCIsw
wdl4wuDkeME7dSLGFY/h/RmlY2Zy3K8/hcA1rfVmXvqgJ9ik3agahDFqW2dX7SQMTQOnbofQrIDM
FYZ//DRvCKkI7Ugq9FC6P+0GH6PQgyhQwrzef/9u6mueIucX0EsEeHH55vCNorGz1gx5wXgQA8BC
2ZmWojfC2N/gQ/msh+giNK65GoR7957e6Bw/IUxhNou7xinPd2sGWAGbPliA1hP6ln8L4g+kgqBT
PmlPPhGbC122gkw2EYxrdZ4Q/BM4eoEQLXAFFtBpLBjRIgvbEgWxWxWtxrXN3/2K1RhmMfjjoz1t
OCkL3DOSYL8CHPmQbKOq5r+K2WRbzebipG1TJf6+Ww2PWBcXZbr/Crp9y6XWd/TeQvpt0oThoD+V
9e3ASgCISsCKICXj7DoWTGsOfDhdKUGy9PXgg18yGFVfSwWfvfybSLZfFFmRntqyMnFAoYJgAsb/
iFO0jsnZ0aCCKAVaE/4vC9J9r0tA+cIS/IrZ+pCdOiIC730RzqvDeDF0R85U/BL7+xlFTJjTe2gs
YVX7IkuZ58S7CKDQajW50aPEHYuEWFCrKPA3c7nQytmlSNJwVDwB62a9i4SYpO0F+41jUHpq0Yec
B02wf0CWv0Q4N1hx/kUTnxNR6GNFnlPFgO0VRqdxB0ghlaf7Ds/e7FlWeGkHtyjBOceI4zfhuBir
H8SSPVA6T1ci7kWnbOTiBDsJiyPYdW852DnRYGaWjOLlE4KSN8AruxPDGs3+sJhTx4CgSauROq3K
D2ZPgBN781yGx43loyIDFJCvNwWCRum47ShDqwROZk2sIr5z4QOZnsLD1kwbNZ6FkNfS7YdwV/ny
BV70v7kqIaFi7QytG93H7vIN9q1+mxr4fC8tQPHPIRNOxiL5mEg6lFsBVMPpBn4jFN4mdrbH0eiK
pfjGDqvD5zoRiZLtOc5icfjWm0mKRcldhl3SXJw74brjTCCQihnXnVvhnkioalYJXhoO6VSJiyaa
bAMw0JwsU0jQMHh3zMRC+O6fsUQRMWd3wSPrYQS0qMsqgrfbQ+sz6Nr2EjYgIQvjamYjOBRzeMLJ
a0UO08wkqqYtdLI5o1pTYsoLnQh+elIuCla2loj9ADs9SEXz0fRPbveoMkE9mLzyUPcUfDpA5VCT
ZCOa7OdA5uCC2HtXKsqpxi1hiA+6+mBkUAADNvbAQBKt5IGhkLXd9xarD9NkpHIXC665ZmPB8TIw
Fx+LJdAt8hO81ICft+r6YP2HxrWz1z1aBwShQD6+WIo1anP0oEklBnqwIo9rciqbzdo1LGCKMcRB
mTwQuD9615NUrSj49fLgk8uukwSAaWa7oX0Ow/vi44ZydMZvVWcvQzOFeXvjDMbt3PzeUL9QGOUs
JnDZSMQJ1gCqDeKDt9rMTDAcSXOo9Ml37C6ib4fIMcJmY3OdtUnjBT5VG7V6W8/Kn9kjODNlDL8T
5O3F7j9ImDuaOm+bM/3jeSjzh48AlBJIW6CBsN6VT+maeHbD7a+PwXJn7g62uY+O/JMvv32G76FB
BxlnvkS5j46dfacpaoH7sl+gM1U4KVxInLy/sMGG9uSUQPR3zzfZETMoRQu3Lx8mbX32YzKK4yQJ
sAJPW7TyMzuaNgwwxL69RMz6vk7wlIs+pqrzlZLQkmhj7B6uUV+lS3CvmWRJZLspesEjW6RU2uuC
WYmLhmXfEEUXPHkn+HuRCWKxV6DnqPfvld7wQYkdxxJ8BAzeNB/VsCYnOsOjrCyZkLAkGo86sQuH
k/F5Ah7YXz7uMI7m0+lB4DJtIhAWzvOpxkEY/ffHEKb6nEEaE8LhACFRf50++Omsbx2RwSBAFb0b
OsPAm3Lnw0qvtO2JcsXnIFYrVQAgtuSzmkTOLHn7MLlMWzFYtmf8u2CS9/SnTbyCBOeoLaR+lCfZ
tK8PZdLGQDZPT5H10G6lBw/E5xaYFI5YGVB4/4loXE8fIaEOxibmPXQFBYdiXojDbNW4Z0PM52YO
NPlHNCD7vZzL8+FeEL7oRYwVFAw9nIpjDYQ2mtFv9Toqgbxg26EOVhV4GMt3EzId/8YHDfcB6xWO
OS9W8B/Q8KUPGSlPvA2Hcknm1u0eq3MyJ+eT9Ry7PFTnUtzhbU+S0ZFF0IFzlvaeUNLRBKNTxJCV
E/vipx3uoQXqatewmPRZQZVw2FECfNMK3pRwf1p796TCwyt0YJTuAqmA3IHBQiK+8/0S9rZThMNg
0cHOVOqfMLX1JFJ3o2aW4nLc7BR7GNEkMtiA+zM3bNeyZccndhUDRYKpabIOeq6BIF0SM7HJodTU
ByBA6D80o0VWuYSK1fF5hHojhgUzjTKiRprBjFJNjp1+hcN1QsxHZGksrkxhDCi/GW24IWf+BS8U
1X6jMJNipHlvoUFILDFza7oxCzDVc9QhyyaB6hujTbW8/wxJeXXpOs4zlQZE52PlRf/HgNqs194i
4ADvWzDvpf6z7aRBl/QHh1wpUqp3TL4n2vrC/6kC7sJjf1ziAKaJL6QbqQ+ufgBm+zMEIaTRRYJ0
CoqasjflGJgbup7RdAjBffIYoDIhYIIWS/18T9y8CvyX/ISH8elnhb2h/e5dgT73I+NoklJV3JF8
4QTd38dJ50yKHDiOzqwTyBISAtBWxjIq+9yrD8dG42JG994FIQkR4u1+UGNFvCavZZ+4JkSyETzm
u96pPRelGyPeEmwm+eRABwre/+UaPJQDmWTnmwRzM/UeApd368EkBf5sLM0vnFtAYAHnJ50Xy0kw
v/RVaYGtJJTxiRmmhZCtaKzBiamDzSaF8pFcoOy394zXethdkDHB14jDZAvZUKX0GNziF+bewsrM
ZUbvai1NxIkpWHJEIQMnVVLluTBMy0VDWXdktqxR2b9XRwb/uOxJ4FkNDjFtFgIAIuNjh0zj4Cst
+tCOA/75YOhy/teDRv7rjFyICeRkPKHsm4owGm5cE+u7UrqW/0IgTHRqMhB57D1QVxlssTb/Y44q
G22n8oKFyofm/5Ap4XZIm3M1mjnOMwfzi55nu8nrQLXv9zkBXBPQ+uw++i/x39I9r6GyYXusEF48
VjgHhHesASDNnXtUGgzCn6/cLL3YL84RTvRnem1WKN3Izu/o01KqfqYdDXBiZ58NP5dSxhRyfbNC
lLTAVwOVOtXgOhJamjZZ4iJjG16li8UnoPhNIg7F0YOXKCjxcCDnKEVhYmVSFMGBJkdYkKdJiLFY
8SbfJth9t2I+dZo8FJ+zLfMScfCqKeSP5bnFNq/M3EV3qyacsH7HpMfNnkCL8JyQe3XR4+MEqVJ3
raWEhhkBWBhM3nq7bPvFuU8+2emtL+TnYAgSgsUozXR1REngTHNkztE/hcfDepSnVX2jKZ10DIiy
5BST1iJ7+WCIbo0VvTx2LA68R78P4F+MIsC5mAcbg1klCde6RenRMmsASR8E5b67Zhv+dp5NxkKA
uBQZnbxZ/FDYIACaWEPBroCdQ7RueYt1bj9mIU4ASIXNXxAy29jAvJM9YFVCdELEFZL3+tA0p+OZ
OZ7kuWczT8gWe3dfdBsiRbSpwE1pDp8HeINhN08DlY3Q9LOWuj2jUwUYQkHKHlLB7YEygmKBK7e6
sytf7gaG+5p53rvGMzPJc5hNyvaGiGAD/gog6xnJeqi7IqzoNUeMrZXAbRXa3NMECZPUyxOiO5bh
2DXPX7IInqnCW0DjW8iFMzRsqf7MChdVrzexjnOBtefMv48OqGXPi4DWnixFOLeU/1paidb6v7U7
gx7o7vXIcKahk8no6Gt/SPyGPFXhC3JuzwcECrZy8HN0sCb1/S55DLxeikynUdb5Wd/Ho4dtZ0FN
N4gu8hroJKIEkJ7w5/hagPxo2lr3Z0L/AgqxK7f5Jwg9bxR+oNVAAlafzj3nXUX87dNfm5GMAcQb
hdVcaP+Th53bJdybf3rP2Hvd0nYtxaAD2z0K7k1lHnPCdgtw/1oJteATlCdKyGn9LlBgBfA+QZxU
JH13KcKbOTdWsB/5jbIbxjjBhVKluLxpdItNypRedJbVmfdySaqHnOcysfInCMNuH29UKghMWe3W
caBTt3WR7P53vLWqu5QuusSfrUr8VEN9kiIAdzuLiXq3zQ+bqEaTtPJqq8YIqJ3KrbJjOk7d52iG
eLn4qpJT+hzRgzM4K7jsjPq7FL2WjTGAljWzufUdER44bN+csX6Y5X2ypZuNHpOXS6jFVXKR+V4D
oViPpEwP4P9qcWAlQwokvFp7+T/HRt/0/shnZUySgTrj8/qQbZSlt/HcDTvPLhOCVw0e4E7mqisg
DjI1MlIhtZ4SsGUk3eRMWifBL8oHeM6i0/sKKGOH7IHzzKx9RPUyXIMc7TQSRIEKIyMj/TNzYyNp
hPlgZbeDoRAVwPlerxVJmGGNN8jfZuSdXI6zOmx5SE+1K1YeAevrK1fGTEo7VpL2VZp5GcaPrCoe
cfJboHA3J8N1bLjAA0Yn/Afp37VYG5Efbjm2QRfZUoRYoSHQGgmH42s4L3cu9FgeS6JXyb6Ccf3F
2SAM4EEICxANLHEBay8sDbhydTkjhu+F9YNjuQtAnkvzZCwIa6js9R0JP1K/CrUnStHLyuhUUzMO
HApCetpSAcwdzrLhnR4zoPRZtDvG6vuY7Dtr2aViAhvdSSGBLZeD3zdggLMjDd7Jf02xidmFf/Lc
trLqvEsL8uGFgj6SgYpeHS/zozlUjNGmYhMfBf4j65Lf66XWwTk/a8UVYKVx2upF14bHNYuB3Yfq
f5YzTLCwUmd+610g/sr6xUo1vFleXhItyKSXYG2MHWjFgzKeD+Of/u/De5QXfhj9iVBkFGqHaipa
T3DZFbhLQewUL8r4F253c1XmezAzcs4ymvJZbaJyCt2zKDWchLPfkdqVZzQaFPHDWkPD70cYKH6x
OVMwJb0tzskVrh5+4DwOpSyhxPkcdNTQQBaxIPNNa/ZcITCVANqVFM/MKu6e74xfBUVjLXyL5CGH
v7rMpjdFUgXzptU3xfOSgc+HftCFU8ul9GlFqazXb62iUIvyjeyk/RZGh/9Cutir0K1nvmWGdKFO
yfMbhm5vBCKi1RUUIbMubqEpuishvOJFLySF16mDlSpm5hLPcjhHgRgwLPgb1xJCX0JbfEANPPHG
16krOSd4Zt0b+gXJi5LhU12FPCpdJRYNS2tLvUB9vZtdqa1+ED3I8tZbX0ZOyjG+WprIas65dBU1
gFbExmf/LPQ9UJ7kWJHbgcWxV5nicoqDbYtkInAKyqQUHmI0gbKCkkHKQAFvqFek7Ya/pAnGU8Wr
c8orkwYBShKI53fgDvfEcw7ix0ev04PpdjQgBJVB1K7KqByqca1TfFWTbgtKK5xRfUJNDOjmz/fB
Ds1YGgW1mpRXXshnTlvV1Hc1zftVX3AkmPBOe7RPmP5FQ6fjcgK28OWTKHYH7Ltu2hPW0eAenLgI
yUgpI4i/lBkxyeZ+dnoD+F82bUauT81dVSJlP0nPqkVUSAVDIaiA2a3NZPltwJbci/v5NquOhDyp
sGllrZTWlj2axu3PlusJKU5w6SghSAeLvrslaIdk+jeNDPEEoa2RbAXDlomecXVUetbZHlDmeGnp
V6fnxK5BAapDCIGhk0L4jiYvp5GB8bg3HoFkyUCzmGLGq2d5ltv8E6d2wcX4KmZZ70ariQdMxZN8
qL4FCSlxcbJZ2HfnaI/U6OuAuJrWcTahWtQg0qjG85ZeQbQHgVeWhijbpzWc28wWiRJ8yJ14oqEh
Pa6mLtkueOhiHa5MVT85LyRxjtmVguobdLDVsvxP9tl/hw7Zal3UM47ZHL5NYyYRZV7dFx+ybpYw
tSA4J7OUGA/F4drPj/U29+PEWHm256b37oPjoK3RYNvbVRutLZ+XhyPSUW+O15d7f1JtiOcEXSkr
IQ8zaaNJLBytfsh8HEkJLlPopFA0ZFZysR05O6KCR41ng7eYgAXW7d6TdVv6nboqquHkcbb4gtCv
BW18gQbiUt50Cr95BbI63z22ytDtd3PdmLeRUbOU+8Ok2N761AlxMgt8YuEGQT/Ltsg9ipyxyF3J
eLH41CirVer1753zxW6438LM3XVKHnqvGsb2ejKWEGx71E1g8zUCemKSoOXK+K82IiQWGX6cDAb2
2IVmXrHaHnUmW+kwf5GBil9kFh8/diKzbBD17exLRLXaUctM4rs2pfGQMEIaY9AJbJk621sl4geV
Trd2IXh65MvCuu+7yAxMKAjvTmQ6oIWus6yroRHGTMazfdjV2Zy2Ly4wxLfw7xT1lZ2OjjdyX/n8
BJEsYZI9yrOu9feXKWkTnJpvl9qHH4KG/px3I68s4tC0JitUULEdfHHMUHHgueohUQN8MOUQrNxa
p8IEQ60oO5chwWRaU2AtIAkrKVdQoK/Vzi+tENlnzZ35iArd4fjHoaSgyLe1AsWpbZsBGgJ+NB3V
GC1r0dmWSSRdxP5UDwgDFW+rOXsBrRzPUlqws/xHgU6N5Is6gwNKM95IdBfWWph8bNEDx4daLK+7
v8MiVxmdyFZHvx/kDo9aQkwMqZchjJ5s/ZPPAoUbFWG7JJWsyoqRobtApEUMj8bZ7STbDfpXYxgu
yUvjaaMq/UB9ZEM7HrOzCzJcL7FHqPVHo1yLvIpnKDglM/i6jaKZgAy/PY+CcC2k9DYVAjZUV4XY
11Td92OWUuWuhOtqALuzxg9jiaSLv4qfwFEdrlFhIAKmY8Ugd7PlA69394OtBVuYnNuzxKv+1OFe
UD5B8iGlYoZPNaWa3hZMFizCncLAzdlwOhVrU6Qz795ZhwoND0as8VVbeUbFmCkB63NpU9eabLC7
SasyC7knRwlkDh/QYzWhEzBApyoNDEZpa4dLu6cF44TQlwp6XX2gcWME5dsICF0VAQU15avq3zcw
9NR6W3XiX653M5ndfSKiglt25nOeWSVuwP8hNlhbnSeizSmaJvMCuRV4WD5rFXVuYl7bos3THr35
KspOU8K6F4sMJ8nndJyntAL3pGJWxJoYzanqbiGSKxo/itzWdacC2NT+RjQ5ZeH+qJVo86Eb/6dx
lqzBXlV/qJcJfwKzgfOkLV0ygt2mlVNmY5wLCd1juSZvUrk22CpMHXyOd/hdfF/imsbqTeTHa+UP
WMx+dbSfPtH+16nP7ydTIXhCcCkmFUb2nR4RzBU8WFsWfD57HkD/3KBSi7yAgQX7e/j3PzG+7Qpz
/0ZJrnJPGRyAEhCJUSMX0eDxRe4eH+P06M2lDKa84Ghlu+AbeDNKNBTI5U9ee75AgK04K0TZM9m/
P6tTG37ncOJSK7zt2+PtpwVQ2HonZ65Ix7J6Nv+6sCymm99lzKUb/PdOzNFiuGENkLCb04bOavUG
CJnOl0qLBhy8OMe30FRPSBmIzGPlC4dBe0sy0esqvsf7aVCESYR6hqwYgz6KTxe6N11clmQiK4+B
Qndb8KoYTTdM9ykuf1Q2GJ94CTeXE8QMfVxci6hBqpVX3u/VMU6Q27AbBAL0z71Q2R8deoUO/fYy
oq5KLCajqQoJDE3xFk9Ou8tDGraLzPvJoPogdR/7CNehYrBrIfzH2mEX7iJVc1z1nb+yqbcxSBgb
U8vdgHyMHKyCB71wAj2vmjguJtZXe0UzONwJP8kEklwCAGaygWcqvU7YSYwSADvTYyGi196jVm4b
7eU9KMFddbsHyL9kf5dpyinQw3qb6L9nDEaWi1hfp9l9WzhusorO2U+pOCzEpJOFlJ16oKWLnAbe
tLLl5VQSjjWuAkgqpa7+5euYbTGqPJfTsyLk8MNjUnkpvogPNqVrN/tLm+oylMFpujf1Lmdz7yWw
6+PZmapiczCywH6CuEnwVyrQH7rmCYgv/Qhxsik/REksDzBYDLkRzaBnholPlrDjIV/KLauMwkHO
fLgx8j8cn2PTZEYCpsxtWuJefrLfy6uBmsSfrCm7ioSSwF1vy+EpfvGGMieh4gwu5doSOclB44SB
8Ly4XDT1cQ9R4vcxM61dUC3ivKeZC65Tlif1+ZxpG6/VBUZditROD1ptXA+E2nlmV/IZxIhaERJ9
dQ+Jp8Q4sUlcDpMarPLoJAJW1pvPhQMmAdHnp6RwpgmIC9XIf/ol6heFJMbzleNOzleDq/YYb0ga
XZquN22gaMbE8+0XGkQOMuj2BoTI+GAcnzkoH0+jPqDYsY7evGH6BMzzLkN6k837YDzBK7nMYlc+
6sVLp8Roz05C3+ff6duQfg1GLZ+MwQ5lVceBgiB4Rm2dnAqumx4LEe6+nerN31+XvO7EsDWHQ9Oy
HK3cDlAsH2XnL8817fUoVSQCBGJ1vNfCpxgkpMO0OV9oVLAoiFoBmx86N2/oN+nsJuM1yHemc4iW
oot2ZzowRdhp4D5bX8id3q029rohOuA8p7N4a0DdM4rsD2ox1ZLoDIYwI96EkwuDiaxSlNlhiDe0
8jwUOZuVr7qng8KI7qLvxM4a547Tf35S8XnUFeFaBNWuh8D2lPmLlkYcIoYB6zYkeKon7agt5ZHC
5o+6yGxvv0uxawQrSWpvsr5pe/hU+ElmqOHNZb2Wlu8sdHFGfDemMGevn55JNHkbI+5TKSqeztz6
5yN7dkimhLnqHangNda+jME2f2D+xKtz2OA7+0m5h2Uvw+GSIqZUQA0ROXUCIExAys64KdUXXQAo
YrnFdg1vIqCxxdke1s59UC0GmXL1pOxw2at86HY4OfCqBksvDQpWra4jWbSaK3Xqg/XxFabuZ49W
NoqDG2FJO73q4Rzjy5aCpyJgiXfU139zwCbgDxVBRgPIlzR5sM5alAFNGdTHrjpgDZWB/iEAMmwx
OFA/KZvjy+J4lYBj7rrlTe2y/WwuyEsee8WI9qgYikxS/32ZP3luTrtrZsF8pV4bMrktXeeAr1QE
MO3t5VMMA5HEGCwFhBr5SGTrU0Zt9WS9w8x8wK6XYaQnGczY99fFIegyL/kN4Snfu1RlSBQ0AMDi
XH8yKTWqVdo8Eg+n7DOdeNNaEG4pyUSCgyDW/QuVwH9gkuZ70Zx6BXgvc09M1ZySvCVaGNU/vSqR
UUU4ydRo7EduHg8lv+l21z43HDKhgLIHrmlDyADX0FPM7hBrxK9AMXZ7Jkm37idMHRnMQiWLU5DR
rp73pmh9rNBxucvAPT3AuNogMJsyvQ7P7fdWUvPZyF2+htPJQWJSAMyvJ4y2AsTrlNlwsGoFDiYb
61G14H8gqzSszCnDX0ZMWslv/JE0dOCyw4bUUOTF6oO6KQMXYyBSXFsUfrtUc1rJbAA5cRoPxWyJ
qpFL5ORVcjPaPHKUv4IEv2Dz2s8SK668ZPMggmeDHKlYcttttUonzm2ISa4+JXiUCOfldGJ954Bm
+zthkxzwwzF9N0DF5epFExPnFgzAkHe8uENyNRIS0TyK2WIUaESYwqnzXrIBTq1vJGnAqA+ZNkbo
NMy8AqIdf0dnk33kPl+u7v6nqoYiOkX0tmAZ7DVt+zmB2Rc5aEiU+D+B4ddUddGqwt23F0eRIx19
OpRVrUXOxOd5skqa2+qEY8GqCTWuzce0d9QPCrtca0WkkmV7prBZi1wmASr7BTc/5LNMYNqfLzpG
+D33MsG6ohI2sye+fXyVnyC0G4fiLT9IOmopo2RYGBpWP104hT/iEzbOxLK88CFqf7FdVmrFV7lF
vSreQ0cEiuWyeN1siI5gxY2owb/h6II53X+ZQKE/dP/8eXYvd+ZKe3xOy1RjgFhvj3/EfMQ3YTAT
2Xy6i8VJTfEYsVqIntZdsES4er2IGv6i3Bfm8gusiR4c4OFnIFgCqPUAMRgR0aAoHS34LiHD6L0q
yT+/oyGRCmyKjcuDU+n87BHiLJwNbz7d2ASjUMF8q312MkkOX3wmTXR62zcmkvFMKu2v7HZ+rIBk
HNjoFuljLMMGAqTwAZS1/tzWhE8o4opAcuVf6OwO1ex0zGSbqsdPnG3fkZBKpJVYUShDpQC3UJTK
AJhx2QUEnwJLA2U6MuIlfWo66qbmA55H/sYANv1XF2+JSqye29ZpsuCpQ0t9u3UDiy9ekvyoKFsI
EAmCCtHW3Fm260/ajEHNlvnNnFdQYIXc2Ml4TTkKif34J92LInMgzenE8sfewKZRRMBJ8Nr0i3lG
7zEHl+AixIFnLu2WfzV2VjvH95Ktb+qTEgf18VBjNfg8bbLhbOsVlpwMjTXx7XbPo3y5ayxBv93c
lUUQ5qAo+d9kaljqeDGKghMWx8MB07GWU8wjUv1wAwB1Am4NPKPVpNpxMHSooMX9EM8rjpZD4Zps
b2abwgy2n95BF9AecE/aA+bDTyNhsETgiQO0pnkc28AZI8lwdCqMuWxs8oc/lilKec/TUB7T7YfE
a1bZ82J5JpNaDFirnFTYk+sNzNFY+fbzcIsEo6TL4dnuLj4JKlYU6858FYlH63fn1UkCuXRRUQZz
GZcNSF7eb1aaBW/L59tFzEJZMgqfQRaaH373tEXshXGPVGleqxFksY2d4gxy/zp3KEVyLbNEmqyM
iAL92imVDEDIMCoMOaZWXhWbiA+RJcHmCwjjG14Ft1ivVyDCoonhtUaK8EfIuhDsmkfQik9gDrGN
bBnM3HdglEp+UQPIobnyOL+prMVkjXxVXMlNwbz6P/vKssBbPb/YdYa2vFad4nVSz7vyuLv8bJ8T
I2qvPraMoEUQM0l389YFM8QTTHzyImMMpA/dS8sBknSP8+25Ja/JQ7CjEp3KfNYYqPS+16XDL80X
/Um0qaxEFgkwWevEG9pgPGnsMbrmoDESC59SP97J0PwUMS+8HXrnTzDDYmisD2ugHq0N1GYfczUm
mcWwUAfCNc7XnrOxHwaqcVR6DGGb52pIbnQpnjPuuqKQdh6qmtDGqmWU3laZf9vTWNbmuAEtv97W
xLHwZbHyDfNBDzFUXKIUOiRIRdX/e6ULQYEWdUG82VmqNIhzJ4Q0Jg3udOTYW6avQjcDUYgnqaAd
rl9MQOcq1NKYRxsjjFEzKD1ZpHG/PFyByhkZA6CeKhtnDj7daenDUS9CE4Ju+F7WyZuq6eWsrSRL
POiM5sNG8if8G9YjwrfLzv8UDUIr3GNBJnakWq2TxyHY+mMNsEAmmscaSceFLEznzbB0eQJkHiXJ
B0XZj+y5JyuTAQx7ZrvOy66StBYR4+GueW8dZfKyCf0EQP7k0ftULX9Z5JKfEHnuBroaOZIFftAk
4a7gLOBlywhPLnUM4c+bUJjth30CFD8L2M1mvoUc7Pn/sJVLq1gEl08eQuY3dB2JviCqIMhMoIPY
C059A0AWbL/cbCC7Mn2iuq+fcKfWDExqOMpadWq4kw5oD1rk2SC9rsnfNOt3iZ9cpp8FQzzOGB9o
NZM214DMS09I4nGUw58J9gwEBR3rz2d+XD53oTlmyH4ejrjIzRbc2+i64AH9Q1vrrSgBWs+jOXoc
eUjFGOk5OSXchFRsd7Ct37weX21A+x44++DwZUucZTaEkynJp/SwfwrwgvN4t0y5mI50xy3tLY1k
rvdm6OPwRcXHw07NAdzfdOMklh3VrDT4YxIlOaF1UBqK2qz3XeWk+xwDMpzyWSGoJYaoYsUg7ooE
ZKbNd/W/Jp2mrYya+zt1kP1zau9M4SIZmZnOdc3T4twiAGeHBse/jpSsK2LdKektOFQPTBcnyteM
6sapggbOrZalpgW/xXV8duSxJqC8/SmVVbGKlqu5hpd353thgxoqwKn9mZCB3mK+Oit0bckIGvqB
NmbfL6JdcE1eA9+4vp3G+Cu0FKo9n+ZkCZ7DazQuUX4XtwsxNpkFsDz4OYEp4Gn8ibAL405bsYK6
QrQGx2JLfnrRkOg9qhpr/m5CmYstsXVstQhsXeTWnmZh2eXtbYUuKQG/4EWTriO+OBGs5S+1jnxL
e6lb9b1NXR0twDobExvnkbWtC1sQ8ooN69znqKhQmGqqSmUbD1YAYC1C01eKVmu3QcPdLsS7wb9H
FCIfI6WeA2Nx3sFC7CFFH/nSz8rwhS63n3EijpNyC2Tkcl7oR4srH98eIM7M7KaFaqVij3tz85eY
G7pcxQLZAJe1wxNHJ1U/acvm/fg6GQS/QYS1m1wJj16RLCz5od4R1ZMyJEy0JkGowL78E6QigvSR
rr2/L8H1/pHqYurDrfEiZvzxqsxFXioDJ2M7Z91I1YfBFawxPa4XctznRM8TRMB9XJKFmwJn4yVz
x5FnSawb571kQhHYE3PRfIGLALhmUj0dTkq0vbR4TqQt1Gvcdb9Adu0EWE7CXdOpNSenAn0FuskN
T88wm0ihU0JyqV0uemJlgWWvmDiApyavkrk3x/QC+ZLJKYyl9VO3YW9REV7BL2BMfSg7xvIVJBe8
lQ7aCpR4ilptiMwlTmkEZ0nVV2Gs5+jlOU+7VrCnJQkUcgXs7iIDqNsUVKr6889e3k1fxQXcXtnb
PnKQns8K+ZYeR2I0mor2JFwoU37YWPU3qzzahqhFuFmPB303CD93+bNduiM4OHoiUZ3WiImZbNws
6zEX6rXdUGeNjma0zPaG7Uxa0N0csCVDQr3R2IijOX+XHG5+2EfE8pD+3yW7dOxJ65U5NBy/FyMS
N5FZV36ht5LiULmp5/6bpxgbQPMxoP5uUlrt7bv5LbBKw3JlmUBZBbXY6l9c2QgDNS6BJfbT27Ih
Xd5qnLotOQY02HPBJuB44YXKMYFLMUF4sgZ1Vmmyk0722RP3gDMzJQmWsUoh0xguiqo6FfkflkKP
2jsKhQ2U/AxcMcOl9uQrTndPM5sThup6/kFOi8QUH85/aZwKJ1228FJDKLMNhUp6HsAjaVepP2HT
OeiriP8G9Gn9mzj922JcPAvEGEzib2YJkxk8pGsn9CKmVWndb4cO9YR5hJXuiLBY02wk5hHrpN3H
PkgzqEGopAGCWEiN1L2nJdZ12/POEYDUxjJimuJc8ICc+CpKhXcxbkuOwTAulMc8KtV3lYCWzP48
XQm/DAWc5fiLoINKjGmVlbVo6bXTkXNCHHVUSst49bX60s4ccuORQ53fHMxFjARvoPEvD3oLpFwP
hAAypiMcnt8B3YpcTIOJyXlrVSecSW7s3kUd3Ur27qGP3K8wxzfH5ZgQPY66M2P0ypaTxHcDKCbl
rU+wFOnj/fIneAoyw3TudtVmJnDtgh/DbusULeyh5wTyWEIG/FJgpnVTLfbAJrPrjdSg5JJBUGbV
18DHT9H+tp6p4Vv3QxceXNPDu8RU7i9eLrWHwnXF9CdzeacMCUGNFu+WrjgpZ8yEz1VjSjiKQwWm
DrLRbZmC5pLHPZ/qVc02vTMTRN09JfL00xj0xJyGN4GoVZ3seDM84yC8jPMZO5nfKtFIJpZcWT4R
OGqIb18hYkugjK3dNt51QADAOUlHfb8WCAO3gvCmZD6y0glVeiq8YsSq1JipPEWTNKgqNqydNXUI
+XaHv2UvL8K5HHHan+PA5KY81+yNuNGVh29sJQitm7xIFCwJ6ncn/HKgJGAqYlAChEbUhZzMlbeS
8EJnOONQ7W2Fz+ZWDz1zkTttDBk3QUB4J6OzBIPocJpKYCXG16pT58VlMn1ZH0egGvKMlJhxivGh
sn2arQh61xC3W2Gv//CCEsBG3LomkBZ/ri2pf0upL2IsGf7h1ZQP5Otw184TsfF2iWmjbcjuM78H
65JsD8XlR/SD5ZGHhcpp5nb8+2zVlhwWxEWrOiFOzuu+LkH7+ja3bgc/Hrly9hoAoYb7ePFVjJtb
TJR83IzH+Htp0bnZmqrc22VkpYBf1YgJkS4GGq+U+9aIQgG6/cdWNE2O7ntnDFYnnNn/gMsq2oLj
yd8RE2ZEaSb911hIYbWDZ2G8HfvQxNXoA/735JX511yB7QQIBis+z8fLoQG7swm7Vt/bzs3GZrhR
NSpnQqbU9TlN0puBF2XEtMHJyBDAQ4CrfJrk9oMMyLl6x4plHCNfKdnU6SwGufcMECY9MQ+Zc4BP
ZqX41lzTZZmRYWMRsb6sjVTZREZhen0C/XsjpfuPy6NgCQsLLurbpshn7N+OyTNBu4YBujo8nRyl
BO/9IzTXF8W7V5ZsfPqmHzU11puGGeuV4aHv3XKVm2w2LiSL3bPXJ5P0J7HacQklS1EKnZUXW1FM
4W/VgppFUTpLRe0ve6gbEkQw+ef0uyIDBmURlVKcvGAFBeg0o2GdmDxQRikjUFK/2vmkz2aQwRgQ
qP9pEV7uzBraZwBN4uYwElgvmC/6NU07lePONAlvWFUUfXWzO6QCQiDJhGQmbicdOIsRURvX1k6D
KCUUwrGxgVlfyIW/N0gO8+aLq3PB5dL163RUajcqemg6S21cwHN95X+6u+zRTJoMhEecEcI9j2X8
JuSfXEM9lBCzpH3ma85EjpRWi/b+xqneSZf2JJAO/2ml2rD3ATlNR2lGlXBilk2fBxvxVuM35fJ2
bZ/a5l0Ohudp6y0e5a4Z9NANGY97RCUDIB8la0qepmT6QJmBBPD0jdRpdxKvIku5fLg4FIQ8bUik
xVyHpXqgfh5PwLAi2i4Ksc0Rd+GZMvqqvYB9cqfPEQ8F4aEutDdyJwKw9spg0mFMGuoAPMjxxY0D
7PIxeqqrqJ6vE3hKyNvq5adIlVxN/kxojJrtwYARcnG8ddCyNwMnCLzANje5AAIJyhJKy+qDFT/S
ZulLmW5CWGChXa/pBtHTLf1zZznXyql1xRjnb0UH4AiT1xzKcqggNMcuCYWcxZZa8uMIL8bua2mU
MCxcb0/kfT7/R8Ioh6BgtopDNKoKr+AmyALFdMa+VjI8ImcvDIkiqh1p+2vj1Vp1AsKWrTkq0d5m
bgRk3mZOWgsCLZqOxp1MPEMRTs6qXs50E5oxB4k1hOAxvDo+BGuz/Sw7c1j5WOY6qzcPV4O94IRY
biAUna1GxhoFbxRfG70X/+X1r6kLDBYAnM3XnUiFbnH0cKd+yu0eFfSSCmXon7pPUlY3H3Lt82zE
+K1u7mJ45LaHSdVERbTqdmeA/4LDYGn2EYqtyq95SExVwBIRXaSNK0fk0rI4IjbhM3yeXB++P4hn
seD/CqVsNAw75J5dj93npufnUZHrMEUErrG+pxU9jH/UQtDOXDK4ozvyAilZcodzU/fUW9p9JsaA
8q35otOWmCaflfB0+YzfjzliNcb95+iuGiE5MgtxJaMBErMTfXU31G37C5PX9/LdQxEdprWSPcRB
ZAKYEPCa+bMvIXpa1T5qXVJr+gH8u2gkeDZ7klBoCskhCVW1y6nXIlmdwCpHTYlLymjoITDlAFHR
V2jb1fEPZgB/G+0UgnrIncJF9xXJHwXQClJZWHu+XMVkP5BEtVZ4I6h0iqPUMpVSzaFh6w4C5HAE
gULULDYAHomWGmXWN6RuH/HKb96czvV/USmMOaZo6j7b0elnwo1E0WDsV+SoDaRKpWHQmKCnAJHk
ObpOFZy4KiMua0lOp57Mgl7e3m54KCX7d5PF4vWrlhVzkwFlGFsjW09Q7+YWVwbE4zvR+3PQdF7q
gRpT8vnPHp3JB1SAZEfBEFN/QXEpXKfrd+jhf97axNgzu8xzCFNol2b7FE78+HOPuFoW+97+WidM
9726298CiP793uB/7CLimMvG82IDi4yYWazEqkiRcCbm/9g/XDsqhIs4ZPSK7wgjLXopgioj9jhq
jFcCmN8iYY73E7dKxCnh1ExkOg3Eq4T41FtF9Z6ki0y3JiD9CgNhj2ZkuSNV5BJIVS0mPYwY/G6t
5ilSniU/X8kUCYdESWXVQdFbqxtc16YQadSuA2y/cenh8lM9Pf74BPpJwtUA11jG1jS5JBUwGgaD
OxoAavXEE0NSjy53QuqftIorZtjwTDzqM+j9v7fmb5BK/L+hGUK/XC26crPJbkCsd/C3oRiUBrMv
P3VN9/XeIYMbpXzIkpbAXatuutGBVs5OhClbqXNMmmqxBQtgvZaKqpVk+ka9udePx1FD+hytvpcd
BTjORWrCRTsQV91jyVnFgUhmCDyETCXys/K0GDUw9mVk/WX06yUD8UikmGnqcuy70MM0+3h3e+0A
WaYaKQB6zNALE0u5A0/7jtn7ta6Vmx586mn3Is4RoYu3SYpO/yzLBtBrZWoGl3N9aVGiSV4vaS+5
iHpXQtvR3jjnlC26+64MDSShl0DJJOtqMudWkrQ24a+59ubXCV1IVYxJpRGPlRMgInk5hCb152z4
BYRJzWi5ctVdhT4u8LiGei6F9tZCdJVm18eRsMhiRaU6Xsr8Ry165L1/KrGq5GPmeENPmIF41jqv
qncINclxJB5yNm+C2sw1BS4Bgee2E3RdwQr1Z64gWnrB0B7VxwWhh8HsPfw489xJZ5jE+Ow1ld5G
uu56E2Fgbo4kHhXqIXO57YnbbMk3QsfV9ur/WUfNJhtrACIJF8b5jgY88DFJrpl1FHn7VH1HAzqI
QLQzuSSM4P8bEj2dMDiKT/1mXISStV4SkPElc0vUs3Kv8iRWGiWrbacIJkRaXt+3dF6j6S0gIHHv
5PnTF5ZHhaq0V+DOOwMQxv8NcTgM2mWihpSSX4mxY5IyE8tGKPpX+DoOdn+u6CBxehTVxZ7bzPHm
fJq2UMZhExr1cUDpNEo+e4GtnhMVKRGT7NFCerVcCMIHK9YuOrvSRNWOVshczcD+64nOuOyrN0Iq
XWQL8d+GNk6N5Sqa7ZloGmBBAWj+MTOpA0aef5SW9tmbdnEZC/yXxZ1hCjFwD2DC/mKIlfcF2+kg
tIaOgM8oL00trJMzk7WZvBruUHCsO3OEsBceI9dvPKDcoVug+9hYq9yvvp54vMHTp0g2jLce+5uM
M6n7MaOGJLwsOBOeqXIOIyurRuCnPJJ/tYN5Ko86bOv0IIHvotZR8SvqoPciBTWRXFeJcuVOekCF
LUi5+FEC3658t25fz9lnZZLf/oAaW+o7lcOvUOas/oGHh5SYxI6Vn3u9VSbm52e2+eXzB0VoWF3r
XfHan+5GakV9dE+sl6PeV6q2EWtxz7+JFgMOjaBaG/c3UJt8aYn7IwsG5f/2aODCP9GwzyPkhBhH
EdU6BT7kLG+ianyjwtNOHrT4U6yHEPQ2MsPSsnTbyPm2TErwJI2bKuJCkH1PQ617mISdsRO6PKsd
yztmo01tD+oImTBHcmltpgLhxgGe4bd1fSGPdazdjhDfq2wNpMq/Dgl6RSCwVCg7hM6dyCR2HX0L
btTyE3eZWzr0MyznHS86y/xrhcr9RaEQNoL7qKqLo8rvDiv56/l46M6b/KSIZLl2BYM9oph1obQX
6u5E84edfNw0+caay3A1qVBgdWTOJzKPgr1W5WvYRhHxHQTMIc8j4ZZjW9mOFbUeIHa0XbpPZ+yk
fD0opKDD+MSiVhDHxPY6PZk2ZwykFX8Fu4sbzZWUBZKS+/Kao2A04uhErzF8o+D88kSLE1oQK/9e
ohhhOU3/9ABOA33Tm5H55V7lu+ublioOQM6bnIYR6Z6ZXwN0/53ie/W3EXMGfGOJpqM2oiaTkpeI
eGQERv12d/ZCFdQqK6Ps4Zjz0sSwqLDIPsfy+uFi09yuTlPK5kGq9t/q2nI5UU6hh2X/J8bNr5I9
MZ+0yWxOLkJRe7cN8rf8a9D+IAoFSVi5S5HVIK/5/fKWeQO5gakQvLaNNuNXcG2QSiU2Fm/budpJ
ealLkKeHzS6baTI43ezkjjBCqAmaVV8sROwmYb/fu8mT8+QopEUgeL2IsnMgGKzjOB/1ooIQobqj
XWKk9ZXh058Qgo/Kw9yuRiX9ulhW3OLpaKn5tzC+j9UVy7isUTdOgcXAf11DpeHA7i9UCPdFEdeC
EqINHvOkLHAIq28a0Y5WlG8ROqcOPyXzhZfuOJwTr9gXzAR6Ipm2l/5nKxZdqYrHSVbf8/t0VxMg
x3RZ5V0HD0qTZD+b7Pa4ksN+t9kgTgff6dKXdlNKN6KR59UoqVXpriM1shavTAIIvjql1QWngLkP
zHVItWCEMN6vYnwr3Uk8njX1FsIv9sx/EG+Z56my4xmewprNJ/AfHO+BaWUU/b5Eg1DR96RKWuyo
XwxOGoSAtFU2R6owt9XXN+ETfez02HS2//s3zsFL2gxBi/oeD44wdGirBq5TLFEEbEZdjFnWACZR
HdEO048674AHfKko0lZcVV2jhbReQP0Rdgqp9Kb21phoQtMXD7AnuBSS8nZmntuTwWHBKnEMCQpb
NGLC7tHNqb+0L8Wxct0V8OlYD/btvIWfp2WpGB/9QAvWa33qjDgsq8imWgTK9T+jHzXLZIwvvJ7A
yOtScgWWmegUKragFaG1qC6/RcOhpBbS9qRMm65G5y5gGstpjZa92aLwkkjoF+0EyYs2epSe/2Fs
lLNZ5wDg25DrcYKP+e6cLMj4Cv/qnk8Nt/40XJDXLmHRLFEKfYULpCMIaLEUH4jLsPFr/iVAzeoH
3WhQjZhdFi/55+C191cPRMI4dswf3r4IxqmDOzBvWh8xkOE1UR9OR8q6BOVvMg8ULYBqfQjGPX3x
49Y+9f4dEtLnaR0A9eLfPcZjVcCT7qny7YZG5q/38PJBY/Oz+fBxhLArtgJJ1v6L0i+Ew3pmc9Mp
TrmsqiMczq4vQI9Uhck+Q0isH6mmdh29RM14ce7VmKRao/RIPTk8fUid7pTDwTQOLF0k3eR3HQxF
NCXIn3wc3xcmslQ1xPQjx1M+0vnLXlCYkzP6yQoD/Jm2UDkKGLbo+0yuxXYDq0VXWmrrUX7x2rcl
iKlOfMn9h+RN6g9Cg5IWzEKGwMKRYg88+b9Entmy2d76BxloN61He9pMmGcX/M0o6Lw+AKfWRNqM
T35fdAHYQTa1lu/domIfvyxpPzBMwYJ700NJsFhKY6NRFIquu+wDpiZVug/jHfXmQNaVkbkFGKXM
oBmdpHgRrBFIQ2fdjKIVHnXKG0XHeGenhpFeE+fFzu6r6u2FB/H3/fu7F0eWI11fUPf9MpIcVmUv
jyWFAr9p1/nmz/LOqC11z0C9PocrVunZgJcqVnJFM3+zo4AhSjrBPfJgqB7Kf7FDYjSuuPWyo98X
tAkY6eUJCHCtVM2hD05PgJIS2t6MvLKiSeXrH0Htr5//f8IV9/YWaFFtt6WWkmPpeITikOr9remh
Jb94Ve+a09590zftGe5vyM2AjJSvb05r2+sMEA8vjvV4pArC81rkEKAChFnuFViWNedJoDmW2uEF
WJhx3di5vftT+moDnJmEhEitGn1Z2DyA4XHxTrjj+gvI5n+8VLrjeBrAD2ot6ad+NoP9byY55jOR
AqAtQPCFi0lQYeRMbceztclqg0VbsFBAuzuRFxHFAgNMBWFyfCcadima9OYjiqpZAMgzQ/FI/j0l
99IsIjgAwgCOA9tfFy3QPV9AkYDxTdc0irHE5osp61UsdIdSoeHXHgtXP2KW8vNI8D4B5jVfwc2B
7XDk8WjPNH/LYB9590uwfEuhvi2FjlqnoLWnj0JD8e3h1Qz29G//CJgNkLyn5rYjLt29Dr6pfSAl
rYQXq/r74mwNc7u/xtJZ3+GYfL9tGxN68aXzeiIKbXGQyOYzJSRRafUEjJZm5st5OQicczeXtUxT
ZylCrJBBov8Sp3k+j8WujFwBjEZQvuTyVMW8LuEd4RZelgds/tHQYrg5UfZml66AWFosr4re/9hI
g3WTNUqdJqSUIBa/AmQnKX2pmnsvIyXkKAMsbnweLpV0qGXuMRAGHdfYqOSa2eqTl706YE1r/tnA
stb2NHWvHSFiouXc1LDSHkAGYkG8ktc6AWOIAsIj3ReDNiUhuuZvtMKI5FYg7V1HHoEcBiZW6eSG
kGtqz1g+6Y8mhpT5+4mmcc/gqKdPaUxLL0mV+u6ZApaH3YFTnNTYN0ChiPB7U5gihBunYXrcd1Wh
BesT4o3Sv90OsV+azfXwYOs6Cp8JtcGAYIA3wb9D+Gnx42yWxnuAVzUD0GE2QP+Xu6JShMQ2PP01
A4IO6C7C4pvJ0BBjFuI05An0uatNzwo30+lHqinsxWGyBqEmzJordt0UW4DMbklUKc3r8kBy1EKh
0bWS4CMQi2sTnTYKgnF0BU0BNIPVaRYHzlhFt0wMs9WVkSgp8aL3iFkQBoqXdxXt0ae+IfW2A7qG
VK13kkkA1N7q4qri96CVXkzxZnWnBRw34l/znsPw3SES9nVgpjL0Evo0TCut72TGs+1hbddabiOM
1umfFHpC/8nrY8hdcHdvXTvSWsbi6egohJN9+Zd1Scmuz3mbBS/WrSF5+XskipUa6yZXGzxqdSZn
bcSZOHcIjO1NHTtoVUccDcnLazIQ1P+HzTfMKH1vF7Q85w3tM+nxMS8rIBe5fcT+py6KobicjAyK
kKfk6olHA4QYJrmClky/G9yB0tPdiTpmfg6p742dwXg0hPwN1ReDfzdiIXutgwaH/6sSza8pwyYU
xrhPhWTmASTxxfN8KNmFdBuSmmFPBla3hfeo4NqzMHIG3532k9avXzSFfxPatUQpojplP2N9Xt3A
5Sd6KZec4JSHxc+TpYU/zeTQWz1bnyzErY7YmhDPMlmQSUWltVT9lWqttY7ap5uqer+/tK/FnG5L
ighZDfE7KPAlOccn+WdKYlV3YNCCbxqMQpZwAppi+j7OKwgIkFvsRTQgVwN2xyg47PmgSdlf0hD5
AFxZshMp0nzIdNOOSiMHIEtsgEza3NUfKf/Oh2oR2B2IJ+zx6aax4AHPtSUDd+jQF9L5xG/wLQ3p
iwgXnJD9kEs2agt9YlX0Ie4eJG/I1LCeVLB98vExyBhJYOAvun6OOI9haSt/d9snUd5kU1pg3Qcd
gVDGaZdR+CC/3k3YfbiVoeAZrBL2cv+RfhEaxD4ypZM76vaihgU056KIj0ajnp3dOO5xNj4B9fcy
Lq89sYx/3Gzg2ls+eUsl+qO7eEHlnp8CQXr+zorVpCTDikvrjwqlFz66o+5/zfFvLvau14mxGhRv
1MA0vPNqRq22VHfbFFp23ma2FhIqnakBkhrNm9IVT9FoAqyptazzKdoag0QO2gUaFF1/BHsEvORd
u2TLP+KUeEIFGSPhd47OEIUxCQOtezo8xgzo6ZsQWrUImvrHf0POWszZab3kEFkIHeeSbYZyKt0E
3WIzlkoT6iVuKyyIiiHAHhBxfAELVnvt18N8VBSi0YnJHvo6arvkHAYpf56PCsNKH6DARkncOI8a
dcjpeJ/qgtVr02L9qR7MXv0o/KLb++10CWsxYEtL0RxlqnYJ2j0I9VUnQKGSrW2N79j1UzH+b8UC
AuUkkI2lxtepO0kfkiQMtdh+pgr9CcEa3jq6hG6Uw655Pq1XsdGFGbHIUZUwCNxe6K/2IzI/1Zu2
4jqVaUSVB7FPWU3gZ8J3fwKLgSttINV+frQ4M5xutqs8QqCuXUm4dw2rwnu4B/Wx8F0PNPyPkMUV
SCINTcgvbUqjqemSgvA67pK4lSRApJ32ZhEGjeKcE3KusLwmsLzpQvcXl3vmLFauum6OYL8AeaN8
+5jpRA7Arx0s+WvfAllwAQhWWhdJjPPzaKByA94RlSsOsEVYgH4fbFgWrD+1r79bwBXtrERm+MvG
ua3q0SbL8ZNM7UnG4ITl5oiYpcfW4hMJfjDEx5Q4eLLomIZJnj8haofsohNJlMbvPCP6f7WjU8BG
BxIKGWpGgPZUSX2d9sZ/q1NyJJ6ofdOC9k5Sb2aNuvdEZOxKPvdN8seWopNafhdQtY0UBvnW/4On
6KAufmqvbVYFd5Gx7i/OrEzwuqUKksy9MQOq7pd8CnStAnmm7enRgihZMBRo2GbQvCHd70N+DTx3
t4nOgj6ixKUMQXBFzbiSbdIy5v5QI4Rl6SpQrnaYxg3K4kBzWeQdZ/E6XaUy654qJm8EtETiAWnA
dJxWWEp+nX2MSpO/zn2DiDeQsdfV0vCjsf+wxbPXnSU9Py9+GqZHGpYMbyeSBcLPuTLVOCZpumd7
F4hEk2qCYtM1AQQaAcOPYbiYBjLkeC0X2oS3M/olKwz5CFRi+x2EUTIJD0wI/04q3RNeEU7pKB6J
EmQEKE6pO9QHk8bNWRSLhd3qeJYfjQ53MK3Uj+tExrPbXHqoOIIl6nUM+e2B3B8OjmSVYuJ0Xbuf
1qymm8699YVsMPbJ7ToVtQgz0jV8aIIBAF2pTLvSkHs1r2ZkxTBoG+ox3LkP20EXADsika6kv2Bt
BZGh+N0fIeXBC23Um6GhROrg1Tj08C+i2R/xA6+KMjvcDKA6p3k479CuiXPPK3j/RKDt88tiqOs4
UwwdFjcwK3bMTxKBc8IBSHqp6Z7DAajmoDuGzej9nn+9jrazakkVm5qz5gDFmTYaRxLNyem+uSwM
7PcmNN2n/vBA8s8R8LTNO/8a+p4jWonW1Ryd1PIQsmCni3EZ+Twb5LeJ/Oz75+CIwRj6LRGZXleX
SFbdYnCvlYYqYHgLX6KOvVMXi6SC/RkMOW32F7C5Zz6g16kabeDwej4TbaoMQpY+3nfjiA72aRvn
o8bOOGumZU7uApFo469yySf6JcpPGp+rh8KmANRm5l9w/R9YM2+ZU12/hDyXrdVbh6b3/X7+K6+J
Ququ0mv5/pAwcqbes1wz6sRFx+3BnTeyIUwwDSmpHJU9vmgCbEj3cDLeoApmi4ofEtom+HJNGFjy
CVWzCXQNYKv00cCgy0R3xWpNHzXIpKEEelxpI5EL4fMBbaDHNap5NK+orvaCFJ7alrvROO3TYcSc
Ec7omkqWx0/PAM/fg2+9wWyg5NjUeALEx2djX7xmAyQQLUQwYtFEJ98TrQT6Zmj203EuqvyUuwzE
6yL4Mwr6YL0D1am8BehSLhTXGqhnw2ndjiaaQ9BsdFx5yptq0uSquWGLIYuP1zlIhzgaas0s3Eb9
HWWAT+HVY09A6TnRDmILztkdH1TUHqwhH1uxPMoeIHMGNxGcbtkF++Ut9juRYO+GsXXsjFwa0Zj8
cO3B/0Ojw+wKMZomOun3cyCRHBkszTEUoIolT/tkAVrIxBmpZkjWem5HU72idVMcey5ZzRgPSo7i
gzE+aFM0mzdFtfg+sajPtLWVgdJMwMsB8gwmFacLzJtJZaVw42I4usypWiWxGD9xoDbmvvxs5X1C
9weFK/nyj3pw5mBHswYygzhCx8cwuGOoP00h7HkjyGWTQ4Zx9zl+hAGQgqtwdatC19bmBDzONvDS
ADNvHgkYrwcbEAfisM8j45yMdYXQi/gba9CUZBDQdlZbHmZdDCXfxb/hBFVTQc+/Dkf2EOj9bKDV
KVHpHI1yodYLlKr4dlqtZR7+GCJ42HHeDgMlwi0jL1Yc+gdqoYtVM0usdenpZaYmAa39XJIUClxl
SExfmz/vqliMg6ftZQ9TwHE5IwXz785/yByqIcrYckich7GPdQ3V/mrfeAl07akgycWD4D16U75l
spP6DT0ecVGpXv9IUnq6r0WTc7tUQgIxWszbOyio04WDrcuNV+EUZcxBAgTwZkPkRDvK2JRMfpo7
oUf6TU9ODrMiOfdm7UidYLUHva9p2QlusDdXB78SO++/eANWlaiwwnTtKx2Z7Blzhnw1TxziwreM
ZYF6Wd3wvg4mFeARfM0T2uqYerlV3/PGSOwxpFXHedGionaPFSaU6W6HEh8ng+KMgiHZhJPIvGY2
TGKNUFqSxMZbBftyTlJkReU1I6wBlu7gO6JU10shiSckT++tpaeUM5TTnXKIprF729asAANd5KC9
yxdYyZjp4wrZpuWoVOiVnDQg0hscOdvWVv3mFEvPirN5+zbsbfGna2z/yqO6+Yl7ytEr+hiyiHf/
CXCyHFcDc6WQn7MNhB3RIATRU8aNf0L9qm41HgPHFGlku5CHkIkly7uOP7jeeJ9ziWbLPjM9fSjA
hGRLQNpxB/o0rFVLJA2yyX5+PTtO0cIKGFjDfxq8MlVtxu4qVcIoLyAz1yXB5za8L81wxMI5JthV
SoDbFKe4t7em0S89eRI0nwgrLOcenMigFjEbUk110evapINyUaNPwYguhq6kzFEjyQcGREfp/lvB
JJmcEk0mQssx+qHGIxBIuJNdy49ZRAZTmyhNpvWXwqfRtppt3SsPhmQJH0kRGidyNV+gYTPYs6wG
thQY835nnj+WRS0gt37NlbYJeVgaRi+ivC4x1PQVT8S+yN5dSh+MvbW2nuTRBFvzUgaVs/98aJ8R
NH2EgNZIjce/5AkoGG8NZBQDcfs3wxmtQ30GKOEFK+D31Gorct+8ATl4MzBp08fC3LY3HXGBsHAw
kQndgxYDpiBtI1qOFSYXjS89Yl5oxBUrDYta1XPfDXKBUARV13jMfNZMoiqU8zfAtU8T5BjdyWvY
VKEhFx+VUy8rYLVXLnTDJgdr8rDkdVffElpumJqDL/1PY9oR+aO7r25tjLK+fsOdnSmZpp0kZvaC
HlhxvY3W0/itieMTV6kH+6P5NmCws1YxdaVgFjjo8e0kf6x4IBUCoPmwVrBr56duxK7b55uheUck
zrku/Qxx37ZOz3EuYgq6zP8pe1JF3XyJojisO8WtyC+1du8C3chMdtAm7X0iICp6pq/hpjsPJSiN
ooPzVTDo47Zs4O3URqNWwHvMATcnwaUdP0XLTygrsH/jk9Y1QMhqgeDFjQB2rmKXEBaxZwxjz9pn
5lxw57GO2EBXaGIo7FaAvEcL1JcAGKvP+qUB7q1vKmih5ddvjpltdtzv40Y58nrHZHSo7+Pg6bM0
5vuRX8eyecVmD/g33qbXhPHfXCRGC3a8Nm3K+7iGhZI1ozImnTtox/lxOvSJTblcKcoQboUKixZd
u8HwN1nrKZopTvgf9p4BpEPuO3GgLI0St3x0H3Ozooslkd68knnj4chD5nRLCI0sW9a1W5jU6ZQk
xsxpmewegrsoFFAGlYsLfubSgyKP/rJDv3QscXPthh5fmbyOqIA4PUPbAuUEgazK/2FCH2/e2Sag
YLgd7EbnmnP/xlJQUTA52pUBdxiz3edOGWQjttZpj0LU36zy/9/MT+4T4ybbyQfoBQ0zsPInE0nt
Q1gCEgUuc6Etb4g4hGc8wGBlRyLn6VcMDNGjShidTJ6azLOK7djI0ERmG1sI2nX3oNhdoEdnhVLq
H8mMVSA/g62m5sg6nHWzfIxC2bohrIgXycYeGRdICDU+mtGuTRr1EnKdV/OnVdYMnimLLnfsukyK
97pn3WLC4V8qnwcJ4xLnXRYqwOJQBXHk8Ngcqp5M7RVYciKJf2olZyxkQTC8Lhe78KYVbCUeWEkb
1/JQmoqlLv7pbZSrFTBuDpQI3DcLqgObXq2WEYODIvFnWf8uygAlMwT2g7E8aybJxxIN/mOPBI+/
Zw+sPFrRYTmEvNecvufFQlcFUbTbkecaSf6WSmiwqvRkSQWm7k87kk4ZQY3r0+tWLlcaQotG7wkH
xuMBeM1bDNtuej/6e8AQsbXHowMWUSNHV/oOIQBXO/AFUWObl9u87QsOJVaUOIW3j12XC+HmFeRN
41724LGkeEi5XdQGJyIdsUyi1dyCRZZqQxZrjmnSp2OkLTQubmhwpQjRYIK5Q54Ysgw+zscSJk4B
J+1+nuV2yPFeyyu1At1BiJUnaDj9QAB8YeIobX/0CKqJ9PorYaTgkuDTXgaM89pzWwaOfw8SLZ1w
lsXiyfJlZ+5liQW1vQqvBaZntgs19u/QQW7Oo3offK7FFY0j7OW3cDxUcohAq4ISizsjbBmyh+tE
o4bm5DeA5tf7EMk/6LyFWZSSV+WzhD5bdjkzYqn5hf7ITxmcYmmOX3PyljQAPSXTLrMtqPBj4dYT
eRMNQPoxUdwT3KmV9eOZO7WFuQe7b8e5e33T2zLdpLCc8KzcilJcX8A5zlAlDDA+5PfF74qNZz4b
5GhhU+GFyFQZkTgNpw032tdQnJ/g7pjRq3NaRROGjEDrHOj2pxg9chn44mRlHaenEEEG+HPigMi3
K3JjHoCLeAsajKXlCtpVrzvsvEBAN6duyrkVDXliHyZ7zixJwUkpOg6woa0NPBGWrC4zTqeDv8I7
jIyGFasCmUt8A95vWkcmXqs2M/xSpNl4Tmm1ThGHzR7Egl+MzLFKNVqGlcgU6t2TG33G7rvb60nt
JFFnntj8Gl5ry5ZSaR35lOpPMGec9h0T5Y2sCKym6zYou9fmko9sJ6SPy1VjsI27F+IRO2kVBQdM
c36ocJQvE0PuzxiObZMI03lbinU/AXaZ1scmkhTFEAopIBo1lhSZYCHboxE5kwHAKe3gf0V2Ttcw
NG0KrgrHV3LN/4ZDVSyaWTSXILZCW4l+lYfkCGI8BSi/rng0byqnJnUzWi7OosYsdnwAdaF5bP0H
jntSvCRRwtMGcu6R5n6hLlyBrB9UonVOU9MCXhfkwo2++VmQO8At3321j0YiJov7oeuAswRBqO1k
Z8KjsgkbBVXwUqTq+G9fcxTDGJwjyzH3PC6eByN11399hmOlSV8g4XPabUNRrvNL5pKm1QpPI5bn
ii3J0OA1mv8CXEKmQbXl/GOB3qQoyJoKuEEIQYv9143zWpks4DQHq1tTCMOYmePJtpyR4cUSjZui
pxJiuiEApGSgvFWWlMtAAbh5pD1AQGkEHXf0/mJV7V+xLCE7xYZppk0x8aMPCv4XAG3yCg0eP3qP
WLrjIgXel2ZU77xInxIeiF9TH8bNj43gPaSPgc86Sem2QH3JrYBOnxNio4ncj2uIUCPkM+BT1WB+
tHv4ObutqvoU8lesArKkpNnaQm+9cEKiKglj+oapzghNtWUZoJ+JqvPmd2hAyOmy1GoTGpw2nckE
z6wb5mIMNlk/6IOFWBiFMOhAkMnA3B8j0W0KUpADwQsPmI45kL+480QO7qKdjSIohUQ86d0Ntxlu
QA20cYZzlgarICO7vol/LT4MHqrFEhO008YQ6qaETs1Rk1XDL9Iln1KmZ2JKAeU8rz0Q6Pewk1Yt
QY/Y3m0poLlZgIFFrTHuIA7s7vP6nhv0meY9p8W6CYGvV1JLE4YyPNb5+hnM77zyA2cmAQXGP1bS
AEYtL1IenRmRm2nQEVMQ8eTdlznkU5lCu8LQVvKds9nvn1/slRQecun90GnyEtWmPev8mu5nu7kV
2kcjmWjUN/xIGXTsgIHeN6ywSyNlxicMAtUE0gg9kIldB208/nOUaX4GRktIPTfuG5O24rcIoT3a
pzCXoi+CcznNZtY4qwL6EOPRMRWjluf6fJSnL3G0dz8l4+nhyiECP7sp1R+A1KMkoSaRofGFcp6n
FgVd4g/BAhjVgtuuPfmxnZ9QvhoXOSLMb0uscTHy973MmEqfH3WyeDqKN1iN9SgSB7FwfkXYF9k0
auW7HdsyhbsLVBANdfb7JriF+vFqZTs84L8qgsJm1McfbIsDKp7WYzJGszwmuDuhvm/IlZZ1y45s
OdfE3tqM5xUjzcad+nAYB+ej3NpfJZXLFGG9Ms1QmXj9GJR1Ll1l+xrCQXkK3HhhO/a6pmDiqcS2
2LtvRiVCAqyOP2NQR8jNf3wBGnKiFWJrFAcWVaYV3Hi8flyJg75HkZs2K47WRCcqQ5ZSZh5+JOye
cB19JzQ0czjihJJ+wv8OurEmV5FMLeYSokfHK/23iRggx0V5LOcgNiqIkCuoysdjgOZTQIDnIDbJ
0pu6vg9DfwNyEqdkiA3p0SyQHEyaj+a+bvWB+6CfIk1b+bEb1+VdbsNDckx8oZC7jb+HUUvbfsyD
6W3RieB7qeTagAOGijKXxo3Ksy8itwRA+RTHV3a3O2gWurOjnMOc6NLn3t4auVxZxgn/6rWq84NH
EnHcDviiwxBy907jbPOet5NSaPWlEFTITCYtGgGNSiIQjtbAPGeK/CIDGdY/ONHzBvXGAz3g+QHF
ACHQ0LYOjrkSqH/zGLXvZz69GbYmIaEAINPQf3NlapjhYCelZOx21ZWqUcZudw827KN0l/2oo483
WHdVmGnhE0xQX/75zGMYCO6DMbtOy7Z4jjT4pYmc7302n+bI1dzDyKAeStmGulHKau/czca+ssQe
BHABys/k1VbE/smoGGAnk39gV8FzoKCaDqNQec0rqV+Qk7lbceA0/uFCNlOE5+6R6z7nWw8bQ3Lv
jyZCJzMq6GFeD7Ye1kDmr+Xwft1a+t8gFaCZ+RFvc57Jfnw7KKL7SNEjW+pNZrlBuH5qwxto9EmM
fOLrRz1GVsl6APOCyGZJYh0M/e31RBGTslfaejxiPadBQNOt3Jdvp1So0WNnxjsPFTeOnjDK9mgf
byDHRXA0qjw8h3ePg0EjqqHxmfX2O1CV9YsPhYtJ9Pd38ntDgO2MeJsmrnylK5SwJpKpRhhpNX1Q
6iGh1bSugLPQa50u7+kPXhYcAQ1qYojKTZBNovytf4pWmq9gHO33spCtU7teGeJ3V76RGiREhE2i
s7XC9s2nxzzTi2KbyBTBTJZVsMo3ViDKJ8Mmx0VYNEofwBvGMUTSIwwm3eh5Z8aVat9zdq3zhDJ0
ou7lvAxX6V/d0WAfPaaTq+wWuc9W47kvwtUcdjEdKJNj7KrZ7XSwY4SH37rc0SDujX4RRrqjGg8F
UGNBDrtViY5GkEKgVsVXO1Ssa4vEHpRqMChzHPLlpSKFjfIc1Ntb88959OeawlQb9YHfcYgYMFKA
IM8UVdM4rql01/lRRI1EBBfOaVoBL82iJ7M1YymZb7BbpJdaB9JfsyKTIz331Vuuwkf/Hr4j2v7W
amwLrusoNYi/qB85KjhLTtL/84q+IE9C90D357AToVvBfVaA8nL/Y5MavbbMWTCOn5zpkBmL5Or+
K1nw1WytsWPJEj6YPqek8l5Ff5gs42U8+E5/Ye6GzK5a+XnH2SoH+g/OK7s00TgvLEcEFbFrceNM
0c18DDEBz1Gibz++O0asJHhPwf0HeNOI6z8x+If/+7a1bYPXoX7+rUPRODY72k+7AWqO2sJhDR1s
crCgkeecGCPYwtXW4HDlbb8NhS/Y/O5gxJv8YDosqDfkUSQmrrAUKHCrFzN7ERo9HMNUvt5CBff7
i7yDsN0lpipMFAgdHS76jVO2b0qT15ClQZx8ClqnAwho09T9XDDlL6tN/UsW4OaEyTJgIGnAr49/
REMm/9Qg4LZPOzt6PkaD8i2XvsbRly9kaPk0UZeo9FCC/Vcwm9gL1iIk+YNFTnQDdNcPOk3Zm/ng
F3cLAriwoTqLpOSstMzBZl7F1jNMqSeoqoyJUXvqkTbFV+f6XlqoBYMyAgmrfajc5N2x8wsb28qZ
krfsOLN49wmmoJIep73QZj9XIwnw1ixqABtKxb65idFIWO/MTWh4fQ+LF5jekhLdxm+SFWQUhX5X
ajOpiY6vvWuZX3wmXLQfiXe4V89dOfucUrz6n2rJ5nbe70m0XPnRV8rJNvggpMCvLF73TLRr3X6c
Ole6KeOtMLWHOxJ4Gj9xnLCL+476Ex84DDGWIklP3fBMsSxki4CC1M1tRjwiBxciq/EIbL/j2KVt
J3jtgvQSjOBMuTXpv7UghlTP65SwdcOY+6N3UIGWzxwBX/KWkadxcoPMubeT9fhdwTRAgluH5/MG
kKZeyZ5PPWRMOUhJzVRQzhSwYqmu2gzshtiJ5CZlIg/slc/3WczQl+66Q03ARcKWqQOJv281nElp
v0deA8k8X4k/QW0tSDWZzEJoK96Qm2hnJ8IGfRofNR7uDxEWDgMbu3rFrCR0OXbCB9H/IKcR5c62
w5znbOv/zDk2/ZQjz8hC4Uyoje7nOVfhrjMZcduQxuKIUbMnPDmt9RmrqHhlHWwKVS9e7p4+g20I
ZUSgV/lqHYBNtBqjOyE6R6BtJ6HYVqDkXHkMnKQSTpxq2jVeJZ4W+qoTHb6WbPmR6xPwxcuwaVi+
CoD/++vYJumeII3uTJVIEOxOXYGkRlG4N3APZdsEvvx2XW7J6bWfeJJJozgUKxJrMzXVSPjvE7RD
GNhQrEB5ThPuOCyyHmmn4GCYZZ5sN2vivOWnkTROVwxW8Cwkg5cNYCfgOfQ7LipPbYjNKuM16+Hn
uxubCGiTytLdrdEuapX8dUTbJWxF5Ll3KSpgMnLg7hH2AUcXz8zXCbHd3a2guVtqOrlntKWPdCKz
xhc5zRnobGEtucIYhbGvBu4myZ0kjGrzFDfm0XIv0J3uU/PBvx4fib5jU5ea4rcW/v837k8ZtXx2
KLPvI0bsJp3I8ebSB/+7I6LdmCKmuyyRjfsifCBySuCq3Y7HKUDK5MeXP9t7aHAnfJLvT/PM43b4
26cGbPCPJTLWokQePTm+aX6j5rDjVMAKSL1USiMslOZe+HDN+4qg9UnvfLmR/nAiSj9dYSszwAYf
+KhG4jkSpU5Jnrj6AGg5JC5IDT2hwRR1+p4LB2vvMXQTeXOXIVKFFVXnQyvkLAErv9/clmgi8krV
56A2aBaZSmTqxY4cRd4NwLCMXxEumht7O4h5MMH016P+IfAa16zb4tG174Pp6CLMnfvATDk+LnYT
IA8WgH9HGcFC+w2DL40HwWNSx8Cct+mOADksdKHQHaa2YKb0N/VcOM7CNZgrnTCxxEYIcYKVed8X
SgvL5qEDyiLKa1BJ/tRpbx8lZq2Q3iRXgt5Y08kbsa5ArWdg7vf6ftlc+N94AQchVijr2OOq//3r
+oND632fCEmm9OKXljQXzYwgYHjribiR7EjISJquEEk754SxLbdVmGqLOrgjfkJ/gOJNzXZiXq1z
HtutTnKLxOg7U0m6Dz+/AxfXGx2sC27JrYXp0a9uO49f798btKCYaJjaopdoL60HXSmbPweXbJw9
bPhotKY/CbsyFqv1fvsd8dX/rPJTz/TTmWziaHAyLJY9pRwhxE88Qe86izla+dfqRwkqaRB9unlf
PM8V3FCLlyr+cB/NeSySR3pt5s3J0hLwvKQrQVcrEMPz26TbgAX0Be48MKHrLLkb5Xuj+kl/Re25
C027W563Rr6D1zXCXZecNvtnHXLnah+ndt8PQAXDukGqX+2ZLfibWqxk11A0cBLPMvDZG4MA2Qqt
282lr6N9EtwkT6CTfm3qHHZfhd3xTc3h5o18FWHmQzyZcQe2AG4PGD3ehVwZA+x1v5z+zm+F1Jrt
ZZkCgPq+gwVjAmhytwagPdJC0BDOxLoLndr6Z2UoHaeHPAmGVACaF9vChUddNtQmF3kYw6yx9Yri
aja63R0MtGNVstFBsJOKgbveTyndVvFgY7fmP7/Udj4qbf+aYAggnP+H+juEP5xR01AeuBTKbAbS
T2oDyYUPVzSDIt/3W772yRhCTb8JuAUvGgPYu2YhwA/i670FRZnV5MiGhsDOMY3htq4ucqtSRaVL
lX3VWGgyIq8rFLAPZwg42NrCpbZrolNYkyBlMtL4mCh3qZYd59dDnNaxQzw2OW5WtXtfrFUWEUHy
X6jVNFsnBe2p8YrrvHuwDIrLn9wj3u7SIxNIAdN8dIqd63BYYYFISNDsl4k6PwoS8jFuLxchfRZj
G5+/ByyaUNGuqqC9g8ew1njnqY6pgf1zggepK0/sOTSy2O64Xqhc1hCI3ZpsJlMGHpkV+DMcFGJ9
2KvAMeFxA5fmEnyansoBhiXofT5mNdRebrxWVhZUeDMcz1iuDfaoa5k7ho4gw63/M5oQSlpqX+1m
a6Aga7l6W4fK0ypjZIGg9FryO9w0wbkTTeCKb6GOnwiJ40NMRcbH0UzUImItdRNc2CWr0tz5OX/t
LwW3n32JOqmyT/w5c4OkzqviMxT/fWFlDEHzg3JaVg0o5AB367RRok5H7lykApBR9y+/8sWOYyfn
4cjy5m/HFo+TeFAB6MDhZ1NoNdCjbj4J1+66CAw78/ivWu5s9uGsiaQLA93EoBKRG27A2gTpQbKw
P+JDfWTeDjBPsDGdDGR55GXaf4kNzLXI6fQsASkQLDKyaFIbs2h0N0MJ2yytWEzxoJyB4RjALoK0
TVCjfjDKyAwRWyIAyYr5jyJ+qw/4U+r5O56He1tTQvkavWCFCEN39vRsv/ialNd0A+eoECKiOevn
9s5hvQRPp8ufGP7RJFd9qGVIPnAxUDjas5BA+TlcxFFHjp+OgAXZQkfkvKcgjAi+zXxw09dKEtho
B87iLx+dnq3+hRiH89HOBxHM6BM3CPz0i/SQS34a1hTigV2o9XRg0Qjqn06nvmShZeaOWjSQkGjC
98ZqCRVcXctfKw5Kx1lIrAa7doiKJAaQu+kofHz336LqRBTmh0tIwzz6pS4h3DaPdje2Xlj+9NO1
kxbusLhHq4K98nUwb/KfUgiNamNfTYneVtqUVXQ9V++OkOFB3bIGaT8I71be8IcE+ikKynwAzAsJ
uvuVYYt0blFbtYAON5rdkTM4WDA/oxohdEzBPomWP5CogY8KG+om8DXCMNGBtcpAL635Hi33Rkbv
PJ1rOvFoyCUCTQNuOszbFv1FjuAXRHEsHhdL7MfCjALbFfUaqauzmD9UN2/mtmw46/xx7SaO1CQ8
YYNiiyV2HrTSpJ/QWlTAeEXr9HB5iEZZL5pO18ixLjR9NkLVlKp0RblWMsCt/eqlWcXHNO9yf2/E
gRQVtQFlWXU9A7VX3nuZhIU/5d7FB1g74I4NWCWVUviVf/SfvUPmsdtA+Beim0WlaccAeE4KvC0D
LzyQmYxAG1NhSBI/OalTMG+AiZUXBjNNZ2GWRuYdMdsq9DsgNZGBHFweImKHbzsYJvbO1LEWecqy
nj7v+BwMnMqBzWJNuRA/cJvQWfwPxeQlapExuKP+JFUONCOhgiBh2joQs/aD2jVYgL+GW8bDy30g
QzoCpi36JIQoG4RT92RcyUmkxQnlQix72nGJc3/4LNCugePKM0JOMH/iLySxPJhTMu742vaSGaZy
sJ9oakSOh7lR66lG2nBftwbbbhV4X7CNQCGOArWcJGqWK1qyicP1BxF7dnFtUzot/y87c1u2cg7e
nNfk1TVg68JJQPKQ1aAik0/o6qU9Ux0v4eYjinGEFJvWjZGYnfAiibZSiZh86h/osM3+kNXwluos
+q5ZEwHgjh7E+VmsmWQHTX1UlP7Qo2hC1X4pTr+hpfpRClpXxR63DzbJNLnGZ4CXJqZzLrAGjQuB
xs95MIft4V1MvJgHamvOIfiswxTa0qCR9/RC3EqmU8dkpHJTgokEDUlZRQNOCcpWkEaVsXDZB48S
6mmJWiipm9QXhWrSjiQ3MtwPcpcrN7FMoAwa+dIRPceEb8nZGLy9vWQF0X1zk+jZjHO64BMIQJo9
RkYzUW/rK54RutsL2JXCRFSANG9fPkQI9e0i0JimPAVAwbW21ze33yumrq+BdvKQ28iuHZvB4SGr
YYF10GCFNQ+MSxNTPItHJ0L6p4fGel4/rPxbIAMVn2nYyL+2X/Be6OEs3Y5MnunBr1JmjidekwLE
uyjS3fWF67xlw20lyGSjb6SxBrK4JqNwLDPk868WLGqV2wOQsW1G/X9aU4dOcRnIm75sUwTut5pZ
0VyTIntllnJ5PiovkhA0c/4lRRGpYThTuBPz7wBwpdZ9kYj9eKJIgWsFxSwn5BloXAs679ibJtqm
KKsA4PzMHzCZBNFRV/jjKeS2eOG4uytSZcXGS08lMP0T2TluiLqGTClo/cn9USqDU7r2xnty3wxr
1HHWmPTo0arT92mqSQft2IcVkiEcxMKIY1TXwmcZm/DosKNSGpjvQ5xJWLnJnofzgxSp6XVVqFNo
e6aTMIkU1pQ1IHsdFGbUjkQgM/4QICKHktsyCoODGirNlbo6xmnyemfFj8DuclnM5+ncWo2guqz6
4JWi65O+QnmlDhxk2D8IAZCLdjzXmilvYgyZetYc4ZvA6cL9VrtuiFP5mSvChvBz5ZCBHDTeiScG
W6b6TIlurNgtnT1WjVgufs3mL1WNo+rca/kvx1Q5LZHmNZZBA5nFbwwGZ8k6DzvGwZfNjFeJFAca
N3z5mPOdb2hzxVubuG6qn0A85j+qIiK2HhYz+n85IkxPedzSDB7I0WAVP6IlPcL3YVoQlc2ZZZ8h
KHGSZo4iG3lfS7Enf0j49EykkLFGEweWldVF1YNGBPJg+JsznZ8oC4RSVOi2X/69YSQPKZ4Y3592
4dDlO8jwbnf6Et5w3mlq9E9Ace6t3xzHyJLLVk8h8cVz+P2kKoUUYaW8ajlrvQhy383gzZ5zzTSK
fnDZWuqCaqcZzlM2+/bGq93JPQTMtwn0N2vnB4fNU0jneYadxw8uYuOUZoNfcmBhlQx9EInct8pF
9jTY2kghhn6m5HfdMdtCsdyig51UzUE3DeQ+3u//f2PBbmy1sjcvv+JlkuYKR+ox6y3ozy57mP8I
TKhaVyojR9CmFwSmy35YmOsicTM8b6Djz5agjoMZuV9BJ1FYdlt3KTzCqdMewhXYj7S2qJ+wS049
MkQJUiLXbNfGA7Fg5RTF7pbvLRG2pbnb7fD6qmmK6dOOOpq+edRQuiWpHTf86JnQ8RsKUFHfPdwq
A2zIpnTlyas+MoyNcB9GmY/d2UkX/pQm0ieLv5PTXGl/SY5iqs2eg51p4MztuGWbZX0AvXMbBHKM
drW0q05cHn4z7tqBoyzuG11hbtwIO5FZxlZHJcG+ifstYrigaq118m3YlPQzVX+aHfuoNmPj2DIn
Er8MQcD8XCdqtdzntgieDwseTt340Xo01xGdWp1rwC2CsbndQw4d6eMwJacNNc6CBoIjxVdYVK6m
Jxtu3DPhXeioxr2i/kn3HRZfUK57sa1umleLaNgDLSbcf1xY3A95je0jUGyVDr/JnsbXFUKDwTv6
yg02BtllauYCrYryWNa0T+ouQrunOSokvjBxfeGf4QEzGiiMm/a0reXDqN4cfzDlVwxmoqVgts11
YXPrLuCdlUgx1mqoCMK99osFot07wUP79Z0uyjY9zGdWLAXC99dDTTqCRqvGN2RRdZ6qT5EGgFPK
QU688rjtNDqRGr74b9fYI2MJd7WbrYdnrni2bVqCty2x+0Trq9NXJX2KbvzA4Ou0aY369e0ESCpT
6wkcBknaLkkY07Jnf97kNoPjQcBagpIHlvp8xRoNm/og+eNOL32Jhk0RlGpCBbSomk9KBtBYzIjf
3FNSBdbN8d24a6XorvEJxB5npsVwC46otcw49eTm7Cpzl53wmF6nxNIne/vNql4W8JJlm1b4FWRj
Nt0jGwliVIyBhxQfGrHTd4VZsyAw2czU/3o8+0p+0U9CysLyWsI3HLWoD1Sbw2Q7yef9MABlqAqe
nwRYqLXQv2WmSLFeTH92T09D5Llch1m1JARlNO1nM9mdp9Q4UN6avEujDp48dNnyRp2tENSgyaJY
32WH5cCskauaPrNLlXGdG6yDTPpfHLtlstKg6198w86TMBM36Y7EC2l/J4IJPKaTgPlxsFfJUBW9
fhoEvixXt3s/Lg1wRwoxDsMNZtxxaS2jlcRkj3zeh1tHZsUPlSV1pRKdDhuk1e5PMlb7tiz5SkE2
UX6SvIYqL2sdTuXmFt5m/+Dq2YvM+94g8SL/LrHBG6jDMAgRnxPWbbafY0bub02ukl07qM/o7umM
kHzoYHvN4mll/i6hEr5Qh+yuKoPWYCJgjXkAN1DRxd3JXpjTwMUey5ump12wvQBH3outFMuMlsVg
PDW2rsuOM9WYeYzUMjlGZz7lLr33FBESmLFUZsIp70J5knQAmEwUP8cJ7tedjZdnqsBZveCKUiJw
ESEoc311yNBoQA7Fv00zTfOBboG1KgYP1VckSyI1l2dDSwVvpnCHWGwCbLSguO33la8ZqdRGHkA3
qTs7vmDJBjuz4V+Pi+6BUcfINE+A0vF7mbgAj6n7EyJRtn7i6jk3Nv70MEtKnVI30vqifbKGX4mI
tE5l6ey6xI/KKWSsLj5YjExdAdBcjBYJV3nYksqR9x7V4AzjmMP9J/Gb9PhhZjichKWG3yi1ObxQ
mBZP6FAjXVv+eQtM1urcpk0AVLlABK9/kcmzxfnz5i/FqKFGT9X4ejXZVLMvPauBpl5uVv7e/DQl
gfySCgOYCmDO+Ze1VSyG0olTkyx7cGUtennV9DdiLXP5Ugg3T89zl7onur/bdQPMxlTCASPe7Hlh
60pWPxyEAyarMCnUCBsCoc219syMJhuE4tQ1S5Y/GSRjItZ0x76c+OTr0A7Hu2NmAzf031MKfdSE
hBF112NDV5IgK0z14Vnve972vTw2v2qMWAmmey0bjUqlgNZOKFJg34p6D6QxRT+akI4VSXWuhc1d
sGSmgEodvHbQULnE+8ZWI5uCU89YdbH+Ho8Qw1nTu5klbQSIX4XpqlLK8bc6j07fvSUYiJD45HYT
eOvdSF01JuFg4Yr7YymmPidIkc8PCS2CRTfm/E3F1ZlX2YUIAMAGytiFzilfFAIepIgq/Q+GH8jE
2zqcH3Pg1MxyMKzkiv/6I4VfAbgxcTV7NAnYk2/b2QO84VWEjzDfMUhpIPJJQHGDUFBW0VrCau90
ZnPzQzvRQxZWeqihLrPUEriS22rAA5uB6n3SMIEolIHKk0QO3d9lPMgmGeLaVS70COH7PipSXlQp
eVXbSxXnlYDe4EZNFz/nnYP0gSvgNmJ/ph++QpTjYSLPLiVitsaf8emfgG1LUgdQTW1J1Z1TkFf1
jT7QttmFISqL9mOAwr5mazxGcuxux9cONuS2b1rNfguoqcxrivf5irJ6CcBeSpPa4w72ABskt4Wp
lKE4y4aSlxl3q+9mYgBTmdf2gIsyvLG2zXwJ3kRDiXZgo7jAN2XyNRbIFoBq3CAacNrp2xzASo+q
Pbo/NnDH50UOSXBkUP+DqPd74v+bF+u3rwxb90gqxPgWqvsbFlzYsnvnn2luSklv/Cbux2bS5Iqp
j6Px2BhnuMgXmmeuQm2TbWsnvHEwELjyuiwFjGjnnL53o9Nw33yzgd4doN/qL7+xOHlubz7EF5wi
QHz+qA+1+ttqjSHaM9mAdkWFu9TCOAOXoaHHEh59EEO8jUowwS05fOyAgOnKXb169Xt1okFBMoHZ
+sMHu1ONPkJkZIaGLRShsVzENchaVUOXIjGEDbnT/c0+VY+w8iz2IO/4x5xZLprTLX6zjoBRY2Uk
GCpx+NTAdY5lSFDC/ux1ShdHja4RtsiaeAC5k62QPF10AZiVpQL/Q6WR4Kz2waFYsRU+vxjkzcIB
Mdx0x5Tsg2ldxo0e43lPvlfh9+RQVw86geyNJfDF/j8Wcr3HmcP3OlsJNi17EnFIzwzHfhd7/hLN
NZEdcebtkA2uH6uL/mby/Mpy02bNrccOrtjEnA6bLP3tEDQKDbU4tfeIIsDiINWgx562KaHANO2o
gbZpkg/RRJMub+5jkQq3/uY3iPR5TxJx1R5H+FR2URuJrdVLCr8mz/y3m0sEvS30wHRBc+Ynm0si
PvcbqlBSlZb2daY7L/rfs2nUUfbSrfBAFq9tuzGL8fU0h5Hz8GX3erKejVjKK9ZQpkzTnPFHVHfR
mOOJ6M/N2fgOrlbIHVNd+RVEkGNHU9xDeEOYegtGUrbhZKVXs8WDD57kZUmmNO+xVKusLzpVmmJb
EcVD03gnL/0HEGIkWlvJB8jFu5hLFPaqTLE8ttYg9HWlx4LnpOZpStC7KWdp3yHwlhlTmtsSSBTJ
tyVoJbu2x2Yr+2yVbdInhtf9TE6ZuUXhADdxP/7VSmaQwvubCZuxg1kArEfA7sGOz4LXBoFmo5AM
HIRFx/wLEbqi1fK8N5gsX0JhAxiYsqpbgYcN+fYb+2grboDz3Y/knbiJ0rmevrP1jRnrqPbgU03X
YyAe3NBNyLRdJyxY/xNYQYNshXjNC0MMuVLDQ+Q4vaiM2WxUy6p7hKrnDtKPWjS5s3TLkzVnL+9E
yPZe30fI8BKcIBMmGoOxcsGJYLS/iC2IWfJ2nyKlh4KdNak85PPAWxfoUSfWrDqcPv0MLZFiW7wL
T2k4wAg6bTnyTIHZMe+XksA1xb/Ri92LHr+kAh9zBUsQspPw8Ki2YyWPUhCuWuwyV8iQ+bK7JMS/
srivW6WCxC49dc9nBEMH6rv07vRjo4pXcNAtv8HiHQCwsHMbJjTy2WE3XrgIx8qjcnYStaAESW0+
auMyOHw3LAl+1Oaaf2V+Ql2p6mWbwB431Kem2Nem9O3bqLw/PYsU/Frd0FJdGzvbDU88TSUndjOV
MqvXTVgRL/CSC84MDKZvDLjZAHmnY7rRwwe2u8aqKc3risBPgqeJ7+zMEZEH/gWVVrWvGAlIa6yE
BGndrw/vLnq52Nf9aNn4Zs41+7SS3rmgZev0Lo7IGn3bL4guemlB7dtxH4weN724hrLH19xvawZ/
VRiJ2X4T2VVsiviYCa/ATMkev4OPj2sOIKyp62uVdJa/v4ru3ksD5tmzNFj2mjuPFunuJL2lLlTb
2/q12bSb6hQJ55CvimaX1g3BAXy4ang8QTkaZoSjxQwW31rr/lB00SXLfv9f2YICI3QXrVEDqVC3
QqDDqr18/4g5bL7gDoaUHBoQLhSd1c3N1djJRuQ2vx11MYuDiI9q2Em/E72arb58nnXJFMjcx8Af
yuEXHL1G2/ZZKdUedOUnzRJqPIyxDSHTqPcJw1apUo5owJTSgxc8yWzHAdG4Vp9YLpT/oXS0YqZ1
mGPPGClxbrMRUJzH+m5xiPA7LE2VAV7ZNJN5xZoNgeAhVOF/ffQWGQX6bi232+GOfb4ecZR1EDk9
8pAFpLblDpWlibyrBU4QsdpM5z3pjeUsJpNnJJftBFH0tUlTEGxnX3IgGUupuK2caafVhs3EoQs8
DJZsXEqO5zH1dW0NVXhe3wmcZzralLsQiEQJ4jQ+p2jZsK3qxJsz937t3bf9N7iAQF+ftZHRxOiJ
gi1vg2XeaFvIbJCOQH10c4F06aHwqvaci0nRxQDi4Vt3Gjp4SaVwKHrrr1KIaMGSQQPWQBkh0SlD
mUpp6q2MlG/DrRHIRPz6s4W8X/kMN8/VZu2//g2MVei8g8Sz74gmspiWcyk+R6QUEPWJ6z9VeFJt
M952a2f60yuDLTyI+bqH/HooweFAI9Ub2CKzFHhLa9TQgTk/thvGDBSI3pAZ+G2Bf5nz3G0dY/Gp
idwtySMjlvKQGZ5eUp4IzqhHBSQ5NQvsq2D/5eWeXfs7PXPuRrcaLayr732fSRr95O1xXb/HTRYA
EBQ/BW4BEMsMZeFWjXdpByAwLzfNCzNPg9a3M6Fzn3VuSi0lXJV6bOFDBDpukNNzQQ6iOiziUFgy
XgO8PtTieo42cEnWDM0j8fhvdqR4ZRfIAbmHtliV/Vt6vPLwkD7KWWvdVY+8sY7rPN+niodlwnzb
jgmvxJQLEQ5+RINPkwNgZsWwQXK2/dHNsNdTDtMxtTTcEEnQW0vim/QJPwj0SSj3NYUoj+pBJ3b7
ulSPWuJXS5rj7p+f7A7tIAU7TV7YzV59JIg2vrT+C0PDQA544De5OUwHLxvWkE3ZnEWT0D3XuTf9
dRlOezcvS98m+bRBiG6nYKZGNd334aC/B9UwxpDpO1FTwLdUQRGVWvJcorV8lHPLjuj4hmrWwPnb
OynqiyRp1OYTXWMEhXLGZGQe3Cb9eUq6Q9nEeeSOKUbrrGkVnzmJAaenJ7OUGt90pyszQQyQQwG2
aeMJSPPfylaoBNJXLk7+/BG0GXUJ8I1O4cFTxEsC9PdhqrA62hbKkXKWixxgW/F3ggN2zR/jz4LY
G05FqXeEQmfcrcTw16kMJJSLnPwhpiUZyhMv8+8x9mHS/Fem092qNKpu711SOflq+TxyXVt+0wpH
WZ8nyG9pY12vySr8l7w4QFW6z45XpTCu73t0aocjvtfY8oPthdGbt9PixtEltXJIgB1o7IflOQH8
TVzAu2F2M3SiC9HqqrloQp4TGQqIi1oDOuwEGbrPDi+L2RRi79kBVlukZ1Y2Eq08daae3GHmRaOb
tOYgnXV7GSdahKTe0ZrFCxZMXcKpWcqqVY+UygX31LpPkszmADFbJirGaPo5IKgYg8Z28pzI8tu6
QnYUeuPyDbA9ZvTPeeE5usLrGSHs06OuFiQWlgZEvOHx0ZVhUaA4eG6CMSFb2pgCzJVSS6G1Pa3j
3cgusGzcZV4og4aumxb1/RooTjJ+eXnEOyokAanHFIXm3uY4QAKGqWQGdASJiTd7snQ+JEnHeWdV
uRwAYIqEl+siq0r8ZKg0SWo72a0JBtfBvtQnzvW+opBDBTbKKcVc6dlqcQPmGbYYFxSeqFD6ISff
lzF/trPU3LK6xCx08AVcQ6DC/7edomdpJcZ6DrfogKB+OCP/bIE8DmukbN6Sln0uLHcC36IpVJ5s
KiSOB9TYjOmd3bbPnYm1kIJhmtxvhXpingVtdfI4qN7/p9SaAUQJcLdkSjLcIIaLdjC27IXCpw6V
+y9RViY5nqbxbV7ZuL8HbXuQOyudDZiHhF1RtBRk8d3bm+tShSkXwj/zO8lo3Wo4Ssu9mA0llgP/
ggyAlQsLb5r99zhYBDyUpHl4yZ0gzz2g6CFdJzUjYeqNMk0h8Evgwt2Lzf1ylaFdIAGQTtY07u1q
Kh1jCaawLRYup30Z9egaw939zL7IOEE97c0qILriw4TgYpqto2pSOpRtJ/qEWGrskVS1EWpSTZB7
l6RzwrN0rb+ZR8DIcAstZFfxJW7ZETvgu9TQgGIuJq760Ar5/dplqrC3MJt5mB6EwemxjCag65bL
TSd8+cEJ9Vo1Qc9Oq5gJRPdAoW8petirgo9tvbB8p8m3PjyUAK+EU7K2GuJbStBx3TZdmxpc7z7f
h8MkPJrCsxdQwDR2GjsH3SlXg2nV5GBtQ5dpngrnkOqLkR7pRAyyVrRjeeNIbCBKgWeuBy5QwKeC
xZbGm3nnrUmEP9f4q32/T/d7tUhxs92uP0RZ8EweICz4BZ+dfh8yI8Zo9XNAXVufM6R1sh4oSGVC
38MT7C9qD9od9oNyPwfqcRPM+sjAJ6Y33M2ji/pNIDMDNjijs2YBbIwbUL4jWle5va89tBryL+bE
Ub5IGcB2KXL7Q0ttB7m+1p91w2ZXXUTFWatCIaD87vWBqpjUbFa3ELhDYfQX1N3OkG7c1nKOGitR
cDhfg2TpyBHpHTqnSXY87cUYqzp/YZCGtAsf7fsolbwYJtwko7iB//JsDaPm3yo8LoMoIpKZSoW8
HmFjVGxXOhGVWCuyF6UIgkFXaEX00LkRpe9e0mq88gAW4TM0XzGzQ8tjIBbtwelujRHUVfKUMUtY
UHf4VYS25JxS3iY4Wxv372/prj6fWheI1DgkeXoELX3bxxCgCIkmKXltABE7le8zDhH67izwpj6l
7T10dG7hhYoLEq6HyifeCW8VhltByrsk8HP/TI8NNK3oNM20m6YkxCGPYQIL8bFx9DxioJuHUa0A
NppBMKbIyycARiJUyqPwQwcifvCacuVt4AuNco6t2sWHX91s2yBAqQNTk3X9qr1F+seNP1JjnW7a
oW1ihJtyDv3fTEPr6LY9Z9Sxm5GMQb0Jwx1aYWL651m0RNImiD2GvA32iQfYQb+0Co0KSkcxaEb7
K+PC5gNtBRHj2/vBQ5dpCIPT5eCG03rkVrksNxwLGCj2yT6wf4mMNbslSaokugWoiwFA4x1pCqhW
ggQ0RO5GJxvmsdCZq+k2hgpWL7IHSCjBok0Rq+eiA1N02MiZy0OUxTF33BYc14PciIdkp+MwhJAT
jLS0czd95UcU0Pab9u5Gnf6F43iEHqDf84fN55YWuo9Q/25EUxp2doLwk0o50jO7KLnPgtHE9T/e
24MR/69hj5DJ4wTrqf7sUNElLV76suhhivXFBkaMy32oOTFjy4xIAssYLVuiJx19ido64xLZ9zp1
bNhbOmJqNqYRUe9a/Ttb3gAd6TIXqEGUMMvEk55l6PfDAvuRqjU2aHothsXDUoO9fJaUGQAPij+A
Rbewil2BSPtXO9adBmzzFHPCKLJxwwGPJlsfYxAmbh0ewX8v3ixYx8d05eNWHyPVI1qM8ZP+VVTE
CzRmc+ovJPzkgDO8NoUFEuIP/kUJe1Hi47wYQ8eJPSOiMF72gO0FU3vC1WEiJekfLSIrGAn0x/ke
WqpNVLaWzZB8sysviugigLah35lUlsclA0cFTaDw5I94oEa3dlUH5jYaqX93tLa4lDhzf8B/+qY/
senL6056Da/dUUAHmFPZRSPI3+jqZzeg+J90VERwpgD8mur1dFA1sw3tbJzw5/JOj3G3ov9KOirb
mDecap2OTa2njncMiXOP+szUAJkmH6piBbA2n4EQbhng9HSvZCOTw9meht7HVErIIQh9FeubYNK/
S6qWod4zrQnEhAtUW+YebcL8TQM34ltkGvAU9+FGHgzIMeoilQKNS1uBq01NbCVnek6Rh6l7z5IF
hvUa8fcJ3dc3rf8AMVNvVZCCQHV1yYWV+k3Zy04qRR/xsR7NZHwf+Ua8ylIHsVvTWERqCxq9zODa
1R2nLF7QIv/XFCLPmja8t57PeDrHROTbf13Bo/9BMO9EQ0oUNyP6PFRh5ecu8Dj+Obc5lPbQxYzQ
EelIrbTvN+tAWWjaeR4Z9LTS3L59wObd2pRehffDgq0UZYK9EiuiuoCQ8lcK8/gkOcld8IoBsZw8
6yEw4fSdUOSGjxddMouZkWEMMMNoCf4PZZpcwRflS2yt1mpkriVfGHK/cgFqhD5x07KE4hpqtqh9
TPN7Wo47GD+CuaqoQAffmJheHk3R7h29aPGMUCGF70/iR0qoxWo3z1xIE1htg+wlSXb99/ZObkuF
55WIh0o66/dLrUg3qFyTmhSIKj5kkAUFgrbLBXOwQ1XhBi1OuCSnup1UY90qJGYZL+RNpNsuIb6c
ypJP7CfM/kheZwR42ebPEdti0kmM73cJtC84dATKVEmlKcoZEb3iQaK68aDcCR7Or/Nw2fwYxse8
hwJa6cM9LwI2qmELTvXrrsCheI0e0AUTP6b4KHpLoR5fGb7CMxtMlO4M7xqWO6WxERkj5kcyVT0o
/gr5IkE1wzazdS+fsf1UHjLgREE84+esz56JA/04i7eWSARFRzM4SYSXDXDyuW1tK9pLbS0No0Y/
ydbtikwjWsjuWzKttdmc1bU0u5nTVlzZEnzA4dr96sLPH7aDt09/tvRxi4mEkVTIxkxAJRjANP5m
czc+rXYotUJYmurQxZJhZCX5gwU/ql8Mfllh6ikhZDwELTrcdRL5vQ9KjkUb7g3tEvJjw04eUT1G
XVuwIBBbgHOngWnrOiNwL6K+/axg+M/lAcpKhK63zq5LX1wXva0PsOs7pMJKiPobkZJ19MxA51Yr
avL6XSakP+opk3KA7sMoSb/YUxiEhTLzlATs4/bIzepB91ZU7yua3GJUioOb+MAWhHzW7kJcGtar
PCmgfMcL7WReO62EnicMJc6btTM7jlpt72+ejXxNksGUSIjIDl/RLc5WOJu6xnOOHmLZHya3BsTZ
2iBHOmwN2M04q8klrj7u9rmlkrSV6I4P+u3/XIypT7OH3xsWvAWQyqs70LUP6chyoDnB9lTXy6Gj
d0tAe+Sz+18kJAiY48gyHFhoSM9DIFV97SjCk3NQnbCWUH3Y0Kfj1RBqlAwOGjZgmzxP/rfObMUY
4X4aR/XGm0mUW7x6vO/f0lL4FwImbJDIqeQ2hTv5rR6ARTZnJ5zaFwL8vhnqfMeyPudDPORv4t0s
UrAs+C5e3n5ulzcjhAgdBfYODY/WC2GDeX/wJsm9u6qdWp64vg82nSmBZ4C4uy+6Lz48dm1g+XO+
uy/mJVQPYjQBpXPIyy021G45+lvZrx/JYS37e0kuNTRPl5/x46vEgyqqkgegTIFe+3eYwaIRbzkd
KMLUNsaYGj6gz0FrT8zmmhqBk3kWdrXi2o8bsOHG1PFXNrOpCGh/tERj2NGKRlfUFM0Y5yznGL5i
uDDerJd/YG05BYcwl/x9tU5Z8bCQNTbfKVg9NHsHx/liBuocqfrsJDENT9dvjXHsxrIheN5jXViY
Wwff4LxfjR5gEwr6kW7Xx8EKxHUoD5b8cxP396vMt4s64xlZh/m/eKaVibH2xGBUzMwGeWrYmxjB
vtBED9zf86+k7fghlqe5xQqbCIiI2god6FYSe6LapeX+2P7fXg31fBMph8dlJGsMPwTIieH7fgVQ
Lf7V9S0Bru/9zKRZezx+cMCaKx8N/1u+I4RbmmW3e9svxWNvoiljZJWo7VY/reh4QWYGmxStR+BH
jRF7NaMoWmo8kb4Gf8nxbnrpoQTy2OVOINWaaGNdpz1aohEL4V8z0oL2iVge86qyUZ9C00AS78O9
xAcRAWbRm/Q4eJd3U93sQGwq5NWGHQPvcXH8jdnmMdG7Exd8w8MiaY8lYU+FtQY+UeD4mL9Q9Iwd
U2FjnvIML0tmENtdhEvfCyJBRmtMQlgyFn8nqjEM5g8krDis/RPSINMJTDPKGvA6pHjoRS4Z93NU
Pe4DbRwe8dVhoQ8Fe7W8U/xjXQCEVNIADzJhST9AVUUW5GL21ww/MpZv7ftwLtkgLfANiVn8nJoW
GUe8xXD9z+6lpnHTerK8+6vGHxru4+e8Lu/lu7x+vxsxvbFEkQBanNKddiVfaaa1kiRCbRQOk102
QcjndLoguFayVSLY10Ya6V8cnIV1BK1dE743xskIGQGuafYLloYcVeXAA9padw7y7qWQMBsj+11h
GixjHIhigC10KDd9tnFxISitR1dKem6ZZggctiopqIFJXuqOf/xzbFEo9j6i6yGSPqyx3snCeiOa
w6ZLEO5JRIvtUnIUqNP6iTsWPsKU5uoaEBZfpRPsgVLOB3oveOUk5zfjuNjxshauj8c9ZNNF+RKh
dMhxc1t3N3fBk6TlRkUE8T2+ok2lOPU2ZvRZN8mU8Pnb7laymWLbsRxrYMBEFV5MXVQNuQlNuY90
Af5EApFgjgn/xYIJUhTI2wo24XSS6t66Oenlt9wZqrkjRQg1cbdPNlp5mK+RmCeE+rcljrEk6FUp
/MINMkj8p1HGjXkgLs3pdPLzHTvdaaCBYjA+3GgyixqC52lonsdnR5hGt1M+83GsigPio6JMyWYM
kuTb1aVUftVjKw0ABrJkJvlaFjPC9eHZoX7EKjbVhOD9qS4X19gRHwU3HeOphE21qM5JV5z0NHrJ
BBmcRouKztjQQSW557NcBtQtp6QLWolxGz81cq066GZECGh3+MPRzTI2nIF5tjYryMmcTcYw3GDn
vnzXpBhqjQig9/tl0O5ZEPdISI2tNe+KdSISfkSajRC7A62BeOboLFj7bWn7kiZOvNwnlsRIEfB/
+Gzrn81sjP9jOHSXrUTlW891aa1AdlPUR0iqayHm3gg1zfqtKMrZM4EKKRaCpdWWOF9BWRBnOoYi
6xHyGONY5g3/FX5zQRKx0+2VWHC/QTRg8KrffANngwi7UJnHc/m7LUp1i5A36bNyX3vsk8Hq5uLr
kGoCmlDurnDiPEYGzdCD79ifA9GOWFr6Id0rp/c+PrJWuIhHjxAGf2GxLDideMvgTImLsCjFuOzG
H+onY9QPC4y0sNrFlKnSHcXzMv6LHgWLK8kWWEktAqwd0Re9iYmO91a93UUrMCB4NHCEXJhUtu/V
xd0FIiUiswxOzamYBKmaYp8zJ3jAkhoHwtHdZ1fqoZQkdip8vJ3b8aYqmmnj8F88KElIQ8XdapFT
Smscq+FNfRqx+2SaYj+qIpVaG8AcKTfplo7PVRaxAPAmJ6CSDyY3YHW0lwVDdXGzYGiRZezkYYBj
9XbvgeriuJvs/+bdBlLw5At66c15d7aFx4Zv2ys0vslagybNhq2Jl+L4m6HA/m2l+QxQXqhgKXUY
2hrLh28NrbwgzYMC3nBZLc+/Cl+Jpi4hWFM6tAhlXb13+BKtn/LzutxyiKmFxIWFjdzm1MCkM3jy
H8pQDr9BNaFDeOzSemQLMrdAoCNRE+afP6MUz/gCbrnsPObB4N1nVo/kCpmcE/mk3BELb6zfPDHB
PAWRpqizSd/l7PVG6tx7PXMQDge2b/AFhAiT/WH2mVxWAaiOlAJW+VuqBCLIO6rg9dFa7ZHNFWHY
nwjDeQ6paRpp28T1CAMVmOhDhb6cRCl/j+H5opf9t6b2evQuHHJ5zJzkFdhWC0Q2uT5fen5OkJJu
32kexTohPcebsR5ZobbuOfainNKnOZfmJnXpk/eh3qik4uvB695yapkayv3tJAlMWKL5kWxiskIH
EfVVEjjAqlCGUw36o1fZ+1gvtRIPhRu3wazi3lCW3hbOg+rveTUPtMW5xVkh+IbdKHOh1+nrRxfG
gy0AFyYHurg2WL4OwpS/GnPfn4Uz2fxuIAzzaPpdtiFrQDEAfh5kBIRgmJzNhew6v9veDtiNYn3X
EKzbkNGWpfFZfDjZGiKU5lgSUYNftIk1ZYMHEfD8fe3iOjysfLkg+Kjvt4s0qjuS9KYylfQCuNns
v0ekWMWulHwJ1bU6fDipwCujZAZVrD7xzFs4Vr3c2NEfIpwv6yKkw6qb3UM9i1PG6IGUO5Y+G6eh
TLpbIepA+H3//JNypQYh2QL2dlvSzZAjs1od73anj6us515NfTew3fJN5wmIcmAvAAxN50jFl2aD
i1rVT6g72gux3GAJLllwc2HjyCx+RtYpQbpjYekWVm7WQB7f3SmmELKUjFNL0CaH4D9Zrx3V+PXZ
Ri3j/yjx/vb3ZXVZ2/Z1kVvnaneXvRhawj0qbbvpo51mZxGAhlLWbAfNaVYcwCzjs8PeiGGRGxtr
0fij2WqRQ3S8cNrST2+AoPDK5vISnRThA/gehfPKYQqNIOIRBwWCYZoGq7xbsirrgSlMqILS60Cy
kf2w/PSAaTyPcQPeIY/5wrXx84JBmXwPpOeH1WkEs5RpMR4XCpL1p91C67KWosD5cZ//+aVtGIQt
CQYPJ1Q961Db+9HiI9XcIJeWK5/zIpByNoIgjKClC50izInr8MK2jopF5QZiODOPNGCZksW+m384
vTZa8HPkycjDUlaWD9gptVAZZfRRDE+yK9wPbBeE5vzy+gA8jdNxYCqoqen9mZ4kB37AY5dWiYKv
4Cv6jupJWykjxsKasONd+UsZwaldD8CPGrQwmsc/mXAx7JvLU1ZIZnvsprmSq2WP8PiaDzfDYEyr
+i/qjJ8NKibmR/fk34Wv9gz5hZYOW3b6OzATpSwQIKdXOP47ZM/60fU8nRVb5+MOfvwgpP4USRtc
6gTl+QIX3ipkNZFtOxXyZNjdIjRpSw533/jubrHjjfsP8OaGXGnAQNbTctlBLyeZEa7ZD5yg8cK2
Bc0KjIhjIzET0axsw/sETg7x/wTaHU/mbRP7bqmlNHgebx4jVjJNE9Yeq1bLZRM2j/hjzKYQDKca
B7pr/CYKtJCeYSPWeElVn71O8fWiXGjXwv2z2kdg4L29xftGFgcdAjIVVVC03Def7MzMMcIdlMwi
DYiGTgwgD40Y2U/Z1qOY5ekbddgyn1A6UKA5g/dUjUQnz3bLQkdlvzkRtkYUooTZzhonADT531Wa
z7WbeEe+s+Eqs4liTgMpJ76oSatnLK6FmYOVLtFqgj4UED++pCJwKg++NECHa63e4wpd+Uamg8Q9
ptTbaDvNCbMjkK8K0J85HkTIejmtuxV6ZRiFIWgqBpUWTaJptPgxac+K0PlyCD4QfxwsnE4jmJ86
E1ji2njDia1grq5UnCUlGj+8PokpchslO6+beXU+3/rW9X9uSC5Ccrkcoy0oEMcEKRn7GMe5Ap7q
chc0BGQe7yfqkS90xenpryjadXtc40wwFilktuGa0A3w+yJKv3UkgcyWB7mpBblMKIcMSEsSIcFz
/6+VbeZcy5a05tJZlQIoKz2UHIz4DCfyesW/Wx5FFFO1q4ZDcHGPjXUsKcUFNDlFEA6pBpaGkPn6
Oy20q98mvA5XLfvDvhnKlHxkYvAn2dD+sjoupcnxZnkTOb4x48xNPEFIADCssXDa5p/2ZLdpkUvq
utow/G5OZfyKMvqszh0+clCL8sgYxT3O+vZz5ffKlkDqo1rdR6OkPWBU9TnrzgXtw+okEXaO4gVM
9SRGN+M3wfETMiBn3x2xXkZO50HmZW0erTHU0mQUutVqXMOOxhecITiIw8FQ+NAhrF7bfY54KOI7
bca3eeebqBzwipgSNahyOhnEcM/uVw0Asdj0jVkt5n9j1yLAClZbX0fEN97Ly+hZjiBvfWkZzziD
PYOfNDuOWVHn+B626+Y2rt6sf0XCYSRxgAyCMzkBJX0tplKVAUD8j2WdTOfnDw99iZAZANWp60Ir
PoX9Co8p69Ay0GMWuSHu6zD9++BynSPGBo1vCBGDl+EFOIobeKMpD71M7ynI7b7UE1QRCeBF6CEC
GybX5zQ7W5FutiAuCvWEFZbrz21GkmV5e3RGRV+mOgCmMKKjpspLLmy0pOHz5GpZPf2dWr9rf5kA
wiCJiIZfXb+FBUe9q0Y+Liy0+9Y2I8eVlUEZoiiEYP7pOIiNaoa4TyO2DDcgkHxz53OQndKf+Jm5
zchXAnrYK+fN5JxK/3QzJFE89pFCStb23A4V9oYyvRfAVl5KmOkarSKJlEzCP8uNAyEgA2faQ7R4
KdnIxoooweFO4P+nVDxQjkRO5G8Q/c62WrPc93S5QPt/Jmo8+25TcJ01cD6SKok+IgShYZ8EEQ00
kl16kAtfLvQT9janXv1eKgiJ9rS0h0zNIAFJSJFOXd5ztLQnUKG9wlPBznnTW62a1B8LKqB3oaeN
3/B6gE+k835Yc/j4QTlp+0cOTbGgrkcQ+LJXJV5Lr1xNal8++PObrZ9alDBAg94Z1NP6vl1lCujN
aai9+dSWXV2NfIYcnnWIY2wkF2TtM68iSzqCMu+2mTcLI+ZW/bGsaEwDci0ECUGuXgrieODyZFYB
UYngBCMgOvo2YvQ9FQ5IHdWqN/LmA0nZSLDeem4CZ/obTwXcw3Aj+L6vbSUdKANsELOYxKnb0KGm
JMYhdV16iT5+2Hb5y0+rGKDRke5pWGdQoEJE9OWXYaBr9Fh+TsxxmZsyA6PJR6A9Z6BjfFjTkPS+
vgsYvicV0Fio3RCpoWn00rt/U+QVtAn7KvWU8R8u5q5eYJAI6T8nMc+J97dlBwqSt8HPYR315Fny
QmLA5n/i4BThyIAac/m8G3BMCC1p1t4N4Qz9n+akvEAnvEZ92RaFWczvNSdlcxwLJsQjlmdwcdta
OwTVRP+GVNub2JHcsa/YMvrDsGa6+U9t7r7bx9UdmYHGN/G3vBLa+uvjDVX6JUSubHyxcJocxuGH
PRwl1UJtZ5N+QZI5p/Di+DouzhJgwQWjzTohT7LI2SMGfQxoPtIRZxfp1I26KbwFs4iv4CgAi0VW
cQvuZ9grJosImpfmEfyID4BwtB1CzLDCAWb8vt0xojnEWdhtB8FmDxKF6NA+6OBrqdQtl49R/sxc
o/bBAYw62qiHgNBKsxdLbv/+Z4lxX/n4Rya/Jx3d1HAzfQHnZRSraMDR413etRkFk9w1Jah8CyPx
QyXJM4lFn7y/3J68ZN1HKCu/EGP+Zi+RYRtB2rOLWIMQYrOYVPodii4RTXMe+o16zx2gARkGgpde
rvUbMZwbkj7Ygu1RGmHr8uKYRPCPKDx6iRn7YAVy5NOQMoVqc5do419v+kskKlqyY/jKw86hDnNs
kvLRRPFw+v4OUc+kFHmcLQnfhVRXiGdZ1US8trzx+teABoT2WBFQaC4khB/nshUFXeOwf+deo+/M
lZ9XRIDKHWLf6i9bxmnmXwg5pheFCLIskzYLAKWE3IcZuv2zBbrTDPLF4c9r5kfXo7Y8GGNcHs/T
JhewqdUTR1QC2le3brQ6SX/6Yy8lGIbra1w1R4coy3WXxN8hrIJEcs2mTk8/rTmfhnX17DCOoNjD
xxrT6L6p/Tnm52b1uaCQWFmF9fD7oaHHiV6zirla7Rws3+yf6wyPwbhw2nVXqRZXrl6f0lrdWex7
WTYkextoNh+DXqTGi4MAvYf+7GVBZp9Mvt/Mf7b8eKE4irpfqeuZ7+EU91rVIJe1jsat7nY2W20n
ABkgdsoIalxuJ0etoGlA9dgS0YddVkl8kKGlggxUX1aFHilUKEGDHWCKmumAqlHL+jkPZ3ngUCl0
b6ayvYJrv93Yu4pli1sUpOvMopgcCggLL6UjfucxrLz7C45bPfifoxXm2dMITq1OMpoxt14qa8OE
fS1YiQ//nDmCdqK7sW8uez+pBVm42+LWba3JKnKdJLkn7CxecjgNGF3aVayvIEq6kXhmspTeJ/BX
NxqGoRo0/Wwg8ZVAlaa0T2VzERcnDilnSjWJz3kz1gjKJtX1PZgpyAbpTZy90c8KDJOOehpnlNVQ
s7fmFCIVnaXwrpwzOOW88ro6LR01y+GcVGD/X7i+TDHTgsI5NcF318CrRHZuR3xXk83cy/BNjAAB
3yf2TyugeGu7eIB/aUBxflU8UhJKDY2razzXDYT4UIKNCmyivx3SfifTIUBkSv08rA89Za3hYriC
x5DfUJynPzY7v+zzMh/TW9DbYcxH9/PA4KRFjLEqA0hO9+tI0J8i+dkrQOZ0SbiXlfrl3U0IQ+sp
EtsqmOi8NJUu1Gw0CGQn95nrjpcymQ+hr1S7VDhmoALC0MlQ+/jTRCIGYUozOLpAaKbg3pjDBWM5
iuJ//+mzkDrHmTmXvm6RUcQStl5s2MiTVbZaD8XrVKRqH6WwPHzK+qyboxNrhHfg40ZsMawUOLz8
VHoQz+u7pt7WIP/JFMq3CNE+JO26Twal/w3DhPmkh9/NuyUiABZKICJm9nt/urN7Pa6wuyWB071D
d5WOLoqA3Rm45XDh5EvNkLMltrSSLLQEp5hbn9uTg6mqwBI4K5qyZEsxdl11My1cr+I/TxmcyAsj
2yiLKJLJv/qUAQx1Ya1VN8mKC3G4YOHx+Y8JS/MQTZWwz0HTboKD5GPWj23v12ZXrq+FAq0nxSgE
SajFAfdg15FNa7cjEMhhcqbp2CCc/7t0LUQksAp3+rDJuju/n3Fw+PTcg4xZiIhGVaNRViMnVfcy
7yGIhwd2a3O1UQ/UZgpTjQaWWKBzZcQrnBd9f90iva7kDPj0ciB+H2CsfqS9ni3pZSU6rVo/lwvx
HGiyuvgcinuq74JLa5AkHU2uocnatZ6LweJ8OwgGo4ZzhIl7RnHtl0MFpt+dQQ2scqiFj8oY9Tze
/JQb5nY7weHiuSteDdrNwC6l3ZTZnvPMCePD8ILyuPxaeZwbgSWGC4NOzHSNjbikrvkCj+c/99T9
LhScWCUo3/4wzpJA+Sdrxf9evCJqcMRLor9zBWCzJyE23aN5BS6Uwhqv3+uamWr60gzN6LphYMK6
1H3OPX6+vKo8z8HW7on+oIdW0fJpm+zuvzdwNGQzZXKpzlgSOea9gGxq2HqW96QKhMIwPQChr0FC
YHGlwEiYKdCYPrlhTpIOsvlydCftJrF/LbMJohf/QAUxZQMTkHoJvK4E2h4haFs3gvQ0fIUgSEHD
qLUiQ/OejCt6qCfZoSe1YBzQDnpyAuPNKFeIKPt3GaAgaowowFcSVcx8Ny39pKrV2cO7oeC7CkJd
JKKtU1q5qGc+bFmewgShwjQrtSCYkxwCT3it6WenyHEjnFHe9UTFsEWVBckW3xGt3EUV7KYlwsw4
9T6wbF8Vx/Dv1JITW43DYzkA3ms9Tf4jUt96YEWUoXTIFPNOGD5Pm5HQwbwcW4tyz5HM/h9R/eOH
nFHjZ2LX2aYnDgY1y5nd0t+EmhxlGOdjaNuKB7v5Tb15lyFIdbWu6qH0uxvoL9M1nBGUUTPchcB0
goK+OlM/R9Xpzh+aZGXWvqM4uTXCgWy6vKjqVkz6W4KIfPUwd4tToZRuZ+eGL1EQPJBGRVPJmug7
R9hmVOU2eSeXGjcv7UppNyxKdrM2PtiA0SBN03gJNV5Lcc1Lgl0YxreGjGagTZNsQsOvyFSsLsFo
RqNnLTDerKRhR/CyCCeRCbCXNyHYULAuzMQvpIUnTseBk2oW79zFZ3BPtToKRbKW/pShabEN9+9X
Wke3RVIHBkW/8sVmJ217Q2on9VhaRFSaHFepDXms9o2uSrq5HgygsZYH1ezpl+MJBmrY4qILbaNz
GhFOJzVHoSHIvpgMggy35DimzjSFkRUF/BllL2AEyxDaPlGH+S2otB5iJJvlty/0q5tfcfQ/AMDi
SceoD3DfCmaURMeRa/iSc6sPfkt7RjeY+6skK5a3g5vmkHUW1qE3SzR2Mnlkjwns+zq25pGufPgv
VLUYrdA2K0IjyH2LetJFG1KgaB8NGU52vQoA9DEKPVmUaDQ94TQjo/9lhKKXYqj1WP8fKHh2NVA9
BG3tpMA1dvvLhMF2s07pFph1WP1MK/XY+x1CP5utUTzglH1O+WjT1eHg2ZOl1tncatdgNG75bv8e
lg/OjO2wEeyI+T/JSmnzv4RS7zTGgVBiaX2ZZHLeXbAO6yuy0pgdSVbBB9rV0zHiTVddNyHJt0+d
O7vpyadZ2a7IgFiyrWufSi5dncFt7u4Wj7wFV57fgeP/qG9/2OkYCti6WyMynpWgXoIvTTsF0M3M
zCdrSo1N/l2P523oPROUp+16f/jN5lS2SejTM9Q79n/ribAXjAxfBJkS69uo+PkMZGs9bJqtaJz7
VzLEeoHTDnSSoX1xwtfI7xLTIaniKpEHG4X0VFrkMvG2i6KAzFe7Zet3rbfscP8wCjGf7/roLV0A
In3UK0RxMA6NPnx6ip6vGsSHr5fhQJUXHy35b6Q4+l7VKvh/k+Uw5+025Ntr98zFgPCV4xd7FhN/
Kg4XFOtp3sHexkPH5FvqG3OgEVyt+ROi35cVmcs3iXGaDbRQQ264jsVg2fnkijMThhYPFSyMKU9K
46IFhCdyu7tFJ+VZsDRpnJ6x2nMU4ZpqW1f0zCVCpke8sEyk12Q7VAGV1lnS1dEZub+JD0+IQTy4
OYbHvc+PZrMzeW3lzoQFt78Z1HahwyiZNtg5scdyy6owRf7LAXUJqA98XMNj7bQIXPCf+d2Veenu
qvP9A1O9GqH/5OiQuxi4JLvPhf4Mlf3us9dkofeg4qMkgy8hfiBdTNi/NQdgnau5eHxE8iuGPMQ0
NMYeXkXNKa54SvwtoiXNEoF1Qgi2RT6THH0G13GMwWxWYPvbT9dOF9NvyGHsrOIp+aopKFz+13kC
iiT2ZLL0nHun4kl2rbSWeBroKKN3bGnSKnlDHhLVfJopfiPA2UREQHMSNa+EVDXt4wKUQQpUz8FJ
/pXm+86B+HVHs58W5IHFYiThCzINLZlyth88aPxO3jxHurYPhc4rV4ST6BZt1WvYrmhJOz7c9Aaf
hsw3wCMTtz6h7RGWJqU809wSxserCG70DtUWhtNzMhfWslK/31uKU2tRwwEJUTR5AXRpuCta67FX
LfDSkRc9mA65KCCL9nP+RbpBD79zExISZ0xtItuoFZ0BYkpSu0r0OQZJS23sdmJISlo8JBIBZ0f1
bsO9Ghy0oN6QQ4sdZJyp0Us88zAuUBvtbo3btnB7w1c6uNjOBq4zQ8ncf+NKP0ncULkzo5lRC7NM
f/XBOD3qel6HtPzI2HxyA1x4gA2+lNuKE4snSr+nzyeNyGiGXwGqKxcF1FJisu1onoOMMr7RNnto
yrgl7tPrSXVmoyo+zvgYIezZjT/5DzgMdstq0pZ098xpG0ZpeNEHKjTudu3uKGsUYU/DEaRTiHtS
t96uDIpu6ychWegTJ2Raq6299DQzajfV9m9Q6m5LKpKaSTqbNZQMzyQ1W3nbjIYd8t2JBfmvHxtP
1iPNGbuO4j9zr0Eeqiivo/41eM9IbYqy5QxkaZk/3BhFhqT+yUUCrP6+nk2UnYiZlYcPY7KasqSk
zheKz+X6ZUNS7Gpt27QgCmzkFAsmiHsZ7yn6HmjRIsi9deFFpR3YxEO+O2dgi+0WlWjFWRW6YEYa
i8Whu+/JliMTL0EOvOPwjoaYQ0LizcepWgbeZawXsbQOgMtNNNRlRGsL9daqzcTb02X7ez424an+
kC6JUQwPdAqYUWj68lopLa/MTeBC1z5x6Fs7y4LP/CAe9md1tj3gmQBc9/M/3E62ninmxccJ1Qj1
5TU4+70B6nBhfaEg5VfZTztlZ1eaBbFmwVHeHjNfd9s1iZWQADmnx/exp0/TBVuh96sQOKeVkjCd
otPtyiI/W/w4LOjFtmtlcInghOkN25nr1Z+s+0kqsi8duWfgM1w1Rov6/Z8X+v+qaSLqa3wOp17w
jBVvFbefaT3gLVBm2DmlMyoa43ksXj1XV2UK4RFi4ngNwOaEqavD1Mtdav/lFsYHlvXPw2tmYttH
wmVYLNcxPbp0LQJvapj6SjifS7ROKG82L22+9+5mATSCGvQMbtPyy0RrQE4X9zXypLRS7BLMDTRJ
uSFemY3lWhqYRDim2s9S7WqVP8iMlrP0uj5dNVO2aofy+T3nCu4Ic3Frkbhm5sLKPVbvTBfr1mnI
dU4PxUyaD9jGiu3cEHoE6SWgRhnxsZLH61FYsGfApldxFdq1zN8m6TDOH7vk9vmQEaOh20PtM9y7
3Hm9lShmhejEji1IFS8JtJPltEsdI/4uVNFoQ5U025kVSm1mbXWnX4w2M9+SbSQlFzRqY09/uwwB
Li+9xEIpl1wO3mY3rNrwVzdeBnQkbbd2yNrh09DTMDmBz5FQLVP5UINtO6oO+2R8U8gXZ4wuJ4yN
woHr9L76+l018TuJ8X+Wjk5DoCXDzjob9jnXhG6YEdrwmViIxYLjHs+4+avMrJr9jsVmnM8hTJ5p
63PCL/x0r3e8hmSqA6SV6131IV5fEfHVoOQidOP8fz9Drvn3hsnoLCsuRpErexxz+j6x+zdKMUdy
DQrTJH7qKtsxXNLDdnnHsqI2y1KfIOxGvztoYDNtHCjH88uwP/NWEVckjzpPYMo66d/bY/QVlQ1S
YWj3q2YxTXyjBKBFLmE5Rklmpm/PXNr1zCgX2YmV4JGSu3GUWdbdct6V+7Ng0st7ErCHrHLJWlGR
ZLfSHtMFpOkUijC5IMQOlSSuxvrc7fEaZ6uH1NfDJ8w6kadYntXf2RI6i/1UoAFDm7Y1OJBUAVzB
DfK9nfi7FEZw2sosnPSSt3UGNBuFrx06at65tQvYLvr5lFr4Dmw2btNwtx8tRbw7xK6gFqv9xrqQ
VuFOcSAWwqiMTZV9uJVryihLC1KIJKpFJXszAZ+g4HvWdY7eUTiz6ZTfMHC8SFy4aXZaXMSOHhwr
byRJGMBvYM0edmiS350MC6iE0LAUXkyltKv8MjK5ifiLGXNrKGriKx/Rlc6kgopqTalsK7RLqAgD
3vNA6Zoyhtw0oD+pp84B+I7umaT+7fogv8fACyWrxMUO1S0dxJtkl3s22M9+WymHPJpkTbCRS5s4
Dcv2X3F0MLuZXwukaHg/Ek0lg+ovvMrvBCntItT/Z9n7G1zdB9754CL+jaY8+QYiKjg1XD2ccykU
KbauTzgH38+nM82srMlvJLiZbIeCnza77cfxn2pdhNgeAuzlYPd29CnKaLMmTV38ru34xFnS3rd5
baqjv0ok2U7C98FFOXnNdbETW2kwNfDVKEIR8S94+99MewKXHsYo8t8/L+vZ58qimW/IKp7sieSt
PcGfb61yIUuNi1hk0jto2qoVpq3cUb78Dm+F21gWWW/PvNFuK/dNk3b15HEpeLjf7LdIzaMbImHa
4mgrT7wz8EmC3VtFmFk3KM0/0E2t4ydKsJrtzRD9m3120kb1XxiCM5zH5/yO4X4S2UrhlJyBgzQY
7dIDCMrdr6fYC9TE5yKEjvv5ZvFfSdkPUBwu/MYnS12zfZ0EYAXUqE4ExmKEb8Zp7RwiGY+nnuHy
pv/i62u4PoeWwxsxRU2bmTtvvoi2sECorTdwxKvdddVeQIrkYckiBcbMTSOlUHklcTrf3M6F2YSq
dH5P7kckO99Q3ZbElMzPNgyGwZOBtSfJIO7urfUIDyN60UP3hHfpbaGCCtkrez0grW3ti8MnP9Zn
o9bNTyW30sDvSG9MfXNa7v6+MA1PHj/jkIQMHN2VDq4bW4sfQpa1m9YfVAbuEEnKAYq66TSHe/2q
R1ijgIP4CcRrMevzE+ZjDZTbPr47GglEEMa1I6j9po/brPkdj/ZhTSDlowd9cfjywb0AwhNshXIE
UTzRHuyJwToYqwHld+DJBv7gdxIngykm9zB0vO/aq1RRAKuVOVM5TeZRNLB6cmbfknH93SpUA/ex
A71Vt+/X3/UFPuGSVh3jO96f3JNz4goRirPN+IkGRjEEyeUzc94ilWM3zd8H7CnKHKczBA+48PNg
f86mQ8xiPftB+WkaJbaDEi8pgT7iRolFBUSajtZMWxwHcxmafbMMmc8yAdc/AOM9UiduUnJnpn7t
h2b8Sm0uqtyRi59NOco1ImGa2wvqaPLAWw6G90DTTng2sjKk50Q/M5wLCGnIVnPye3jIsYWnkl7q
Kona8ARykyro71QXad9VWPuF69cypMhu1MdPjI/cnVvUgY5Jp9S/Kfo39vghsSp4chE7GIyf+tsN
53l/d3YeLv7+vDaaHK6rGIOlwCF9Lp8mrI/QefqfwvuI79eUvzd2GIkjDyGkk1OMyUVd1zf6P0Wb
DvUuEh6wmlA2Az3FjzA1Oi2SlPLRUt/5EreDlld6JgLio8zN1zgZ43rYjgqt1oOWWoNOyZ9Q74wY
9B+IchtbVa/YhigQPMt2gm4m9UC+J9z8taWQj5I3RnH5fKUGi7rP5uBemAJv0kcL8dsb9p/1zfd5
3tRhsuRhJ5Y7SnLqvS52lSR61kO7kZJW29yu7px1NvidYNmDZ7f/I7iCditGkOssO0fdD6FaU9cd
CfVxNPHjm5aIHq1oA3XKrozH6hzdsVNkjbEX3qebRY924N0maAaIaF673dYj3QvXgjEc++XrZV8p
KrK4jR3BuVCvOXSH+z5qm5SqyKEPmiewovG7tq6VPJCbQBcCwikBhnfQMwilkJGmKTsQAOFw8+/2
VBHbXpCtxeQMYnSwJ1bxRY5iDxBH6kGOnSh0KVXUlP+IET7ENg0u9czV7ZHL2Y2ovH7o3guzFpnF
7d4Y19hhK8Vnejd3BVdybozjp86MsCpcoMmyt93YWTe9ml/dV9KTKKzkskqcF9MuQ/rXejLPC0me
SvrtMSdGDnsR0XztsAHfTHKf1HB4sLEUXXNlrU8t130dJ6/5p+ONEnCDLMVsqA5zE43zV+TejOjb
o9UAVGsccZkx9BBjTutyL3AzwcQZMy5+1VgAVaKYeBC1nWYFxBTkQicqjbEGZjh+pSZ02IMDJLgy
K5D2lr3WlWYAjo+cxo3F+AGmVL0bW8+v2k0IcVnVJKMF/EXap2jIK+TShnhaTzPgijzhyI5Z4Zb6
lf00etJYK45uUm7Ysu75a1qcGdcXXDP1W/xXL+K18rYBRpDH/C6sgAiVrjM2u0R5t0GLNZvBXJV6
ED88xdyDNvy6+X7Gcpzxt7LZWISLCHTUz9MweCKDLmq9JZrfQfjiAfHhPTNIEN+0quHYOKH35BJE
2uaUBPNXrFBnIcvTAF5PAj2TQiU6acYcWxy6JkjcZLWJ0r+2QFh8TAeVqLiY1BHAYDrkX+rZju4A
9f60HsOde+JLKKSnBRfC1UnhfVgqTQ9I/RhdqFhucyT1BP/QpFHQaCQ36Jy+sm/fIUxhrFfv2LxJ
YEojwapusJRmJE3JHt+Fr1vyfJCStXpowAc7kVpKi9Q9qbPHgdIYm1Mow/8qMH4tQnt8CS0Sd9uu
7QlA8zxxjXjDjEhadTfRcQ+CEDedCT0oWRwLapR0b7twI+jNGN1LPTfciz4TC3MaDiepRBJt1CY9
2XOfkk/1irVaxGb8Ybd1Aoo+Q0N5f1rEcgNfcsoTEa1UUY1rgQZkxOMl5th72gE3fLdFX3jOgL52
mXvE3Nhb9IULlFdxPY5THRqDBC5HxMM9zfmxczrdGSbBgcJdEF/2AG/8eRPiJmnJDPuDa4lyHGk9
CTI24iQUTdmnV1ogpNIYub5919nGWnb3RKyEROiqtwhEOaUifL0kXuEqvUUhZiZkRxPVnkeFgn72
iGxJxC4yS9O6uCzIwyKN0dGRWAQUkjIzCFu5N8DzxEIXn1ky5FYlMN3PzJMMfNOo/83Sw/40ep1t
oWc7qymdci0VVcAdcohBGmkttF2UXNz9FVijJDmNVG/+QGtCKOegkGEsS12EcwyfeBtJWVxZ5Wsa
37zTSChErJRAQFijpMB+BwMKKETCGDkGEWMlNY/RUixR+XILB4z5vyBkjNtLuupv1NFwwoU9Q/d1
671dxeoJiBJLnxYf/RRuHO2YAxxtGne2RE7/kY8UMAmD+2MNcQctYRb+uVaEzenbqPgmdDUIiCca
K/Y9E8MhQEW+6Pr5aKyqthDQpPBusr0kf+vvga1ARui1CaGhrOCt5YENgK7eugFZScjXApfF70v7
xs7BqmtsZzVd9PIO86zmOcNhZN7Ruut721RQzwb106RRU6y54VY3fGaFjxt4RqFLNa3gC/kx2/tw
0E7ufFZ9+7TCcikHZ+cnL8BwNYA62pnwLHsboFVvMso32eYodBgDfwSumZZo7DTrhLtclhaq5wP9
4oQgv1BDEABpTAsctMDPAukQTdkC+sp8K5o6anmlXXWzVa5XjuVHjg5eYZCXsIyac6pdKcF1e1Mn
xXUXRpjhNxR56smXpzhDhzr5F8d89/pSfOYVDJv8cB1rZTDO30gb6yfoMXromE8XxjiTZ2PiMrr2
xUX33CTnetgVZPDlDHNSGOgm70c+XTgFtd3D6ppDknuqWFXxoKEwFp0tiSmrEPNYTYKfkBQcdW3a
/gHq3DpLfDiLGccoIl7uB52qtOgFMkITcCwVS0X/ziPv4/cE1ugq6/k23KZvzhpUo2jzsI6KwbiL
onDWZADZ8C5G6nxXlu8W9AQsvSamiDk2vZs4jQqujtU01RPrnSUdpSnN+tJwsO5PWhQvTi7aGj91
Uwe+SZt5P9/+46KfCZ9MRwG84PJWFFIr08SQyofWKXp3OlzXe1tptV1b0zjM14xa8N6H5TAkdXXN
gHRRI8hICE2MYetz3ukiuYljUqQUmDx+dE5nQ9CmDSbej+gQQ9sAwluskBFiDWbtmjG99Jaw9aQP
MYCuIxBHAlUCnXVe7+Csbo92rqeZ2+bZ7mM3s7LD7fv+M2jrF11LMC10oE4HbtRra9f4qYo+3e75
5DRitHE2yIX7nyUss6HYTZzrv44XzrTTBaf0m4Z+3n+C6E1ryzrLb/g9zSQZvzFcSqe1QReJNwao
DNwIC/EdnScEU3e/7XsU48zR6j9amxV5snd6MeQ+pcScj/l23xxxfvN5PRK+HRv0SGQAL1x568al
1rngUd9MxYalzgWH48p+jPXAJ75LeHJO2iHAkEGftP8II1wkVrPpfaVo7u64k7CMHrCVlgbW21j1
+jy0j2ld4Mm1DJBbjfgZLvDV/1NaStEJdzGvL7a9yhgF6DJff/+pjAZ0u+WEtQkPawONeOPbMiyQ
6X9087B2IB1wxT9PK4psqzFOunIgpouOo/twJd32vSbBqcCKqbmM8cTjB+r4d36361rQYoBUD+M8
8upj/qUkoNXrrggloeuY35Z2+2FSwnAJRe2VYkXTgW/VrDGbvLtQ4euGwfruIwyLS2m457qmPbat
WL8UD7grYDRE4SDdoTEX2knD5b+BDs9KpCTssO8tb91+Xhd1S635qw3vrt/zSNFOhKmcUfNPu1hB
kBFW4xS1nYJ/36KH0NoEgqnj2pUWzh09ucFmCTxzCpXumVp2yMVd49nTGy6/nIWOXeuyYyuqiPUq
qICOeCfIHSRAZnDlfwOOoqr1T6gjPVa8zYLfITA5p9+QyVWrBJY+YQ3r1CQ/1zZqERGx9ctkrzJ0
HJOwNhNSDyjUm1cQP0EdALo6d3n8EgkZ9g04rn7EAYKxXDB7QEg/5AHPt//Te7HlkjFgSxK4uP48
SJ8SSX/ipNuwbH8qJT5pvBnujeX+67WNtBViMht3iTpcT3omst3W6ymJqZdUm0SKCQOf7Nby0gSO
KD8aPkMHCFTOMG9TqHJojy1Iy62pvtnRcoXGPZKGclFx1NQENycJ4e7maJ5NcKdPc/xBDt5bpVOy
gV210biFqCeRECwT7pJm+OX5GS7wUXYXtvdL/ruiPuzRCRV+T0Ud/2BBn0O1qup/9eP/9Vdaz2P5
tr6ZEVMNTyrKmpIK1uNniYLxW6ksCpu3Wuw7ZoVcACWsaLRGIGmZf8mc0do0jYoefav0/zVlkw41
7MKJj2Uk006KbRnihCESVuWdEjp+A7gAgSyB5VevVu8Qa37/1KR/7kaiz255ZpUYSyGi25D5yY37
KGWuT1jUptIJj8lpeWLeeJyI6na2HbSOcxTrYPypEVPcZcOP2UVsnsAHwhOiYn3AwKaAjnJOveS+
e2s7gV5WbIsihgXaB0+HpjUXEz0F9Q+lWwbSN/YHCbNOHPYUMcnc/q8upmlYBIrTHeiDUh9R9rLj
j7anU6j5doCBMbWIS028oi/Ccnrj8TBM3Kji9d6L7GviI2nsd/v4Y0X8MmIvhQedFaPAOSSOnYbo
sWceP3Bjrn6TJGI87aA0DL24oGscBvvd2XQKAAWcowi2DcYdlJZDjmGxQhf60jurFyrzX8xW5Jzc
Wjvhih+P242dI5NQqQIdL4fG+a+QOqtOeZvkoqwLrnkS0IYhfbYtj68/Rn7xs/ja8PZaHI1J87Oa
hUOx3ZzddrGeSEztbw0rTZsVwreui6Ex61nvZV3USiMOsOcdaKIMaWScnFMNXFf5jruSW2bvb0g6
w8XbnJHSLsZJunVLvAqdGSdjp/5P1og+zmzLGAu/ICV2g4FFK+XfE/PM1pZ7x8jrwMlftHqYrmE1
Hm5k8hXR5FzXRmpVkFVb5H1kLzHBgz7EKElL2gCP0FMUXNsfpDVs+79OPPbnOgytwvXWGS1g22ZI
YEzqcfuUm0dEdjR4fiUMrb7HRY6OGd+hvbrN6hdrodaOy0CXhbvuKzXtN9SNO0xwiuP0Wjy8vx4n
vgIGpAHj7NQ7Ju9txq9rNkGDayatnVzVlz235dmF1lf9H3yV6biwX/0tllQasJbob5DcjSnA4dZR
oJjIMcd3Aa9HIs6AHWudnNhleIH1g6DyG2iXQ17UYjAhAkVlS5SaqrqEoCLAKp/l9yMXWFUy/Fpc
6oo8Zp5EkdHuH/eM+K7o4IOZoo+zfEQXn0guYBHjiSZ45ei7TcyLjmQ3mxRIhG3k6QuoY+bcQsxD
8iZFCBot8snMZIBZFsZvp8h5FPOAVS2l/P3WtzekOYg94zYTtd7J3tclRaBDEgPGwzMRgqFFAGwV
7tgLC5peUGR5yimDwHj0S62xe7pB3hfuIerUM47J5f/Z0owXyetLriif8bFLW8v6GkK3uWFc7+zD
4+yxvz3wr20N+Rs+NiEPfx2rkAf7Gj/inH8v0ZeK/bir2jYvr8YV9ExvGjF9XCYqSW0R6ZcebVRx
Cmorft4vBzJbytNrWojH5OGy3vL9Hk1vfjO3wlQlvKQ32kbqdvrUvRW0f0cHKYxvnQlHcWXzT+/c
zIVey6fcAUCZ6+mi7i5JugxbLSrjR9nIhydlOBkqGo07GjuHR2cblfBYJ+kguPoPmnWcBW7XTHHw
O+sPSOUJ0omU4YWthsCQiF8FsZibu4J4Cd4jBLYnWo5rghDOylRU3fvVTL3BLl9pKzR27aa0PEZz
ORNL5X7nLk+bnFIFHtcSsf0c5IiegYEvCy7G25pFnz0F/xKmF/RoSO2JS5QcjUXudZkksBXDX6OH
S6IKtymHAMu1agoRPJuVGOMmDl5QDl/Zx8VGRfLISDlEs2q6sgfhtsc0ls9M31GEkH4uu4IDU7U1
P/q0ttzEm/w5IhYrR7+LU2FfaM/xbOoAhEBFFrdWQuI+D8L521nDTdqCYi9HApJS+OXyW8LBXMeb
7/UplXDi63X68IF8NT9zh/dbO+7ZtxJhlz0vIV2GCO7GTgboElNELNHM0ZPYWcqSKauiteEdedGt
A4iljEZ3K4/IClbmbeDyhoQjTZ2nz7N2SWWQR3/AMmUt8/+3J07KPyzPZsZouJwh+OPo641KyPSF
sNtvYN23LwSgkAK/a8RpbOC+TNIKG4RJNjKTK4EUcuRro6iteKCLlKAd7d6TlxnBNoq6CjQFWSGQ
7JiCZTK16O0GCVXiz1bqDG5RP1umDlZqApgNGhP25vyQKfevPIZVsBuSFplokSewWQz4HedOn2+7
SJv0y6pg1PJRHKbpV8V8HfFYszL17xWZKFY7x0a69+SqqI/++DuJyULcigc3E0VuzSkJf/m9czNb
gV0Ww2b+IcOu5TrkHySxSim5Vvq0kXhZKAZFQTXNHM6hRg6s3l2AK2VRZB4WnDOPr8WQLlqoPD+Y
VDGO4Hu6kN5QrJ21lvYu0LtN9Khhc+615bFldlhWC/sWlALfuR+EqgBchf7ZojpamC7E4nk7g+wD
bArRLjpnLjc1YvPmORthoA8tbZYuQ7Lqsstk3MS7Xw/iciaInV6mXi5FffALKI0AWdFMfDwoRJGW
wGlMfDPEdsVp9KnHH0aj+zyJEnvIK0/Oezvj/VJQKwWLNwqaklVLIq+HdNoa+PneHOHYJfWTSNb5
SmGEz2HxxTS5/RznSUeck0nTCt8zC7d2jPb8I2mvCIajKQK+lM7FGKkMvG6Q4KmMY6VkxB3cLASx
NB0pmDRrDD2KVyvsroEWLcl/HO0qHsd8M8taT9aPJHepVwIpnBntoSlSKKaX9/IeR/G9qEGnWsq8
AEg3gn2NgBLoR97lT6S1yEDNzk53ZUTqsTmTp8XU3LMa5ZsxyE9vIewtQHHzJy0yJQPmJJ5bQvnu
3o4b/fawCKM9ofMg1bWXuyat85Suosb4JFnHOrJO0OiXUiMR471HpUFPIxTYmF753JYtzVcrGNAw
AJJCr8WmrVLDPAHQqLDhfedtaz+CI/9cV3MLoa7lnb6/ltVXeScrQP333Tfi3b8W9LzQng5zzLH9
Qm55dBnG45WfhEFjDOEm+wpDAON2YfP8UTtd77K4THPsWV+31XrG6d8Hsucep0Rn4AWr5wSStVQY
lKGCWwDzkycrk0PXvePy0/fIbTLQV2Ciy64h6J1+2urpMiEAw6CRPIwo7PobdgzCYtbm+qw68qCd
fv0J3nGlS+movOfuRUNxyJadrybveVbtV8cCWiZnFULZhUJLISYBW0LMvC8jpaVvJpYzDJ1/gL5x
uYboXCFnZhNxFTne2Ak+qy4JG5psyigwjWL/EWOZRi8Zs9PLWKMsEOmD/GSVSd2ydOrkqKZZX+dT
28Kp9YuPhGlNOIotE6feDjY6/ywKSzC9FFa2yel2SxTnECY5oYw1oKkRUkmJ4GM5tCQI2QMKlz0J
QapQl6SZPkGVF6SmsP/mlaX82zQQjL9tS7MyCE4TJmYFe5/tad8PFfjZ+IZbrB8ZnyvRx6/zqmuJ
/EigGaQst+kqaMDN4yiplP/74EbEKF2ESnNt9IUOXSLF1hu2ou6i38F5RqY6DHm8VBvsGM0EGz80
EgoyW//pYcRRkrvI/aWd7s7s3zDANjPWcFTXGww4yBsIpxHc2Ynu9JSviQjnfJp/VLLu5k7DPhGj
VFD+TT+W7NSfkwV04wceTJFQQgNQ8pccPe/GS+Y7IEhwoSK9e6RvK5hYG/QX0a7MGhRixe6nmW6s
tj1q2+o8Ny4bzeP87QQNPOsrF+pgjudDHm4MIPdOukZhnlmnVo8dqlty/eAk4J5Nona9BLVn2+lC
ruaN85vD4PGxHbbL68v9WBaeSx2+ceP+nA877spwZLxmwldaQflDGXIhUH2U8A8CXNZbetSCt6l9
7g6d5SnRlhtEKpCbRhTCITuUMppK/sK1cyGLZyVBD/rvLbzXf90Oo+cPZpPwNvx887rCCqZeNq2z
OtVFsRHRVSn7G9BwQPBLGJN6nacHi/ipcHEJ6go4G4kjUYTV9xrk1/Gg5xKzgVI3HAdBb7MhXe9F
f379lhA5g0TYF2ASBCOarfcU45JYf0/uN4NTd6qWr0f37BXK27E4WJxpPCMRUJ9DHSv2arkKgtDA
ekNgKSknQKV88ltWGYapg9u3FbUzejb4uQrAZC2c7Ve/xGlO+3KV6w6RKWYtqk7LdNpnwYLnhhBu
KxvMYgkuD2ujea3OnBURqCJ7RV88AZVqBO7M/Jc569Rx0pyVhFO10rRPXN+zMSedIMIBM02Jq4o2
Q6IguGdddFX/gLvQUpl+6qECTuM5RzGPfbGKc3+vJ4NGks4VkunfPTEOfwReLsX65pvLCp8KSkoL
dMp0ALdvK4TjSF4ucw7MyTay5ypV9f1FHB7oNRrCeBQR+DpHQxUHO2o4srVKPg44X4tUkAeO71Bb
Jm446EIfP9MPgGhjW4/hMF+/EVx/Xf0Wyrfyw/8MXdgdvb6ag4oyixlWUv60UfQ22MYFLLNQn+re
RBbxGbed1MdVnhLKU8pqjjNzecPNR5D+qeRovmwKH83Bq79rx36gjThaFHiMH6tQhQyx8WXE24JG
L6VL47eYp2z/LfLkC5EzQtNsHn78NyuGPJqIfT24hJFvKpeOb+osuyr7nREQiFi5JfjPZ3VunREA
UbVaABwb87hMmdfqpHfRM+4TjW4fAKHcnFEEWegYfA8NMwfMLnOj80y1+miOntljQ29zpa+L9mTZ
jkhe/2HL+f/vCWJtLlE7/YQydBG3adtrrPq3v7Z+O26yXHibUI5Yr6gKWa8jILVxudv5UMw7b02S
idwTHqUQyL4iqpexurVDqmDdSDJFVsbQk4l7R6JP6i74pyWPrgYGninZl7ueq6fhqTMg6bT1hpyw
926Qn3iTE4HdmeVS41myRVvidq9hTyJOqt6oyjK0IOYPKKtNGVjc5uUZVGMwM85Bqd9P4DoGPTtS
JX/LnSGKn33ZvbPecBwLULVpyuwEkP1GgmjVlFir3biuym8rJ5oQ+5/iC//S+YOkw9sw6rp579KT
CsVSFT5qJ54KJ/6uSwH3LFa1cB4oX8NHOqcN6Y3hn/mfLm0YYA+NRyVbdFigzgTsf9U2wDLLloIE
MewWkEgz0AOtwKsgz/LM28ZQdJflFoopZem2WB4HtTdWnnZRAM7dtLlLBBWPgaRw9ttxKX+1U3IL
RhHUi1hT+yd+EADpJEAi6Sffq4g+m4ZP6kbSKItBXFmpx9JHbAAyo9HumuV9L0NoY0/CfDYVyIDu
7LKxWvOZMtKe3y1Gh17cN7U2222d6ZRW9XqasAyFSqqq2lOAJgShWboCXaX5z8kGGV/CgVcWdN6v
Jhs/leondbyBJZQr2e+qMvclcPmNOaUdYZioHIsVQFMJ7mq2V1lIyxN/IqGAaoA1QCJud7c7XxC/
xll/l0eo+zhykpPoG5hVgLVeNBPigRO1Tkcq0I8cDEDohoZk63jC8bZLJ7XPpotU61iH8Kbwzfpz
1N+b/DerZxHPSNdft6zJ+DqDW8XDE1BQ/WOZhN1w6tvAah0UYaoLtdZNLd4qp8y3tPXMSEIAVMOa
ho7MWkayYH4bq7HXaELToFqqHZIlajGAVHq+LAYuN+caxTAkehVuEKfs1Yye6o2J1RKGWsUFpwVb
OOzlBIHFopvxP6+agsNicBACvE+i5Ha6GrR3xRVz+RagZRetKZuKe0KV2rzSTTUCIYZd3Zkw1Ydu
HJsz8/XSQi4NBDUT/pqpV69Ox5h1q/czi2kKCINee4lykUqXx154mC3wswXA+vbxq/H6Hn/90P/K
DY4ofBADckxB1+2VyF4qMDHBbig+ymzV74b7acIUuUaR0BFZeIfUzd+8Ucwni4AKWycrneLpapVj
23O9txV7RJb8aYbv2K8wMA8tSa3+S3GrYxjAOvZDF34I9+wkm7js+RJc2A7DlDNOOrsDgy2jth4+
W6lUxOa4AM0f5QpbGdeawcWLz5EaU/v7DLdMbkzm1ndkvzMuHu0WUGDs+s9hD5MLdL1zSFiYpLVA
jrlbjXUaFuZHSGgUDH1vAFs7njKoLCvp64eYUvpqmAHIqt+w1WwKewyMKa9G/cLH34rSxqmD5D3K
HXmP9Ro0We7mIcbDmpW7/BvHmjSabrnwvin1M/Bwvt+XqChVUNmrVuOJbda7fAz380zHL7J6tWhv
+jI0gPYGX7n2I+avQy55pvukx0fPR5KkDUjx35tuZAbzUcWQq4f7/aF9qCMxL+0BgpV2oypgV7r8
ganvRAjPMAdcTlUXrQHN10Gg2PMdgwmrooaeuCtxadqsbxv0uQcwkNd5K8+MDcczPeajNLfm88zK
YL93uEOkbFTAVerjvxlmulIGpj3xskld9U7ooCOc65rXN/If4ttXdLteoI2fvfd8FH6QM28WX0Ih
pLQfFC3r/SAUH5bLVwMj6vIRapM6gbuoL+Jfrwbu1AOkwFvkNhL5EqEExT/dGuy5YUeOPdYq4oIe
ZwY1cWXyX4xDLiVJSs9b3v2/Xe1dcF0Zv2IWxyhMB1uLTq4Fj8dutBxgIDuXrmdRuHHQ9jkvZeMJ
1LZRxRoY75UV/0kuoNAB47ptJ9MweANcaAIOwWQAXVi1IyN6bBoMpZxCfokYEIRBxBkDojJQ45zK
FJ6BC6Z5sLbhpwQWnsSKZULASWHlXwCRZ2nCu4PWuOLbrhGCGtx0DbdOrc0EOG5WGHqO9iaO+6Y6
0hM9juj1iN0yRNKCSYboEjxPlBAvl6Q8jQYrXVapFoUcDSU2YyPvstgzAbCja9sI3hDGkWYxvPTa
JZvD4zcEk3tGiM4BcWZkPeXT3zz5HnwCyAvTchQq7boSl+jLKp2QfxYUb+/9KfH7tot7Yg/LilNi
1S31AawNb4/OfHN/XbYgwcAl+KhZdmcpZXZSxL/zLt7PXGFhEeLKmlLsZvoizid40tddSu1k8xaZ
OR/6gOMDQPx4CjDdsarlZu/l/iBWOSZ2AFIqL8KqQrg3scAbde+6TXhCgtICjF5U9FFWJAxYTj7c
EpmfIoTb4GwcQ+DmpcWhubcx2fj6F8pjCaKWfGF6BadP6KSDD2T1nQ2ROeFUuM/WRjEeeIEG284D
+NQyAIjVQqILzzpP2lOF4SMLsKlv/MIMUHnsV0WGM9dFlBuhcYovUbCH91AtYNVEllpC327oecP9
U8ahFWl/yRFhn+JfPd91oWu2qCEE+pjMu+7/luntzpRBXpyhsZE1NyIIhsbEKVjy0mOFApBkGGtY
OaQMiShxWxlporKZRgcNEr3gD37NvxdssnaC2BtOyOp2qxcOMQ1Rq20AwTGs4A/izf3h6hMXOW3U
dmtbE0qp88x5x+6+dO8+6F0f/MqucB94FO0CQtMkCEGlYdGv106AzrgnGe3zbrKFi7EAW3/rFg2K
LK6oKqKPooaoJMEThnyohVyDqXvB8YRWvsKzHjGqkMB5EngvMun4A4lne4PMSuHGFwRQF34qZOXp
1Y+UiSHD2EcjaRJjTePuc2O8DPKfff1GGqjzlpuyb/OEk4iB1Js3KeuSVmcT/RKQoqAeJlB5V3ZS
+rDWlf298ZvALElxTbN6vHi2rTu517nbO+iAD6VoJD/8ZU7IPTawbruWro8aQArwCTPnnL4BM7Xz
PBoQZmNruOyqPFESabbwih6WgkoUNkK0pmXmSiJ2Efd3Jfg3FblNmu271powz9IUYtb1cRaDMB0c
+FTkvyDQWmzZcdEqNzWTe1TGTylZV3LYfsoWRiW1VpBHbN/rD5gAKvjl7QxHZ8Anzwg7rwNtPs9u
zorzl5x0cFckKknCq35lpAXtLORK0qCHZT9qdJMK9d6Zvb+iCSGmJUk+2H8JsN2Tw+wSvIYGa4p2
HxIlr4BLruT0njDG526cIShFhawKnZLOcE1OSA3ig/RsDwanw0/QPIpBHID2FYwE+guqLy2tWlk7
KCHun9/1cUFQm9MtyJAbVGZo3QnHuYeMDSfR5Qcr9ayvDbL+S3aCwruSp6OE86kGLfChbU+1y6kU
/pHYReezBNnJt+kO6i09Q6Fl3b09wqRo/SsuLo+c5tCCxEeWjmXk7tODlhlCm8zTlvctoVbmHRLn
SPecnqBHgitGdY5g4V4Tnb2SpW9keoCwNfztcP0vU2SSG0y97Byu4YD1SPNfX4TMmg6wOLnU53SJ
QBZHPyUxBIBIi4oY4YiznYRJOR5KFFKqZcb9MwBAuynXsgMIVMGNfTQgYfRdH4azEkr/8/U0Gsqz
PNKzF5gKnDtXCcJSeV3eZhAxziFVUbb6Vur1YeTllsFe8g1I1pYt4NFM5PalKxrulZHlGi1uPWoU
R/NKtdM0mnyRBTcxuR3O/pMTfLZ7f1gkopW6Uu0xkQhVuTJMRjcKXBGvu/0I+2CDwoEg4ALqjFKD
p/aHZdD+X9kMs7T+ox6vUlegqK93RGrTsAhBRElgiseYzzrTWqBCJX+g4Gy+zn4guUos040hLjPB
vYKBXe3e2hS4DxoqZCTKmP/8f9SvvON8tWdH6YzsJhvkgQTkQIADNGrur5XiXM73PVQPju/tzAW0
3FNdBzLDcPQeEMNT++k9wQ9f/trvaKyjHh/WCvyN8qsXUOANf5DUshbPo/BQbDwgEUsE3Bq7kUSS
5cwf+fVPz8JfzOTQ2DIqUG2P13a7px898JLvubOkpnWxLBZ+Q7VBNGOXc3SwPpepNEicfjrsdsIP
zI0ppO6asNPAvWkzz1zEqT0pUfcWgUETJNdCV9h5bK56zyrkaHrRKdEvJt85ri4G0LnmgWsQdtQ6
ZXAnOhJsr8gw2Y11cfuw1L5dOFUErDhV5tMHWvRE5niztLgKpVvHOSODOPBY9EZJphbyhqbkpD2k
RaBDNlW2mcpBWk2r2FJpYbkfaXeW1Wzf2rA7MGMyMp2W/yg2zF1Hj0TiIH5XEBFzAlbH/LnCtGQ5
vNQMciOp6SKNhK6z71UoZ9ZvF3fPqoSI5t2ScyTv0h5RdUCOxYeK3Fyuf7FSiBdCQyv7Te4sKJ+8
rXOJ19IqW5ruY1PXAEtrBstv498LZ6NRzZJgbyN1RyT/M15laaj3MOjkPucICB0613RmQ+2G3ytm
wSwKT8qpKnkFyOfrrQ+9hJQv2yJJ5vcFHSls97+fyb5nRodJbL+RFFFiitmGJh2Yhxu7YVJLFB6Z
fl6xP3zG7GRvhXj3H/8jVH73UYsHn+JvdAC5WzneA1dM46Zy1UGMXkKLcqQjrYnbALLx1mMws4RO
y/k74yfqV2SHTYJashY8RbYu1JBddVDPZEmLJQpNwxBFIKSMRUM5nYZ1QP09ne1E2cKFWpP46WWZ
nl7RXE4NMWceXbulwhq8ugOH6+IHn1H2tCe0jb6gFj+v0me51Xv609/HA4rRoLiMhxZPMncs3Ef/
/rSVhd3QJXXJckGz0n9318pTzbilKswuzlYaxDaYHoZSxKcfFAIOFp6H1fMcrEozeUlG3A0sybz5
+m35eEvEJyxsARa5n7k08SQ8YnKK0apk+CHJ9qoWKBx/S2NmqcW/08ANEyj+N2E5G+dEShmwhkLn
wfnlNWufGIIThyeqnwsKXQkmCD7BNIECz1HE4PqWSwNCJ8h5aLNDKtsD6PLPUZyDKPelRkNK2T9f
kVjSx8QRii7jFjXri33O6DG0+TIWyh5zimQyQ8DLwAFDWQotDBXDyKzp+4B9XwI3PoHlkfPMcnvP
fLBEMEwxc/+Z6d2t2PSitgOf4cA3MfSWCVknPAonDlufHLP9otE5JE63QqpMcV6bQewLzlVXLhhv
tOBT0+fpKjBSpF7DzuMF3shHLmrifJ9JUuxWOZy29PebxMeTua56giT1o91vyJSY0IkDfQyMYGO+
fL1fFOTPclRh3lAvvz8L3eyXfda00SMbyN/eQDYmBXlClsT091R8qweRTwa/5tzPLufIlTp8JDpp
+pkPWxNytXNvcaOxXGuh6GEyFM1XwSekogzM0XKdTqfndo6WjzDHFeFhdoCI1eTBcrncpHXPa476
HRj+URmgzmmPYSI43k+JpeBPeMTXFIYXX4qwZyahU8QJymnM5tm2NGJqmCabtDpTCf/kzM7mR0at
0h4YLfv1+Kt9tAN5VAn3g4324ZN6Ant4gD+7toStsOnXWiW6iL7msAvceJ96tuV5Wz9hUphcUeWm
IvjpoH6tDYt21S+5JDYBg2O2KePKVc90A3m+Gtt8SdhmOZJLRbOuvA4hwx5j7CxJuore3r6as8m1
eJKl8+MtopgDURCtI7S8xnFRji2zF7hZ0kiWm3AOib0GCzCEpSbAT0qjuFwvtVxLIqDcyw9FWRWC
LSe6ftLFCGt6U0gnXEFGTGcfA5q8RjdZX71Wa5uK/CwsU8pTwFer5vk+cKOUszKbe8JGMqJlv3ML
ht8aIjgPLsr3HwFSazez/vuh3slZywg7D0JlPCRM5Dza8W3tDNNsv4L+BIPft1dgmAaZ1sqyoWiA
fVi1SQAYQBhgtim0oCE1jnhFu396Qr58Un9TcYx7oWo+FbvrD4E5kkKF7H4ufJvO7UIVfe9csoIG
Wj3goFQRwR5ASMv7UIpF1tv2JtpFGSpGk7CNyalR4OmZaHxl4CA+2WNzoUDBTLnV+P6qNjLRSsr8
uqRLPUlMzzpW/5h8kUklAprg93mYmWPa4uY7zBVVL/aIiBQAG4ktXVBECe+hDNuItLaJ7eZXmNDA
bnL08MJJKddmEhIhrMlgeFyF1StxfJHgbUaq+4FOiGVwgqqbjVyQKaXV4CQfkai+feXCKAzUpP0n
lrDCq3sakjkB9gsgo9zreETTydev+n5XrGFkLDftCmyZAjInfyO5JLLy9aE+kJgpQezJckg8WazL
e09aB1uOgDTg4gJQIMIgjnLgiZZ8xBOi8610SD+vOQa3K4zMbq7GccUEEUBs77AioDrNIy3P389N
5HH14wRIP5B0p6+gVfkZvCDP6qwIoZ4WxWRk3w5whYijrRe1yYNDGAcGy9oaQpwRBVYWjJ04XVCD
W86jgGrjoM9ndpg+Ed3yL3xvDHbxaj25NW2uXCwu8zYpw4Yjxk7RnCnJFXmD24e3HKxyCUm/JvBS
J79pIgouRdiQ/cnzYCMBdzLnlwyWF2B3wD83E90eCtjEyRM7ndjQlM+a4Sy9Q087e85yxuxIMI63
Bs24k+B00DsXKXQcR0SVNzItjavhk4BuPAwY8L8+VtIUr17zL+asPeAw7G7SpJ4zGgPAUFdz+MUG
V/0SYvMkET0cWrcjMHva8A0u5Tt4j8BWVUv9znjBBpuqKCKOp1Gbmr/oImL9JNXHkbglqjKc64I/
+m6Ntf20ArNIApWC0Uaa6Xm3vyXNmWeomuRkybjk+Z9YSej4vylhEIOpBp89SSMql9vj0sTxTjga
DbJOrekoZIsftRG6A/XsJEGV1a6jPJa3TerwYpe+XWsN7siXqKboT69GTGxZe1Io0rkawJ86Un4M
lT4CejCeIT9RB8PaGDmWQ8+0zECglBrHhq3uCOFjxMPL8kbDK7/w6GrxMUOdvhQUvFRzz1mNHBLS
7ZOlzmKkA1KOPT1nNZVPk5PN/KaJBPRE/lVxOsiotg9x96WD+dEgwyB4q3HlnwqRvxP05B8lKqfo
t2d9irGWXUJ6j/1X0XhFk+Q20i0o0bgySVugdht6VTgAnEoRlZlTFfjfyAAX46wBCxnnW08LKWZv
tQQrZbIyL3jnaQKzX0s7xnYIc31OzPm4iTimO9764Pxrjb0z7W1LmsQHCY8QoWqZnAclC7SVs3uR
ivuYnFs7hdTK5BZEwkfpre8YmgoGllR/V13/xkfOMhrX72kB3bDvHsVD1PZotqsco526ciWafcEf
cAH2+cWWIsR8uwoS/zz22bf7EvHnOvB1rhvhjwVIMHVwUA2dXfgxO0PqQ7e/0K5ZE98qmWkF0INh
VJ0AG71ROCsTi7zcEvz/XnUKTl6/fSQRHUxLWQqNwYUq4fZj2nAz2fZoH6/vxB3S2xtxQ2ZKFKCJ
eYx0Yftic5/3EVu/BJbOW1MnFYhp2nHNtrCCjfP3+UePTjTxXQJZ3NGa3MKYI4G6w4cWog2gkst1
fh7dBv4RrD2DX50acP+bT7dEF3SObtb8vrFVAy/m1HYZiLyVHuts7K8rVjqgqsB3cRxhKz8J63R8
A6NGNHuAEdS3mv3vEEQLraJGRf5GrLHc9ffYFpmFyIK8UAiSG8eNrhA5u3rIVjb1AabZGTIvUpeB
SqWuM+eqiplB0QQPYH5Sir8Xug3tv4aWFVFOFyRChh6UGbYarVruzx069KMz0htyRNT2+w4/xRHP
09WOU3hsMUO5d0Exb7jNUSqHsPejCG1j3yRf7lTqQzO+oI1OFk71AVy7ytgUb0Kzwkg/pXdCkJXt
TJz3gLk1/Dm50wyFKH6JdKaPjlU6wNrXY6q17hLqdRksttrHQFsg6kfGVX4wd1VVk/Cdn8CSx6YJ
fOoiigpOFq4yguqfzM5KJn+ysmdQWCRAwBGxPhMvXbyv4eiysz4WdI61fuOXtxh0LcdnksGr+JkH
eaVPZR1uAbweOYnq/Tznc9yxf8v0vy9q615gmNPLCxWUF92YADhcuNNhtssiVxdgTcSPjNng9MZw
X5mExjo9hoIBTE5Wz4pyuppZJ3CuagLFGmAOnFU0VqhqX2do0IWRRAVnKBUAiqNCTgS4ixa0bhB2
k/Cril2A7CiRIi57Hdm81qwOzbYNPsEOn+APAEhSDD7kordObjUl/dtE8cXhcKY+5Mb1iWuPDFY1
ddGe+3eEXqrcEjAzKt8rvj9c+0E0iUhxZslczFgnACNN+zqMekua2nSPPv1yb/PSvq0qtWjQZhvX
Rjsf9XqZ1KC3nLex/UbSCVCnOqPuWDXNMJX1BI7VL4IM5FGtRXhvE65/iOWA+gwsHimuyxllWPsc
rMfU0UEA3pmfWWmy49/IVqgfchdBHj7/WrPWXCR8TQv3l17YsEirM0Nd+K8cbEKBjC5CEEH32vaz
bQtBCkYLf33DYfWgdFYblavSEeBjy9O3tM8TbVmkLVpmn0/0Op65CSGlW8zkQls1+myJxE9o8HJH
zHlLNHXDPRpgPm1WYeI7Kk9Gh3XTYuVJ2NWW/VLSTN1cwck00qT/rHtEeE1znMRs+CUBH2Z+QSwZ
mCbCJoXg93AYcBvhntyq8EIU5S7VpLKG5Mcbr8FU285E60F6lLoaxRgnrT5qbInp0slM2Uq5Vm3p
qre85O87tTHEyASV0P0wkXqcF2ZUrsfa6YtzuzvyiUa8NoUDUP6atAKOYN+0NRVeGqcfngsKojV0
5FkSQv5UPqZrY7vaeY3STg3DrF8024oFuqaYJ9ICJUdhgZSg8ITx4VADTIlYYv4PI2S8czAX0DMU
Ft9IsUckyLSxvsJ/5nZUqzfxaa3P0tnrZ1z3JBwfNKRuMwFFpGvjF7GaI4kHspm3ZeFKajxhXQ7Y
3NUYu/mX9WGEiM81PrAPB7DdX/8nv3/3raUVtGgEW2LjrZ4oyZvh1vY0MjWC2QD2iALCt0eSIRAi
6fB9hQCyCPgwKKhuzYGJCGPgyYNt3LHgfEiA3CauHnULvmj9XTMUTuc4Op4hbnkbRcfXy6j5VCVC
Z/y+tX7yXmr27k/0c+kzWnT2MOQYFqDKdIJnNceYlOWFIugaBPXIh34e0xxoG+iWgh9ztkXklFFi
fI5yeY6CSKQCwPOnVKETnSJED/0+tqBG5I/t7Y4ATQ40sMSkSpRp8dCk5E9HqnJdL1n1ZEx0UDrF
xW/2xwBQbxwNGj9ivSTLQ6nxBgKPZ+ptZDTYbTz1kJc6XGQf7Ag+RdFsogw5HA2BI9eX2q/j1n5X
nRhtJukKEGGZOIAfhBpxIhmXh+D2fZdmUWrbi3YvsRvXIoVExl+MyXLCtVA01EZjr7seD46Eq9Wr
6oLXSXSb6tB5w6d4G+er9bypkYLaqQfJcDivG0M1CAEugHHhv2vx1ZrnJ34+Py38lorUtyWGr83v
Nbcxsxa/DV9/1QfECdP5N+lPyPTqj+ZcihFiHxeP9FwPkBKAZp0RUN0P87fialEJsaXWgHUds88j
cMUkArWYWS6sNV2APfRPDDUJiSlzHjo9DShYapPhP2vGULahKwWDdo99PiIsMLMenKWgK8MTy/0g
zew/W07q9uMk654G7Kop7flbyZzSakx2u8u8E43EVt/NTw9C8gFaKJ+mifz0ieFIrgMy2YdfGcbV
S/5OBMXPOUcFumz67gxaF4rbY5c4Pf7jZRAkv1+d0GJYBB4Sh5ZAWpTc/drFhY7OcxF+NsNBc/qf
trNgtO0V4xga01eJW+tTEKsrLBayrtz28fETQZuKv2b8FQc4uWQAI1M4YsZ6N8MZn4sWEo0NBDZ8
89xqs4HHENHFrtcAdIU3dqmYzrdIegtOPCaBol3xWpMVjl/CGlDi//85uqAGfzzpL9h7yS2WrpTz
OIZGSz1q+RTqISTcrwYED9e75nfwLWwVKN3cJ0gBJYtO3MO0GTC98Y87ApEx3o+7g8wx535+oRRd
+h/JJ+J5GbWgpBLxcb3RiTd3Uy0t/vJaRHXz3IzY7j70q09Bh4Std6q+WM+6W1uWmDQ00eK2HZK8
cHoFNMON+MJjt458ErRSzL7HXlLdQD382WTi4SKwKi4E+eFaagEugNUcNGAbMaxYnLVu7IkDzTgJ
3utD1FJWb4UxqLuXLPUgWgP/2tRGqZn/WKYjfjNNG7HJReL1NMz3pPcJK1JvZkDoN8GfWj5cUZJu
lqkfLPOXMrr/QT41Q9d4u1K52Cj5QEfumXftY2fUBGkRUfo60tbFRy4HNhFlV6jdo8oXrCle1N4p
EGnNvYT8GswbuntN3DU/Vu1NtRetNWNu98Id+2prihTp9kOhCXRReGdnUf4WFSaD2kbyqWbdGi4r
NTAwpjIlmq83TK0xPUoYQsil+iosiwt3AR0b8r8b13+6vfszsxNjA2XxsMfkQUlvmVufenXQZnEX
b053kOKmVr6FlJc94EmAupH2FLYG2CB+luN+pXQdl3Wl11HABNA1OoNHN2BfjkReoXpLfWwKIJh+
ly9hN9q41/ZgUOG6lZ54mv7kvIAd2rWDWxdLItbEKyQPqLYWb7/XXHevglR7J8qD84HOhTr87khU
mn61VByAumxrKNX0F6jyz8tmbmpAYm49xr5NIbOkbWzmTY9CW94mDcTPkjHFsYNmIb2ABtvXdYxN
loG9yfHlcPtttAjN4iIpJHpZ3xvkDAbgZGC7JDlZyOWApK2ciwbcwEXaV+GUdU4zR2V2JRJHuoQR
RshFtVLekE9Cwy0DpgqqwNEX46TpC4VBoOBsZ58YFQRfZRxuIL51AUgKDLLTXzdkjSJiK3qEBR0k
DmeOgNR2O8d8mmDAdLZBT8c4jFPjSfegeom+RpT0wsPreW/Q2tC4NQzKNwKrrasOwqvwpTl8GyjJ
7zGXM//sJliXuW5oH2FaKL8GHUchD9hFBPZIkqgi8dtJqEJHM0xPcDsVAC8bUyddx1qZJK6Y/r1q
zXNOM5WHEkgV/IrEClJWVPCLE3fBDuBKx+3l0IqN2/iPJSYgTJIIsh5AFajzkX+uSOMmQrqGhXn1
K00LxvXWua7V24DWTxfWrv0SnLI+41HQUrcpALkbjFz+yOY2Jw7Bxx4o2w9wG0cUtIAyQYJGNGvW
fQFpbs0GgESakdyeX/HbYeNDFHUcQrdp72MkCL45HxaoQ7e/c5AHl9AuZ14AMu8N//N9LMnmaJQO
z83hru8z+HLo4yblp1npAO/Uz75ED7xKDR5kYnozOPXQjwte5xVLv6vW1R2YPaOmfdbjgAzU+k9p
PsBoJ+R3Vrq7A9sMmEaqqAp5n5Ovf6T9gX143jhcpztfX+VcDjoauo4jBiib+y143ACDQ3f1fOdz
fgikz+BgmUgUd1tgQc9yMQVWmAAcFlvHteo7uHWMYdkW4kPX4/IdUKnCj/jid1EOqB5kKIMRfnHR
8HGSWjXyhW4X54eeB3SnYrrygr3w5z3REjH05bmDyhu53IAJaJpOotiIEgVYCKami4mxoAJkKWJ0
C2nB0MEO25O89mnH4uLu8Z9+B9F/dWhb08NeS7gi5RP0pB/TIee67vUhwo5QmJH09Kc62ge2KMYm
SZc2oNz5MIEgtUTWphI7CHxAnwevomtVbSY3WxEr2kz69MwVMKb24LDiOOgeTrUsrJ69fYS9wqgj
5EKOVP0Kgb5DRM90cbF0L44JrgiMCTC04u1HFiRzg/W2k01d8OdjUVoVbRbFLWze9lr8WbbPAGCo
3gqvjgWp8pFZ8mmniZ8Ry5khjlYvh0mQGyA4KSfKtr8wV9SUiD/CdYiYYfWUSOvKQyQBCQDtVN7F
og2+EBvPHNDg4HKloW8B5w0jXklPomNTU3ssrxh28J0Kxk/xN3kYQjitS8JO4DbDEwned8yCkFJm
fAk92E1PBaQbpDP+fYhlD3m61OgqFW9zAu3V1bwuI3iMi95K86jW4CI3BaRrSEXBMvMnvkx8JPGb
0hR623F4V8PsMr2YZc1lVk4ImCEy0l5I0Q7xW++Y4+dh4dg0Cnu8bh9kJIRgJOUXLzQTreTTodS9
crUE0r5rXeJLggzCCyDD2bN3oPlKWRtSR32zqzQloCXq+1OeLruK5esZqZpr8DaHkmzzDxWwepRw
0y0SreZgEB+Ya5Rc5RhWkf/sfibdZjJt9l7vS9CiYlBYW+4o03MOZyCk8+Sb7Q0ZMxIrAHthWAHk
SUkc43KksZJojMl5Uv+DKpXjTDbCMdA/DZGKn/Wpt6qLP87VuS1mHS1Bgzv8c7jEjkdp4XaHYl1t
2F0mbeR8Eqpex1t+HGyAeOoJkQBsUOmaOA0AKxhs9ulVECAoqh6DQ+klcGaNUjd6S+F71ZWtXi2E
jenN5wDYLZpH9rJEtrpYvicWfQ3UCxR+Dzz+rJnMew8HyjoBu4JA28xdCJFcCubfHMo1gTLND7zr
+v2IwsIuUiQPfaAdXSupeS2yktWbIpxXvWM4ivccOH/ERWL3yo6CB5AzQDD/AQniD6LSEc7b36WN
xasXRrSRP6Txx4OhdnLf8Qiex+EvmnyXYOHk7LZbl35QFuxGX3ysV+V9LjeKAjQ9Q6n1sGBLaD/i
lqJOXMzHDINxrHgbQu68nZE/L+MDrN4LsJ3H4S8ZiqvXqSDAVU9pU3J0SQMID4I1hlu5PwbkFIh5
P5Camx7iUHxVYjw4hlknoo2w/vqw7Ope6u7dI4iq2GlFMiRn/k+8fYG9RSukBJRka5VRTDSEZRnJ
Ruw0VSSOCYPLosVH62XD/+ri+eXT9xGvne3cO5zLF/cnWkG7eQGHp/HNLmEtrOS+De4zRKu1id+k
MJP8tLf3wVP6zM42D4URglw4BgeakRyuiOp1BOYgOwQL1Dz13tJMIdwS+bb4oezdde9M8sFT7Yzz
fb1OK3PQK/1DrOS5i4GBK5LeBKgfjKiq/XSJquwDvg/bfQZ3BoshGMpiUWd74Z96UeJ/nLM+kJvQ
5nKEWdSdUD1hoBt+l5Q60b05OZypw57voh7iCSLDMCzeBwzviS8RyuJZcalUb6b9dLqIbZV2B86B
ldlgjMr9aoRRrHB2kuowY6J0JT8U6YLgB/LgiwDbV6xNhezdew8ZWiiHajBjW9mJBUtUDy50Agjc
gybQdgl5bGR+e6dPbBhuk8XNq3liR+mQ7dl0LbgNcq1WJ8ThT1cIpxEUJEZKnnlnfzHC0UBkZPzD
d+pNDKvfSl8cstEHC0cCFQvLmN7J6AoGRnbEc431Jc8N05kcyFLby+z4LQq6f+0eeoeZ0/CaWqvs
EQ/RSZ3MF8COvRzQ5mwBVv5DcbG/KaJCXgQqVFqoG/fDWlYxUhZo9O/149mrVX/VClqj8AE8ZVf4
Mifq7nVKsp8k3PQ3vkVzmlLuAGufadv/ZfQS6Egxr9BhC249VBtATwoMyicr0kv+yNV4KJhwzBu2
zQ1hJjcc8jfCAF7qY169gVQq0xAambfkM428bDd8JMJY3UVYRakkSH9gWacZjtize+VA2uBSwhSH
UUodHNlYud7lOcXmpvZiy/ojDDcyeZnAvjfLjyjPzB6zeN+WkqjBRmt38xbXDwuIDXAi76SNvX6y
jxJk9BpxAVioOF2vLI2LnLfDKjPyMCHBMopypQtAtc00mKbO/AhP3y8b7fkOFmOmO4tOiIPE6IRj
PXtp9Z/rqT+bfNbAtdExN/FhvzlILrpesogrgzacUxmrm0NUXEo3iF+6u9G1nY+A0Vd+U9miVxXl
6ijcbCO1zrzi2iZsfaFwU0yYMdxktpW3ngXVk3kI0mZom7raP1JFusOdeWrJSU9701IVNan0i+Kx
ggiVd+5/zjcDGuqQQoiWNKEtGJ17Hj1ZuadIjQk8fCQstQ7TqCL9Q9hA7ScqYjxbAH0Az6xnpPKB
gMEzQhGEapt/1D1xPPe+kdyYJJOLdA/JjmKGGAcE/5e4tM543OWvCtMsVO0j0f/m8QkR9e4bb3CT
syMHAyM8BElsWGuimDJkHYOd8wtFx5nnvvxmFww6Zhv6s91oYMNdiUIU1+3zgHyIhrcoMj6nsHb1
iCrryJrHHQU6UmWDoThFlDWhk5ckLpxrY1CMc7eLO4XdFVj16zepDCjWqb9J9NIXxBn2eW4+IUFB
+awx0aMrtXpD+Rmx2FLmC+DQ4ZcvNjBxdX48DMkEun2vIimmAdNeqgutV1KbLjxMUzv/ejIX8+ua
Q4NmrJVbwg5/KHRe+cVHY/aPBmEVSjrkp6aivCgNVETo2GE/+as892LYanr8gc/A85+Eerkkwe6k
71wT2FyDMoD3cV4EnPFK9Fe1S9F637pUYei4gE41j76ls1cY+VLEmLapvmVASj4Ca8svZ375rd1J
bXTQnh+iMe4hZd2S+v2g6FrvWs2aNhlQCARd6aPv+2bD9AEYe4TKHa+L9Z66qzsSMbwXHyXlIHkB
/P5DuOiGVZ2xaoUiMVPaQ4m9nCvxb/YVKl5m5zRl+r5cvi5iqE1xKApPOlbPR/Vu68jI/HbQYaT3
4xTr+2AYYiGIzjYV5njMx4O+tj6k+dzUBkzTacIO5k7tr3oX9kAiVZH18jHUhamIW2T8MZVg8tNd
venk+fwHvIYEKxOJYmsucGOxbTe5ZI7CB36owdUiJsl0oAJ069WCzX5opwnSviZdpn28Ajo9vI3O
ZNjq2OeKpLp1HCJPJfeseu0LWifma0rmV1wjunZNl3vBVIwhYYO1rKXQvZEVqotvZeTi9O8G8wE4
DyfM6t+Pv6fOe44U+kSKGr6QrYHPBG1gZaBOjYyVLCg5BD/y5Xq/lJytt1kHeG3jKGIiU82WnWTn
rOx2rlL6ERztqj7GjB+9y8x+FhgtSc7FrcP8fvtSQqrJJFeOUHaar8x9Z793OFN7krOFUGdPHnOh
smpuVOBnHdr3pnpjQyFl+zHgZ3hScrb/y9ZHCbeN3Gl9KFzmDwgCcnPklgwVLX4r3mtHxCK3Qozk
wceACpjSdBoX/wsEhz0Axc+3ncskqJDQnN/wtzJG8vJZlSFVOstiJQfH6vCnaFWNThbdgGoYpfsO
qHa34pH8Cf2XHC+M1bWvwJ+aGs0oWUEsIVG/HtAf4viNA/r/dKQA/KqX3DG0E1iGoh46/Z8VOgV4
dUPZ0q6An/Xz74H/yTLI0h+ulDLwU5Zqj0nBkJrzZsM2NCddcnvzho//dGiqP72IS35PbvFWeCIh
Hrj5FsKwuhkKNV8CULtnYqkPr9cr45e/hk0jrRg+PTeuKIBINMsGHEJqzI8n022OIGNdlmWxJZnb
uBXwBPlz2mYiLDn3+/4foeGHvqAFk1nlGJBV5BVt76Q11TV0K41T4QbgEnRZIU7GiEeYZPc3dZPi
8mitNVdtPQaQoh2Ga65lNIWjDleF7DSzHd66zzq2AdHCde4JptQ+Mnqj+Wug7jv1dl4L+obgqM2g
h2pIZQZV4Kp10+fNZo8pX/62PtiF/odb98oPkilUpS7Tctx0EnbbdQG2qHQCStiSVA/hQZ+qmPpg
K7FxFD/WwqTElz7oVEFnrbx5+HR62jy96Hq7wUj6XxeZx+DsKOxZ5TRLLjVRFxTIpG09yIIQ6llz
Fr+ZI+pZV+o3AS4ZiaUeS9/Gmf9vj9IOZWFvabIQj1jEp3Zwd5EEWatDsOnIxFAvm0GiybhjiPrE
bdYqZHiGKaBep5Jbv5Atp6RCKcaP2C2IPx0iMkp3se+VdwtGIyW98n+UwI4KrCAOZN6j1UbupT2q
ZSAwiXGi7j5qSWsZp8dV/stldbs2YMzN5ity5OB4aenip5NvZn/eQUJFbCOfZ44G13znzbhG3vI7
kK+SR63A9XJuMhYyQIib+NZXSVcuky0lDfOUMLYekPc2fFDK6lxQY+rxkY6pqjFmsjHW8RagsRqW
zafC74LmMOjbF3R+2hodPDjeC4TPLj2nChjJltRQgIAY4f9JwPNp+ZyzISF8GPB8HOW2vQkwcC2y
Oyy6T85/dChArJngjfnEYE+z+yn3zuRjZiDc9aFF+igMZALt6r2+KzV+FdkZOUVCiV2k/8gklYEB
gUAzXOaN6a0o0MmOIsNeniL2nYIPeWOezcaTPwi1/fXfAuPn1NmoEqm08eJp6456wj5wW0JTXijc
bf/uCcMeFjSfbvfr3ibQ1+y5Qh4WV+VUXDYoxDGkxNBOfJwRGdAWSq+xrCegYVV2G6d7MEL2ZaD7
n8Qf7AnaaFAsQau19eUiiWHmQa9MKYe6lOmUQ5pwBr2lOFarTeeO66Yl+YhIGN4sF+ih7jJ8mlBe
rEII0hgJyPLGBiSU90bq8tG2n3H/rRnNfhImDjwmSBss90+utrlaldlAVdNp3Wdb+54AdC+th35z
73M2W9v5LH1QLqCGccXBux7O9APEwyUzSgl4L5lHJC188CJnP0iokKCa+f8eFHw0SNadPd8ky3W7
ZcCwABcn3dTvOA/YQislxCLAP8OREisiuRFlZgR54AX6QU3bZoytbfJaLDFU7259MFJvsbBVVUSW
fB1aCRvD9sX6P+ATz/iPDuS6PYTScbNr8PYD8oKKGF8GAlH16zB/AtGCTjIu1nfbgbMd7U4XivDP
zBz0WS9YQiD7lRXlTuJqFnt6Xh4bAsUINdRzERDl3msLq3mQSSG+bq0Ru9DAXKGc7SoRAjt0t+wo
KdebM1Q78WpnYsleXo3v7Gg2aDr/5eezy1zFeY7eeacAt2MRn1M2/PT1jtdf7LQI8wl2Z1tXl0Nn
/krHw+TuMh3ntR7MheUj3W8h69xHSqybeg5r30W/g2UAp/3FQlc3Eurmz7IbUa9oRdt2PZjZzgE8
rowaccGjCYIlK3++DUf0YVIBGy8QYAtwiPgZL02j/1JHvzFijcoyS6Li7sgRfabJUeuz5jlcA2U2
NjVu+nQRjd4CKwdjMvYTjhHEpLHiBdVNl+phXpaFCG2GX1c939xTxZrPKObEwvND51KDlmMw2Fs6
bfZAzsGT50Q3850SRkv2F1fif8JxOfbawSKbw3CqMZDSuR0TXD4JF4znOYx2ckqe70u8yjfl2GjF
8+spXBW+KtN4SaqE6KkvDKFj9doVfSOJsS1YDHAq9AtUEKRXcOfaYMwiA1UNiGvdKkhEu/YEzh41
MWF6xMtJc6DTX7Kcyq6wBvs37vigYLFfOhX7t1S/vpVChEx9q2LbTDQ7HVaMLQLWtvzdxP+Pyfn+
RzEHy2zDq3wjp4GeV0YdCtTppoz/yJXJIboU0+WeQ2KKTbNtzwKoZyrYmCTQUaDxUf9RB6a+atGN
cIUlJ/qh8p2rY6L7bQaFqSdbIm6rAi9Z+Zi8pxt9Q+4n7/6vZkEfzTzl3jKtC493K69Dcx9YJdlW
JJXd181uUmm/K+Gl/af7xqXiYz9xNyUdLHxy6tANkQyDeWeFB3MLuH5swP1fKOWwkR/IH8O7RqFx
bndIeyRDDCyAOS0KvTN/HYVz4bWdprOvz19NpJ3rJTbFxiH3R7zu10Hug3nNEoW/l0ta4DTS5nhf
7yjSWlNqpGBuEORiuQLrVKxuQzBFKAJT121VgEdjQx8NovV9qdUBGNBItdqfxapaB+Golmqk2f6J
3inmOfnMxNKWn5LGpz9JNasbQIPhM9KCqXW57Lzhg58b+MS8EThuCor4VaAd/SyriR/FMaB9rBFh
z0L1ufAmqZFXtqfJAmeJJZIlMwk75EhiM07bitHB6wh3uaW+HvAs9N26vQM8uU7edAemz8gKvw27
rQkRYNfp7Kva/pxsd9aT7Cf4nADr68KmeGNcW7y1ZOhGg3DTghf7QFjtIRxovWk8/FWrqNS8RpX9
Eftxww4a5W1P/db8wy4TbZKRUVcibLoRYu75aMoQ1gNu9QX5SLf04Cd6IazSXsZb3CtnIo0VRatK
SRDTKGDXBme5d6HHFjOd86fAhFq3FLU6VgJ0Rx/c0XM1q9fXesTr9uXa3GmK7/+49TJp4zXXEuAx
Ga6EJ9OVvPUWjjrOEWxyPoLvEBbt2qWmf2OeEbzUiWeWiBbcW6vLge3lKHDcqSmCvZ9W96axEBDt
xq5whb4y9bmpEpcWYLQmc9QXQFWBccCII07XLzzC6CZJnAZ7jexohP4eEQxdBc2r6ucdVxuCJQ5g
rjhgABUVAwmetS22Ic2WTv67S8XlQbrSiLJfzK7Wt4eQoI/hA2MrQXHCVGv6HyH3qehcYLdh2B2h
+0NPtBxoFtxgMVnn2xTQd6GPHkdF9PMEXLK/ZuxGS1JRvlubZq1YzV6/p6IeAu4MMDUEh0/0ewxX
pMRcoys/PzTrk7LCjyEz1JgSc+XUxO3L/T4xASzLLMQoRQoxa+jLaDN37C/n1FWncpPHzklwchwJ
mT+TgHiTVC/Kmnifb+ML4u1ZulTSEjS7ONAd9/zIc/bYc8+g7B/QHS8AsoQEpbxgTYTtfSevkFxA
ogp8W/cuU0BgDDZmFSAl2xCtrCWWsiTjYzfmzQIWD9XbqDjgcVj3UgYr+sbm0Mo89k2ESyu5wpLJ
rMykyeoyl852YyYIOje13f55Z4r8BX8XuFF+6kHRn+/Ic5OTwH6ytPAHHS7/gMlYheMzEWZn3E5j
mwxppyPAj5L6kKSvLD9E2gBJ9P9c4nTrBWd01LOxEdRW3ybZ/gOM7hC4CSH5RMg2CKJzd9PH/Lri
rQ1OdKyt+pRq6Wo9fMkDtY6xai7TLgkDmHJJ/DZnyQ8J99JAasjzvWM99YK0DpM/Ar5i+bHXcaBk
q/lgc4oKhNPIh44swvZTZVfi+GrAhQsiGGfThrleY/Sg7Qo/ZT0gDa8xcwYcUH3KaZ5FAYNW+qc/
26s4Kq2BSNFpJTUiYacHUL22l4/Fxm6lD57J1S04nP02l8p45jPa9AWHaQHgJIqUxZl6hKsy+u+q
7EiOAMSbhDsbJXmRsnDNRx5SVpLiyZw+xta72ZDZuNm7t4UHg1pXEiPlItu05+t3poWWyTjAFdjp
4AGCmn03RwXti0e+Fg2XYB7LQoyrXEx7PBWMek/oCxozSCvfPb3kk2aa/60A16ZpT72m5wbP9/s+
TfMemFz61c92JmO/21kNWu8Bkl3nU9BvIQQFTeDROpKMJ5B0IHq5EBP0WyUWbxTbqp/2iyKjdCZc
XEr8jMHztO4Kv2E5cRzuHAM2A+6o+cMdNio+g/t2idHH/FuWbT2SXKQ/mOguaLRyLdykTOzQsLGQ
NeCKMO6HL8uiTbDcpDiHgc6O5qcsgr/LixeOp7KUjuesNAjaT7rgds5S0UmPfQPQ905dngvhAKyJ
OAZUP5uvx1x2je0udXjOCggyF71pPsfJlGuDNBFi1vETK6uQlcv1deDdOiFKSFJablzI2pxw5h8n
QgGcOYrO9/hkKKwiQJXeoNoDzDiODh97GecGpiDUpRfCtay+OjsJVij/+RXoJV59TWH9WnzJdcAW
zZFtiFaSqQ/BXfT09HsXHpMKAg/pJspACrdTDUv+ZaW64eWDci1/x4z0AuExADvmkmYM9UPAwmWl
36HqBOTazMHHWXNSYHZ0t1sQfY90hgpkUGZ+6+hmja75MY6SQvrjXo7JwHVvJOkx9wSRLld+ir+C
EjoiCKKIvih/RLkTUBETcsahOUG7eiTQiYIv8qJg2jSCtr/EjWfJ8lWnB9RQekgXeG5rcqvh5z9C
UJJuee7eNJu38wp3MlRjYdm8NEsmTevOSC0OwpbkbbaXfGfO8mNK1N+YMXbcbXXKcGJSHpVBewtQ
3eM82YmEi3DdTmioFTmDqxISkR01xERcJ5zm5I5sE6aM3yeBhyQE1KNMAMfxTFBIdr5H03kMZMEE
JV9gfRUKgFKoV3wWizFKNBf9wH/NpLQq8iqhkcHrqfUD8tAPQZFWruOXOuXWIOAPGf5jgXfSVCUE
DrO0/64ZbW3xm4EXr9A1q2H7MTz7GeXg0JljcRBTozlLQCDP8ksXRcgeSdlQ2GqShny7oBVIXYVw
LsTyvpiqaBluo5K/qozaEeO5T2+YyNuDA5x3XUK7Ga57q8ldhV1dynN953xHl63Sq28URoX45YaE
XS8rKMt+9CfrWMN6+F90ZywIzawD2l6moTvEPVwi8mtmMhov6xGVm2i2x9OJtMFWgzMBRf/kI28c
0tFsvw/Vs6nBVpoFseWrIOxRKjuVbCjaL1+HVHjseLqso/jwk0PDCl3qoc7CTHV45b5kEzzfPl/S
TIbkRgL5zZVPiacpb+GrnTJhTAXe9ZTA/LZCt/H2RmXmBfgR0vYaiCUfwBju4PBSB7zVU9AwDe2+
K5eejhIP0lVu6BuaTeXVHebQ4Afi9jDqCeY557dc/n8Cfo/E4NPY9P9vfLbNKzFXqrMCruUV5Owb
OgqzGh0zB0w7gQE/msnTqakwlA78QUf6H93TdZrZ9wexoeelKL/jIHdLYDyENAs3e+UlsnJBHmTi
O/MvBW1N8vC4EVjQUOQh07suA+7xwO9MI12+M4r6g3MsJyv1XvGp0tU536/JOWDpb4rtD8HJ1kYs
5t8On6bmXXMRuyOvqi7wcnE9XHjFlimcrrVvKvQdkYenu36vu46gwmeoFNYVV0RXFOv5maEW6ACM
hHhJcO+puefJubcTI4tngGiEf8HF8QQGze5xQoyflWU3Q877S4tQ82ZVlznDj/YEcz2ytwZCrn0x
ApEJsK64FHI9N/xegpzs1N/guPUyXOT0jOzdZDGQtRoARLRNrLofuXSLgpDdpOoRw5acmtlffj/o
2d4u0PyWtcSCfqLxm18PYCHY9TM+cqDrCtrxUepHi2hebgPYy8Zv6xg15v/Szs0B20papdhjjkNR
GYy5k1IyURATYnFfbly3mhlyEsC79B6bqUOKcOsBwl6yswkLF14tOoJGDugSPAzf3ULZTZgYOg21
Qu2/lwS2ItdmpgmYODbFG9m1yIsAe82Q8cW+MwyWHsr5q0DlsShY6rcDHzQmbZf1ipp+n1UQcwdV
VKaGwUFgA+E4n38vhURD+5/LXgY5qstGRTGombx+mz4r4eQmAGF/p7Q5bS6JDxCJFh97lJM3BvCn
vGxG90GzJf/kUEQSZvoMvOpfBomFX3MT0l6766tDhdZ92uDechS5+7y7CKnpscbM8dRS6mkbZ4Bq
ZStitjbjtweLSYPpd91z0oCOXoNqhl2pvDoaatUTo3HM35Uz1ojQOekmh+z1XfH/QOqwRtzj6h4i
MaJAG7rGsOXOt4YgwjyJTzYjmroA4YHcrihoVCRYDbWkvYJJ2My2be3NibZhtaN9/Q+GvF2jFTuk
i/gXTpFvelL/LsX3OKlCR2DfhhTau9Ad6SgCyB9jczBba8NqWgoORypCBfjB9RLzCaOXRVKE5gVA
I+i/BFE/f7uIjTUHMesUxQuwJhRxjYMiABq/YlmrHND1eVYKlHcmNUZItLXGg/gB/Ww0tJFXRLxD
Y5j3WhyMRCz1OscoadnKRVe02mCUQgqgYR5T9rvCeN6mAUOrqEKwlXEuCYXMHy9yGCMyAZClwdTA
7D20DUn/ddxKhKmySoWIogMZbQMgsYFrsI6a9eTg39wLghpO2pAZl9g40VGmobHNULQBMC22v7OO
utW8mkxO/xMt1PL8DYdfWcmDXpoZTeSbdAY+5lNLgP4i/ym6qwGCp9udAJpzSQQdMr01dQHsG2iH
r/LUIB3YMWg+KlDfQgMpW/lUjVnZnw65R8bOOjooyyR5ydnu+zuJ1ZBIog3mv4Mjx84QEFMcYiQg
ySbXVjGy7niZrK7JdqfTXntXfXN8kKo68Fj31UT9UPFFbtHyeqR+HZos30y7A8CRQloLaGEruWuN
9Lj48pYRSuU5/NQnRBeQ2CaMX2ibG8Wve2dEJEYeK2thMVn/3/l7NoPPGj+DinCrujn8rtvXZisE
kkQ47JO+328tiBQP7SLgzWOzKcTkTW0AwHT27FJXoZKG7jJ0xOMP8OZakkZxRFk8HK742SGvJL5s
PYAIBFaNdML7BvkmRUdfX418YbNvt36vspqKu8wftDVgujLlunO5MITXf4affepgZqXzrXD9/Dii
ZAMUR5vft6KAzpU2kFBdDVVIpTVqDIWlBnma2rWSAiuatz1ymu3Oy72afeDTmvMDyo7+ujZeXtVB
ewa9nEhYIQ0omzdMQ8gEqnuNpLKyig/B2YE0G5QK3gG0kIUrGR9L0f70HbVYRpaSjZ8LKABtZrsv
eeBZCAL8Rdzf0ErTj1nYkc3aFS8c8t9Ty/EITFbB2XLLRP3tDowx7oQ2V1hJWA5ZhX2xRlxWmP+M
B2NjkTdRKFiv6yvz7l7rRm5G0b+eUuUqaKe9vQYkp9zReJZV7mpejyVk+1tbBFu/JnGYr77cpGG3
VzVnwiyxuMtUVlGO88oaztKP7bwil7eR+5C8p0Z3PkOgKDYojYpFu8G5n828QugCxKNwAR1hYgWs
1XCGjwOElrev/71TuDUA1FZ3pd8oRFfpFgslYnkDXcXRbFeloe8LUgpVF93uqfhliWvMV3kbxg4u
voq6+Yok+sgi0/KzgECOhkmX0CA3g456qLM9uM3p9Lbp15dzO08wcVmSL5YNihJ6IqnpJn6fMzjG
/9OGKszFm8UQDKMdJMR7Ol6m0hku/r3BvQkw/1j8Xwn7sp6ppZqbFBAPSbuA9NaJc5WrTxE1cDaD
9o5kMm2KKcAFX1wnh1WVk1riiagq7YaYv9a2ghru4tmh5UOlLLg5BtrC5kUKMjlS0pdpQXH24PnR
AqvW4WydUUCW6348P1ptyaZpQ7nI9/9Zk2shyHLuNoYmof45ySTstXxxACAA0V3aR+2BxQFtqO+K
2Wd42oLvjCOqbL/Fr9Q8MNU9AhaFrdXc7BuVGKAFi7CPjByZbb35m4Z59Ko9Rz0Mat+S2pGhXhyF
VOAcZReyiNZXLqQa95+VwW9JoEdYjp5c+LzpTlzGpTbIVaAM5/w5CetWUIKgBiBLrZLnbJ/KAta7
TLvUBKSP50k9+ikpcG9eF5T+B0nGjlIpESNAyv57OLSohgaSd6Qu/FZBip9Z9uWQjDIYjyDtc3kH
xrOQUjpfLvYEhRoAqCmWlBJXSF2oYdycZ4Uq+XFlxWpc2F+qO4jKRHZGNPogNgvF9GVL9NqDP2aK
F5sd9Vh98Xkei6cjeNg9AXzEzxgPhCBnnvcvEwm/nfTJf8u6phC9u2lp3A216y79L/6N65xOZ6pe
xXshqhAuMVUhqtbZSWf69xUO32GZL+r6AUM0ZTJeC6+BVF8b5a1THTzCPQDqk3M5Vqk46yQiK38x
MnKnuYoKHMSvUcVAOjoiiHx0ZfLb0Gxp2WvcMFam63q1w2YvJqCWqoeXFXDYgJicnKm29R+YK+YA
Kp7n6MmrYUrrY1C0+paik2HvI8aYXNsjjFNT8dR3D6diI0r/1zi0xhjWGsv09vptReuCnok6+lej
SK3lyk0D8TAEAK6MPSg45ACjlDhfI6UlWL1/1CTJDhwTNLKqVGfOJPDBwalxg7l90Png2PhSquyE
1C8XkkiEE20FDJvaLXY0WfwJfkQ275NIXMaPgtZDZY43OXTW4ipS0Iy549zui3VA/+siiAnOMRSZ
TC4TZf2UpXrHny1qwdTufZtHumM83uYqOCQuGSg7r7jmDAUlgZNpz03UbW7+gbbBYeCyJO63Jlef
vDT9Ur45Itn7vQmZJ9hdvQ9DZwwQz1cnQzkQBDiF1MUIzVGlIwx+VGpsvJOUgmsLwTQ7FXJPifMs
xKOLHqy8xbnZGjMxHw7vpXJv0GKOD8oK1GIudm2PAmkLeMrIbnAXA3sfuPBhIiYY/z9iZM+5ZdjI
JYOpG5X4myxgRf+hR61AX3RI8dos6iZJytkaxhUQ+JgWegEZEnaBZ9J7v7seOh+3AADpN/tkk2xR
72j3YcogJRUS85KkMB4JcM3R3c4L10Mk8xCPXyA62Jb1RqjKdxJoamrP0Qa283f9PZjnd3Rl/OWF
XO1FAd/NH+jIKMXl/BMuSKZwdYdlUEsOcq5JgVzwGYwNx0ah6D1LvrzVTfm8d+/3muG2eEU7newm
Gco8g3FkCuH8/9fweCVbBZIhuAK0UGV5Zd/mBz1lmoNU/Fl8YqHtdTGxc4uG94peJtqorqy60Om/
J+ej4fS4Ht0dkavQvHpTcpGvQ7yWhqAAfv1AD1TDaW5olPwrPbEt5LHX2i9P840JrsuoiOOvHkDW
RsARKvf5TmPm9D01qBUI+mcSy5WEaIKY8mjLkqOtHB/SBocG3XYVhV/dwnMdggeLa6wvk5gUEvDU
4v+1VlCpfRHFWmQhOGQgmbZJ7Y3P0bk2Uma1vASGGcT1JcBQwirYPCuchyWxKaqDdEvmMLsivZuK
KdaQU1t/0q/QDgx19fEhYnoUe4piOQwZvvP3xJx7pn+wSWG0e1ZV8qzGzZkR5V19LnGylIeUo5Yo
zlziVLAWAKhEwHphTtfzgHPGpcbOD4NTTAhxI13lG9Pd/jSiyAsay8g8JF/Bw9CaRJMJ4FO/5pTJ
NDEYMULUghGnQtf0uf4IQ+t5Tred5Kyo4hQoC4uJO3NMtpNWJbDyHhe132Cv0CZfgc+QLLQOCUNN
X0Aai6WSSNO5Wy6Rwm9ha/p8VyO1gijaikplnNFOE57TCztd96/5aYsoBkdrVOVrRHHNQxYL0kjJ
i6QPMv+X9E9Ztf8YA4JQf3yuHwmBtHRu79PWPTf7VS6jskJ5uryeduTvbYqasi3e+t8vVb95taO6
oRCVXg93aqMnHUoM59wUIN5IZHMnQi3k0SbEgbwT6/fLPAY2NPDW/jAYzEYQNVqTyR+jdH1rrvRG
qfWrDB+UHiFfTbaokLWYYPTnzZA2+GwjmYoPcb7QWlyFcgY0POKlXh8MjpURAk57QjTHuz8ivv8V
x6pyV+v3hk78X0IA/Iwdd3EJx0a/gluxTAS5CmH8nKsF3tJjDWkHBSDf2zyE2uKALQuoV/ewIeI4
1IImtShc5rdBWN1hxKafsv4F2DHa9xzJ+0q99zGzNuX9hi+l0rJG1mcxZzZr/F1yLfXyFwCdbQEX
hBWPym8T0ksLTDaCJbu00MfZ5GrohI5oy8TAKzSsPZbTJZoBwGC6Wo6VPM683IS5LhA0U+Oh5jbM
STpvKdRdCLieOmporzqXzfKTqHujFUaZov1u3hulIfjQVx5C7GZkogIdPOJ87qqrGXwiFGjpZWeO
RjC8IlXbUiYvWf6t1x+kv8V2XaSo7n8iSFSesXE2tkv92dwNI0aI1p0UpxLkZYAAFf0xIPkK4PzD
gZ3N8bNNxMgBoHfbbvRHmU6lgX5fAg8P5Ls7m7H6f5w7J6pMH+AH89ehj8h8k8wbV9HBD4WNxONw
LrU3R/67bMH/aBhcQDZiMf+wYwByyaJa4dJ9V40EAszbPR+wrkZ1dL4b/WgbWD+Pwv3md7FtDIHV
fY7MBswQ1raR/bgkWwAN05Ovt40T51i6bkY77MIFDtBmYzZ6MmUoAqKdwZ0MxXHapI1kSjtoLVC0
B348yEJEogk1ahYQtpOfwMOpgLLlTMFqG/vPeDfnN/nFA2aNT6RQkOaNdYLJBwDRdKpRLABgk4QG
9+zYq1b1ea3XU/EDnzwXacPvWMlFAVLfon7Uk4pvGNMnermYeAH4E0yM8b7RSzRyKr1PlbqeSvJv
65Uv9yKtNNsH8PfeS3BjOWAedRhMNrd2PVzC6YL4OOj9OD0zxRuwA39mivj1a5DJK+M8TkoBKzoR
lru+gf9vmMCIjS5FMKma1sZgArMB5JosRwyufG11UfYFvihPoaK85LFF1JtebDeYidM6fK5AgZa7
8okGK/dh4oN4lBTsnpTfPlq7i7CQryOLoSZX26DRnnIhqPcYKPKF4NQ1iH6wmby79aHirFNm0rDn
qCPiF/dWQukLs/mTVeu2AU14mLn2sebVG4BBVKPaYRV3m3mRB276QuUz6JTvHInRSoPdcDsFlcb2
mdnKk5YkcWUai6ulwZYmeL+WVWKVkwpdTB4KREnneJrOk6CaE+V+2NIVv6J8Robud0g8RedmZGJr
mIHST+N5xtUgYwodHxGrB4x02jFMYytc2QTZIvKqFE2MpKnrL3084L6DeRO3UDw8KO8IcWeZguxP
/MNErCNB5HyyDd59JQh5OTlu0lmiANpKgsyANCGOAdTDr8+xIDIGNNOF7MqLXUBEVITZs+izVNOc
MM0u4rLupX6NfU/hRzNX1jSMRXBSRGSmi2wFW3yo8bap1Hi2gCrh9RAccyWMm1XxICIuYO7HGn5j
Sgm+zTwWiXSvzc7VDkta1U5TFZdjJPlxe21uPY5wFAzW4b9TC5KymhsJAf6yhNAfM6Q0mR88eZJr
UuJ32gmdT7vFtl2UL7SC2RmfRHQkGq60vgtnhIYgMppdtkeAiEAh6+jTojl3HZHaEdj1DmPb+Ixi
V/AG1cLYSSZFOBILYnoNvKHhBRxxnK26QSBh1Z1KqIhg+ZbmOuBEO4BpDz10f3gYdlL8SKdsQ55v
XQMwPy3HhjuBQ5AuoSDvY21yNqNOc9lG/asat7ueZyPC6w8pmeSF+XXm0Lfty3309uUV6DH7AC5A
jhlbmOfnGvGDjRy/hUUe145GMDj/0EAG3Ke8IGmO6TOEwjgwK/DROirHjmxj56Ymkb2+EskQCEtd
aMlpJCgxojGizI0KCrSb1KZSoInREaUoiT02bCoSi7tS/9htass4cpZsNieanrRq8R+NTGGL72PC
e1myufFDt/gdGsMayWuBiL66UtHU0iNuHYabZ3LyDGZm9wrLAFhVAzi4NubbTyZioodMLQg0vLYM
TTYPUNq21zFEEk7gYcLNQQkTo8ZgcxUJIexgpfZ0wptS7x9cn1eaDoGMXglli9hcruIPkRcu9BBb
tOkYrNowg6s1h3oAoEe2HHd5E7priSTWVt+rObQLINiw4yJNJMXjFPOQXxsmk3Fct61hlgunQRtR
IN19CdGUVH6XBqVJJlW6G3fStoED7kptKOWMXLaJf8gOLMHYW6YZWEWIDfii4Rn/uzdHzA6NOkWx
bVw96427t5DZYLmGHwIGdzNzaEcJcXafCnPE0dm8HNUzlHfEgeaRx2n2POHme6bgOLIb1JA/vUcy
QQnHMosNn3mTPuM0XVyzgoCK2DNWxwygKZQcbeqg/0iWd9IV5KMVpIfQhT2nv9ddq17zTRMlgL/O
IVxz+Qz6yaybb94vwQRHiMIjCmi+ZlhrREbstIigLXd/2qNMmWYCtVlMKKECP+rsiAuYVPckce3e
/pl90wtgpyfAvQklbbn7AuxuLrQ67/oCHB1f3Es1WRCFfyYp/Z0Kg+CVoi9hpVQiwZWqBmhMJl5T
O/MJrxImyVf1WQe+C82U3qrNs0wUngvZ1Wpp5O4/x0n+VTqWsJmXmMnC4f7A636Mru92EQzqebJD
OViofjRacVO3/FMIrSQMe+3q5OVLrPaAJmkI+F++I+aldYHMCgw2YrFQeCQTDgnHntCDzWujRrxb
Y0fULwSOZfz9T7wYQkRGsAJB2e+ySX9eATOENnmOCJYacUVjT9Mg0qBElGMh0oroBvCXl6Iah470
almjeBB8W2UxRkWs5wBmRGufASzedq9FLf50VpmaUx0EGs0iPhQFneRmlHSd/6YMYpuqB55wVKQa
2s9WnerNpAXXcbLIieWWn8/WTAmvXZSXYxaWXm7uPh645O8ybii3vA67Gm+dZySPK75hvLPuZJWI
k04kXhp5EzLmAhzv6mqqCkmCFofBgNw6XX68pGO7g4IyGZiNmw8NUsVTwuYnSvJrRPXr35ru5tjc
rabj796SaaBBwXxHuQCRHZke62Rd/lwvEkXzUDiNqjVnWVnP8FCIJG4z+h0aPcfcFKbX1WrQyg0W
3to9PYMnHeZViop1PNtioSUe7J/Kbl8ZnkYYjuWJY7EzR1VGw/8YZIqzHyYiFYzaMZe0lVtcgP/U
L2UAGwZQarb6+PnyRNihVn0F2fTCg9gWTFVO0eveCjzwwndutvnS1MRtD31y/Op/FtS9hqsQfVJl
oVhj4npO1Dv2ExCfM1T6YaOxv7ZqjsCQKOu967VUtyJT7bdL0wnUI5edCKZ19ruI3eAXtXvJS5Gk
dY69MybIHmtCHneXcfU4bjOH8dttkLNp68A7PHf8gHwbehKGNPjfXd18JqSmv9r+5aaW/Sd0AadP
QtR20lWQ7+mXj0UR+1WL7uPt0GU9ZlwiL7D1tPVtYn17cPK8euPx966VwiGRKd1K6wiMZjX+EqwR
0nSABOz0ZQq4kCZOUdnmHolRT+Rc8t80u/fqPtZq7K+7uqw07/FkipJAsFBHqCvDiDEcpT5xtd3h
3nSgXQnNPEt08T/kDkhNRPbUq46ugwH3XKNwEcoLWw+AmCCKFC2BJZ8YwRvMqsSwBwch/Gf7gy1j
akfyGCJ29D76owKNUFZz512qg11BmIj2vnb1IBAv4iaFNYTl/t6PYhTWhR8wBSfWzL2KsCDSJ2FO
yj0ltdLqkmcwsTskMoq8XjG68XBjMS3O0RMbXk71GJKpflFMQe1mxeT6vEuK5Zttd9jRT3cfkFQq
Q8GcRrXaluy1dlOxg5bxCCoz+DGNcAYompmz5DzuIE/mfs0pxJds2GwOkN7R581UF2/wMUrJHGcT
7H0YAIHbaAWmAmZ7RUruSKN9MG0dAgc/VIjwRFkkrGrK8BacxRXMYo7O4obHd/OPd8JeXcE0ajbZ
Zrnzl8jGSuwMESEFCjJ75P3LVJ92DbUBqxV/fXjKL3ew0I/HxdNDQ1mneRUKyTIYAzZcBd5wkh2W
uk4w9e2K4FrDL24gVxp5KQTos7MJataeEcK68sPXGynwZ4XFm0XzQnxBqvXbKU59SgGZeW5fESyc
rynGGiHdrGsgFo1zG1b/B1E3j+p34Ny09QJztvhUU2vZM3m8P+EuNEbxSYOd47k8MU4oKHLdgNCT
b/Cb3/z+GN9OKVgbNU56LGquaMy7L8ONqSk5PxzibizQK8PVEenUW3p1cQgImKGP7PnEWY2LvQyC
Waf2jZ+l3Cs19LxXrm49qedHuXvBX9VftxN5FBOQ9YHFVgpkDPYp7FKT+qPh7ns3L0stmuC6k97A
8d4ikW8mXScWVGL9lzsnHd+RXjSzS0AM8GgdHsZPo2t/SlZ1EuyUj/FPGTThEDDEV85Gq+u5DMIt
NsYmW2jVczBhc2qnPa2yoZUSFIHA/mqicz3cLTshuj1zeKRIkBot9vTkPqIsnCrp9rNplmLbW/cp
lT2ZdYazv8fydaDSaLyoKQXZM/LJ6TwzwZiY7rVRi+S/nwca3m0aUfpsNCpyqA7uqNn7PJ2UJOaE
aXu7uTuhVhk0HytCC7xq1n3iDHFUjvd0jrIkyvt5sOYF5g+KYMH5FllfSfYBVMijxmcq/BasLKoC
70Cznb2x7iSmknvHI6Hni5YY0LdDOpmURmBkw4sWa1kMvki8yy2AuhDoBAYM5mlJMkEHwnmb8OcM
NJ3AW4DCzB4Yhlbv5zMNBiZSudvGsY24q574++dcb0ZdDXAKj6hG67umWJCca7aHAbUpJ3Vd0sUf
+YzUh8Nkv9F/q0MWrnbjOkKOYbNZu5VKB4WjJYscgCTnzyz9i1XPVXGNUwrKPtdN4uTfJ/zS0ntt
bVcsCei7ql42nhdJBVv9DSiovf3/b00Afsh8Ok3j2S0pYbo3FCLWeu1OgO/+BWKxppxa3dIZ+IgY
IywP8zcVfxLu23KAmLkxcKPsZ7iNzPqBmu9Kp8kta9fhkBMS0WZIsLFcuErtz6Imb1lQaLPlT3JY
Ue/IPXDVENCUqMyDdTg4T2YttoNn+HRvBm29gR8JBwOj6ce5/jIcVPy4kVZWo5FUZx6rCG6B0/8u
Fj8mjnd5/ji1wPTPl3WuEGdlr2KfPqwoWStBGb51gbyRKaZQAmdOmpzyr1U7SELkJOPsR4OoteET
HkyEoAI3oJ1yJcm8onV1M0yxHPdvBgIBehEmGStpmHaKEWIwvYBigt61PE7LOglgQEYqK09ZdV7l
5FXjuYELMTklPdiSXg23IOFtUFPRoTUQsRIenjquekLzcymJhSnncHOoPdKYvHWiezG71vHoK7L7
Orz2atTe4YCmryD29GP+9WCpk9k+C5pRYm3COVzo8N7Mels/aMxGbqOXyhs8FxZh4NNm6+L8sjCb
J7TSvC6x9Cp9+HX+9WPH7BShrB3is4wU4ZWDGEz3tR110uSUOg7s+bgRHFGV26Zhixb6y5Yj43OZ
/FBAxffWlzkVe59stfkpjd6jAQPqzPUygltQY9Ap8vPPcMAHOwRa+osOmQuvap1L6K+1X24IEef2
nF7wcBDdRwlGa6DBsgZ6brU3YOJgXTqWebltGJBvni1SH7wOd6nhPMu8SPGND7BDA8p9CyS9N9K5
o+yFHOJWZz7ceQ+HJNmua16VNOi2nHaWUGeKn55YA3/xsn0iv8+mjYg6nlEAgTtrLRRY/eezHFl7
G3Y1e3+5Ecy9pdsYQ/kpTIyMychPrJvA7zgODw+pvAIGnLPpQdB6nv28ZZzdCI0bIrSygrj/WogC
o+M81z8tCUkFMM/+2/5huzLaa8jldWq2ai/G2Xzx0JnQ7DkNX+plxv62qQsL67noWbQmAgDOzN/N
UKdgnyr2taHutqWVmNXpuuPX/+GecQYltRco15AwsIshC/Drfa4ep122F8PvwYENfoc4ViGFqdvR
TD0diOn82/fcBv9j9unHPHKzq5y84jSX84D7L3jLnRUYsDNeDTFvFvYm0zQ6hXOjad7w02YW0cnX
RwUWjatHgiVsmCn4ohasRWIokGsuet4fDFS0Gdju8VWu/ZBWbzmxoqZym9m+wOikkvU99Bp6HPjN
eZPdszCzPoW1gQeBlSBu1UIiyjfRmhGHSJER/LwmJKTTjwBid36IHJLDyK7JvVXUHm8zPw9Ur2jH
z1ZajiumJnrq+Vibq4bTx1tJ4eSJLZ09zMMbXa9mCHpEWjD3MWxek5M17D70XLTqWlm5Lh0Cylep
g72mX7gs6y54sJtu5cIeqsp0uDGSlOAK7cuPvBYIJ13YD4LQNxGNdSKAcMp+ysFHUIsL7j4Qd5zB
Dn9giOhfE4+nqQVt+XnIeBO7sEp0OKiw94iGhsmdaoYchVVp/jqF08AXZbzraKEhBxMr6zDxdGuC
NTOHRfRdG9drjZZk4kDe6MEIU1/cAwFH+Dr6a4nuDHm/HXTdsp1Xqb5T+czT6Cd/4uBoHx0mExXk
rxM0BhnFjO6Puwt1MVMEqaqDs1I56kfSJoiF7z3Dbm9BMxzNg76BrCSWR15Uc4O7TU9ujg83zECe
RSBwGdY1ExuGX0QHQ5elIFSJE6ypBelgVGRpA9FkO3PZhRSFUJ8xyMte9ceAxJde+u6FyFLKf5Ye
sg1ecwmHfd1kElT2CiZQob6g9/IqudjygzqCZ3Q7q18qZ9kk2GT33nRmCT4sVhxOkKclz7NoKEMT
pB088Y4N6Ru0gtfFpjPKLYNnRvRLYmI8OCUKHW36zqUAXLxJn/rW8m2LSgyoKHNGppkDuV6gl3VA
OF+HYsQ8mPi0KVA1F2gESkpKKqSuk9gpNJTQK4Bndu4h54bbOQza/yHhhxEObf8ErUfKj/dAplAj
qjdfrRPZ1lBAm1XeHYg3zti+3dRoml4OYBE0RNCKurTO8DtyWxnGZRSdOoDERWFncC79IfS6JeeL
/4EvJugB+wFfTNCSqcJIYaiN31EY5eyDG9YUelE5cdcKe8gxNPE8PXVnJfZSA20Tw1U7rIrrvdOt
nGEUI3qJodylJD4+s0DdLXDnLH/tYpi9kLmlBZus1qYjYEqdPjUtbKcebGnmuVZZVJzfJz67nbxw
z3+B+/Au8kHCWL+axOMORi25xzlOMSlxHJLLuDQGqy7lpWn4GbKSMfvddLuRnJcdMc25PHBChECQ
DBJGHsh4r1gStgsJAz3GBQg2kj+TMeRkEoGDJuat2PVE0Naa2OIIgmux++O2CWLR6wJmZ8/lEjP+
7P4JgXt8+9HsEsrUzNh4PWPrKW+/H+NsqIy5Who7VIPS2vK5ktrHPdEIgXycXDVKLk7pMb2FQXcN
6giWSHXtWxE33/eQrAB4/DvOGBPn3iMR8kxcDkvAzs6hcWa3+9KD6/bWeTLkEK9fUk1nqoTEyjS6
X49mAtqdnVMR4opITZ8srmDpWVnBYleiFuoYEwtDUKAshw6y6ZHrSlv7KF7u7SxsR3l07OGXOLEa
OG8XD8WkKXYwtAq4qr7YrY7sPUvOtjh5mO0Wr5DUB2/aX1K7MO73IkgRVAZcRFi1H8JBA9hxMKCT
FTwHsxFHTDG9PTmStSAo1JkzBtpLsbqEPHJqKstlAQDZCGVpWc1lydQ/ohbe4oTkHGFlt62NI/X3
t1fSWXiWS41sIJ9IIhlXLVpVrNNwxXRG5igLhO4+GmjlzUDottvdzXmXW57sjRkRXISgsIgStOvr
U3T9kXcS2ZWoZK4j8s9ozCoiZiM5RnAPGdh3fHZNCvcbUP95vy4ZfyRAY42wHmv+qIXb9yAHJqiL
Sa9Hw4c6YHsL3At3S9i6Klis5EuMg71SghxAQVxKQvQTZrA6Pr0Fmh1FtxTS54Ev4qiX7IcV41Yq
leaB5FNru8K/WMCqs+G0NYy5M5hjtoX0c7z+Lt0K2PRoLxHlBMJKheSm5iBuMW21qwUdTJQjb9cP
u2ie+FAGywcniZcOVpuCfUZX+7Owv8gXBO5rHBNMWM6Pem08r8V3FIdFGozkdle2lV8UZINZ9XyC
KqjK1sVgb5pnDD9CyKm+1VFclZev82UrmTF4PP4RL1cLYOPii8VM+tzNrO/L11ZkUoEE+9SCDeja
wOc3kxPveFgqIE0WdUggDsbtnhq2EGRN+RwGxpJUDTsAwCtdhm3BzQSRw2b5jaZDHlIFGy4HiVXw
8RQRsVna77v4qVoY5xwa/gYaN46mstzdtFHvr7fiEOL0z27WPYiGTxcbWxWUbGtcGKLevUjGsGTE
ikrRLeABTm0RPcZTfiToy2CPPFuBhbnmr8beBb8lTJN3uy9MNcWQlz7CnL1RsEo14C+pGttEcVA4
PYiCwGssHvS262qwL1RZDdmIgpSy1KmC89EkjC3ncU7bRqhE0rmlDhAp2/R6HLaEq9+Snj4k/Iwr
0JQdbKIVvwmZPJsrz9e4QL8p4buvrrp8he7d8R2g1yPtoUfeAjt6R86B3fVV85gkt2XdVkeY0pWF
tV77LbbyIVvWh6G9A1R2D3zIIsRoRLVprRct7UXY0DB2ofIcb0pGQgsfk9uACggnnN5og/gDnZUW
Aj3utbTopNLspITUtDfL3jacm1W5YFsg61mckNHN4QOI17r3Z858dA/BOxT8I1atRRwuno5U+eDM
FNjCrMUAe0an54kEB5XBrXzXEKe8kUvbZ/FVI3lKVng+/et+n9lobXJC/1Vvg0h/sKtyJejWQfMR
Ii3Psrn6WXtFPNI5CIpAapAD3LBG313yXl3mUd5cyalvclBeu3RvRDGuAFnb0KveJOfKpu6s7Q1K
naBFoFezmfpw1x4eF5tct2ls36Os3GH1B9P6fiFA417EWwKL/lt0OosS2HyOotLGJi5pjnNU/1sB
HHcMdbV2H6saht0BxJAqo3teNj38UMCNHNrg0uS5JisKEZoUqa58iZUNll5/bWb5YR7PmIMguCRP
0VqZb2RuYVhYmrz+0bup5ukMJ0WsLfdo8nAXChOE2jBczlCMIhKSMywfwX7cqRTiEom75WIhmPXN
eGRs9tCkm/pIxwwUWhnT1Rdq8JglFi/Na0xpjAS4Ag/PcpJyCjChr+SwhisX8fpJ6xgfx3AnKbk2
2Es457VNiHD5ofDGToEiQXjc+Ego1b08KE1sHeoap0wZ0jv7bIC08/Fqkt4MY0oaTnuZprHUxRkt
qaV/zp0YmT7HxxBetCpkolwxJAb2/bo/XS9ot1w4IINUM01k8fZriKxlcGFBLEylR98JSwsxC/JM
A0bf6a+dr0Sjv7wfKp9+U6rd9lzn1NnSIfSgu4yHIzskuXpmPBBHBuvsXRa8xaMH2hBAiwTrtnac
fnRBk7x8Or3BuW2HuQzrJgbAKkadVVlzpuXaXPDAQMNi07U2OBnQlp6SxlluR+qE0C3HZgTNYNx/
VupgplKvx5xwJGcTFPKRcGF6mnHw6r+8C1aR85r7Apx+H5lsMHGDm6W82LTjfcjHw/GsJ+AhTLlL
aDXRiMqaPzGW5egjJwXKkRDw32Z84DMi3WKHgtBI7B+cXdxBCg+XbLtz7oYbKYvQRSnyJDO4TxPG
D/DcL1tEXQtCJGM7tSP5fqZdnW5MLCMEwYdFKy/DNLt34exnIPDluciQoBHJJqBQhRggP6sxh0OR
b6xy5ECZHQYLyG5t117bU+WBQY5FWnkLjmQ1dWjVcNDbRzIHMA+EGSj8g0tZWExarbVHSlwTovfz
+bAgVZFGYdWX83YSNdH1+79YPmPl2G0NUGobTUyOef6c8IwcUZi5NsZqgDJCnd74kksFB/Mfw7BD
ZRzmqzl5JhIr6vJ2SeejxiCMOlNkugDrqtFZsP6ooLDG7i7kn2G4Zprqnlw/+o75pO7RJxiN2nej
09tlle/1U/2gdWCt2Jm/QRn9HmBtyMNZ0Ri3PgkPsNWMPrypA0G6MR1IlaKg0Iz9Iuzus7vFK/LG
+8TMHsnvWkDcW7sq780p4XoHhq/2mwrt7aIJIHJgdDlQGLviYw4sqyoyHTYoEU53v9Nzc1VCs3M7
3FbOJUpYmSY36CIBdpQ3m5zuBwhFfRkVSFZLZkF49XDFWhVwhoW3jJCQVEfZdrWxpmoAQCNv0Beo
M590ellcD2vc+IOJD20TbE7a71zmgFRIxc6wVW0Vfv0d1MrMLB5AmQ/ozEV6aYWAgQiDhf9SCH8C
j7seHPhqXqCrknu4gY8bIMKPHcoNaH703O+5AphRRAEBG/Uq1ZD4Tb8yYxGXaz4uQcnpE1A0z8rs
+qNqVyOjfQMZdE4L+IFY7YF1l59YqeJCLgzfF1dx5vr6iDTrwrf6lKzWqd5vvQFab6i6Y5KN48N5
vbO55qfLvVUDMZhktlkUOaHeB0hmwC2m2Qu/Zpv86Ao1ZNmf8cpAf0l5l7T0UV8q/u7bnB7/jhFu
XiXGjka/zs9Eg0RQk4opPfHp6PKEa5SRWSxaturO66vedVuSFm75WjhATuHor2/TNnp2Z1ZBoBrP
lL23X016b+bFXfzKfox0PHNtdA0UET6/v+bX+o/uCPW1WGa2H4X7BA+BSfKRZVa0B7QT6PmJDhgX
tBATBM1lhRlKmTXryMC1y63OdKR9CEYgBVRdHa8KDWBnSJUMe2QAH1JmhRcDMEso/uIRTvLmZ81Q
/FDhHtQLAdC7hge7dUR4GGNjz//jmrxvU5BrT0qQHoLmrB5qQRgeRBmHFAB5Eh156rh74shnmZnr
vQE1GblI1u+Yvrcd7sssQJhZbkYaO04kBMWhcPBlwrtkfl80V1C3dln6B0EfJpyvRQPq25e7A8Z7
I2GFlSbbt/0EyiTncVgnUCRkQgDlEsYC7PGQsreEYxyMGkooijArcdWpSdJQbtzpPSRQZQTHHCcz
z5KnaE9k9oLpM+j8oeify4eZ5ofCK337rPMXlYgjWPL9RVkcW/ctwFlnFvTwANWugsH/xy6ZUcNS
MR97p5dO46bhHwULRgSQ68zV4c83cs2imnchZ5OSp7azOXWES+pDjbU4VcFTyuGFboXRr0Mgh8uw
orPEVxxmwsQPt7Kanh/9rwkUC/e4wf3kdwyELsUHaDwCg2OExeZ8sU0V+82i4CNF5okjuL4dll6J
0DJHDtzunCWcw6ZQFEY9wgQNaEhkgpkjKux0O8mIND70KoWWu+OiY5SzNc4GwGYPlBNJigimgVZm
0XvpFYeTaz+fHORDi69VD6nEBaEmxzMYgr4tATowGGuvst9sTb5XSGbjPQ36Um/65FaztIMzDEHb
q6NgZXgMI/laz7rvmNrbwnW7chp1aSaAb/UF1QXsJ95jT0xJfB9lnJF/QxC/3OXx9gZqvLNJdDLs
yYuAPgNm1wHyWRdQ7I8KXg9dQPywlZwCzMhyXxUsopX8B9eg9eBlNHYiuXFDytMPJ36RtLv3eK3C
QA++YhScvGwIdZYKLCX6sESHRQnH+sjGSNQPYcZEpiinsW/sQ1MnK+0PGxnLdVVk/IP0RkA09Gl0
EOq9FZzHx7uWiQKftPr5yIRv59r7fbdxH2ZC25I9MC3X0lyBiIkVml7iR7vi5WbhPfxRIB89UfUi
DugpRUnQdccv7dmBxK3NkGTYPPGkLVJw+To4fSwWi6YFb1ZCLc3qnXe70SMT6TOEdbF/BMxshi/2
+oWh8ovd4ZryPO1alI6Gr7Ex82tpSvYNLpsy8N6FadATZwoVkfQEMw8YyzK2sbPucP+1pdcSvA7r
WmlaxokBJEfL4YeyEW2lzcraJAZ0fye9H054wEPfKD1IVLqYbO+f6KWhPP+Nl4/unCpwtOe8zs0n
NBU70JNMF1J4ZNZEX5QSFaMNj/vR/djI89JZG3JmYNKCnLzyaQzTnQ5P9gvh9CEjbqykGyTk/DO1
+gZcGoq8EXmX60FHrCjvBmtfsLTgfPIrkyF9gXYW8YgW3a/pNs1nn9ara1iAuAFMQmbPCRVp4hiy
LpsODJJhYRTA3LGq1C18wBffL9Wo9dTt2s6rWPoBlyC3l9/79g6dPWz7fUiCi6POhPMybn+Vk49I
sOMp5LDQJ1wBQfDDlhumgn3BeWhKOuKTVBX27HFg9Y+pk6Gscktl0YOGU5VZqc6bkpKadCuOB5cw
H22PiYVVG82+fx3+cMUX1yjTPhYeDHPkzwlS/9PmOa8ZGnkOw3TpqSy5RTshfTwI+HERtPYS+1xs
dVNvCi4u9+0gft7aTsIgDOxjdgYpp+YbiSR2ENaf9JfOF9vfPN0x8zJj4Zg8oT+c6fT+6tk1IkWj
/skzoi8KgbxiKkufsUmQg9f7yDFkanDUOKTz/s3sgK6Z6ez96SmmJ1rGg73s7zYf6Luf3niRaqvk
o2GA2besfJjTjUFqsMQEs1oHkEnY+XdebA4eaqS/7mMNVaOQygt2C8Y5zYiPGDjtTXSgtSsS8BiC
RicAK1sQTCJCvBd2B0PydyYxS3RvGW96GEmhtfaINkf7l+0k/hGI3lM2j0o3IjDAMvO4Sr8DY0V1
LEJEwLY4OcspKI43TohwnC7qIjvtONZc1Xul3jMPznVQhTcirb2RPjCS2kHm9lFRhDlSarIrDowd
B8xIp8aumcvUaoSNhlIYBRmK0gDr2Hpk3zCgyAMKtjoo23rpml/4SthFtISxKB9aymPfjZhNTrNo
Tilp91GNfVRCclvMM8N9wdbdI+9dnitYrKh+zWxohBe5OhLLaGUAVh6I2zOPRZvQ8XCBFch/o43/
MiFkTgOqumfjAlSfg8wYUR5hvKS5pP7EfVNQ2JnfhsRHksQGsAH4uVulmcd0H5XZSf7LcCSBu+ys
aa5QnNZmwHo1dzNgDRSrs3Rrdt4a/eFmzG625N3vwr7DWpmY2cLNsb+FQBlfrajfBtxTOlB0nSC8
rL5UhRiEPg/Qdhw0hsT9cDFfJ+8kXkpMbe0cl4LYxYjW0TGn6Vd2q3MhuWbBYpMXhcW2q1SZINgp
uNSm6tvSheZBBUpuwgLFTkRFo1tPHmhBta5uAIfiVY7U2WJCEERXRxVv86Al7FcrQe9L34nPBW01
mmyPoIaXnKHnNxpdy0wnZj1tHylj/fee/Xws4WA2QwQi2tgifLWVZrTeHrQjIVByHikpkHW/zRXM
QKNw7juQFA8UN/v4c+a4rtIfbrAju+LZpFZn6WFx5n7HYZrFkpsqRDLQMUNo7iY+7JXd6ptzaeBm
6D9FxC2wFwNJcA8J+xWW3hvreK4JPOGhSufFm9JPEXOPoUjANTqNCk+K28Emr86zur+Rp/EJm3YA
n5/ar56mwQQU65AaC4eDtzmfmK9GU4zV/cL0FK0FdZd0x/69Y2+jiZ6EixXbjTNS6FL+I8r/AfZI
nUGxwdT+IhCN7OsqbUHMJbzjxv/mH2iZ8oq2HJWVZ4R4TAmfjwQOmcbFQDWp7OrRVtW8TBLHME+t
JdeQ7EYLyyN3/mS2VpKs70h/MREGRfuiiQlRrjH3K8GC2/0TxABghufFR0XqNgNoXNJua3RONWuE
Mmr8wlGfokOvppyNk/q3nUtpZ3gWcFk+2URjChWLH08ea+profySlX8x/Cd2oTfpNs3NzWqxdZvp
j3Rz/clmTgI/gtagm5igiPygDEeKPVptSV9ad/H7WG3MCj4CjjGenV5taNti5tZVC7KZtsAYcmnE
QY3Z5QnGTh9PAZf57jurkn9ejydX9df5+vHF87BeTwik1SAWcNqM+WZmXxMOAna0fDd0nlY5EBSr
HdoUzcZLTIHIdQi3E34oFhAA0+sJFvtNLmYH/hCergbiSQMzSs7x0H5tf+rzHg1e14JXZTiLhI/Y
oBrGHtTySUMvJZe1o+LWrLMTtUq7DAONB5R7SpiP0fJD876nlCX3iYmXTYIGzWqGd/2fkH58X9eN
RjTIP0yE7LOd9kjM4RHsf29sfG3pU/ANnmajeJAWAxkxFtladpMErEzbYyrOmpiZvOVWvUzMqbCO
qsaOjcfsMBIRtJJiEUgTKqPMtai3HZC9O9buEbqY2P57qx+nqowPH+4ErjICW7ZLs2Dns3NmSDmu
JwNB+FOalVcvyU/uEfVlPnSHU9OiDMV3UBexEWQuvsdqvTy8MyNZBp5kNTZYVMET0AKnJ44GF3PY
qEmS9o134/4ce01+rNtjzHsp2aC9TNPFrjUSm2veucm9ot42QOBG1XDew9DiVurdYMw+2utOiPsV
lAlpOTojbQ5XiQanlWNxX4IdNYSLpdU071lpDaSBvkW0ZUY7J7AdCS7Twx4J2AHgDnGhyAXgZJYC
YUyV61vBvO8PMQdaTQ2Pw2aUklHXu/O7gYyx4QTaXalirCraoCL1d/6HW7iciCCSAs00zyFd4ydw
qgZ2DnB5aHp4W9glVkABFTQDBofp9zFJNJUvRBMkh+tRwA381YXPJD5GnuNsnbf2AfpAuKNFEtOO
7AmLW0H2dSP60agNBLjFw9Qm24CrT31uxi6NaNvD5kFME/iaGX5nP/cVZtczaxv1jQu4iu5LuqYW
9x5eEsoUbPd4myX2KdQ4GodNijjfql0WBGdbO1wC6LHIbae9+ohqzk4b6Eg1maVkZJ40qEKJjSwM
BRGXdgUIVSadt9+PsA3AOWuxpGZW0uUE/7H0bVpi0PniVjhJHjW6OHM7pzKQB5y1RTvYQRR5T8jY
6XQBnojyQn8ud53shOLuVSTR3nFIjExp/5uXq1b1yZDIDN/Uu6kXnK0056AcoX36oH8Vn81oMb/P
91rhPlJZdax4Ov1DwCRVFpnhV9F8Zs8gJ5LhuetZEeIpTW/0w4ologYThfy7UzBFu0qL3HGutRfj
7hPPV0jQSdQIBVG7Ybijw5bUAJFMsuaqg+EPUIbAZQiS7WcXi8GdvfJ3g9Ur7VC/OVUOzIOGpZhj
Q6p97cWAJ6AM/a6D1C/iGqRz7AX8cVjYMz6Frarx4Ht9uktkum7fRnmTKBhSQOmrptuSlzQ+YVfl
27blwpQlDz4qy4phUXjEhjzbUoKOOxImBA2FzLU6nY7CkCLquHF6McYVgUxVxvDu9rX6giTALx48
UVaeXi9Mwzg3efVDZ3y65CciG5cfLjd/sbWSEs78MnRlPyPPRHKlcZ2390dnMj102+eUcb6GrRQ4
Py5oBGM+QZwOxLEKr/GR+PFUCO5Z+Iv5qNqLIN5oPsRDxD62fb8nrkCPTYLYcpgpHqC6H83odLg5
yJe+S7FIXaFnNh1EVqljYTD5wC4zLFwYooKO14wadVG6zpNSxiMTg9fCIQr1qpot4jSQnUbnd+n2
hAEP8WOBQr3ifKPhaEk0utHigjebrozuTtYwBIbvv9XTp2CGKygoZpASFZbL6wppkH6LTcqlOzPY
Rgrt3CUWYJ2UIDcIWgoUR911uB9WDHkJ/DIU7IlQzU66Z4kazTCIsHwZ9p05Em1t87CgLWJJLMZX
+AzyOBTi0qXiTWKz4oZG1+DDHh8TDxb/gbUQTtzXaGPPZAUMFQPoABkxP2uhT6e53swJxuR9eWKy
08lNKW6N8oQYIj5vKfnLeWUnHf9x6XIFAA62MfSMsopWEUwcwmD14ubchVrZurHj6CU/S3a5OiUv
suaq5+XWFjfvRuWzQf4pHhi4tjAT43zS/5EJoP9lMeKOyAOd8n6HIuPCVno2GnyPeu/MGCQZCR8m
SfzU/FBtZCNh4TiWWk1Tsh99qdqNkFj/oFKFj90YBBhw4e9o5l+pmdL5qPZhXj/V1y0Z+Wno/uG2
+ObkCV1Az+cKxLeBsdoxHZwxdlggXSwuDjg2INvvp+aR4STL6kblbrwz+o45n9lHc3h21QXQSHeH
dhC3uVV4coSwq2i8tMnoOIvHseqK6RQumIKq9O1rQKrIVbKH7C0KM7kqQhnh2kPZEbrg0CFcDOvs
sUKFjRZ0N2AjH0DYxeUwspBnMdGJGG+k9w5A56kKoelmrM8cxod8ehjQkGTayae5d9ogn5vrfhmU
KiECepy6Z76xlFD6aDOSTxXnY01czg9pXqugN7ostTpZhCFH9eawmviA0I7PXBZ4NCoT1hI+KAFM
GBz6a5JWOiBTha4LP1r/XRyUjAEKc1/KbCGyqVlaFf5foLk/kyoQ37QDbVzp92Mb+albcXn3ESX1
U69IgN43/N6hAk71HrObzoPBefp7VyxXCt6uxpHnxlvXiBYYlMMPpQ4VKZ/2gFPPp7uWBqn66Iqd
HCelrG50Hga1PL/raLZ7a4RahsAssRiP5AT1tKUzAIdKyiJel9d3BKS/SQFHPV2UPmguQKHmn3m8
169Q6/xn05uxgCfID44UIUwjbY5GX6jLRZd48RVI4j7scYcTHpuouahXB281SMkD3ZMSrzzFsC3q
Fswe7zAqfehaVRczWl2YlPDkUqu/IfNzIDBeBKhuyTUWWd9StmR65viIaCaBpJBPPE+B757qUXYT
bLDRZE/YeTUkDJRYE05dEoRNq1dx4Mfalfarao8QB9NUdJDB1WwoLDSaxWUo3L6vzCa8ZP0zj6+S
eoFRVMTTf3djsdKgQv6w30qhcWjpwX96KnS4XFMNxQ8p4/yKUgwjGfAtx2yH9S14+kocl+4+l2Ov
3+4XGwGvBMzVqzR3Pq7GJI3jV6buQBp/OwFgmbkgXj1Kpuk3zEc2j0yUbOWSKpO7izX/QHGLWlBp
AYBEJrf/yiHxif6yguGh8uNm90hgRp/jhxVtQfVqHKQBOYpqKLhCnS0l7hySDb62RZErEsxdwv+R
jBac0Zk4rwD8Y66z1Rou2fmb0QP8iv61ikAm5XZuRA4I4Mgei2tQgrROzG2N43nRHBs9U62CJQ+s
hzAuYQd9VxeYeBBYVr3VRIAAzoLquJ3RBCDfqBINj6zHgNvUkR6B9PEhnpq+wTOG7W9RP0eM6SWq
hqvdaMc95GX0iEok9hjCnL1vX36uQRY2qzOruQlj3umDrz1bpz/aLqnc5EpeI6qEzDa2Ry4U4mOc
zFdKZT6p3LI792rpO5EWFBEqmf4huQpM7TMvmHxCM2SsQuiE7NwJ6gpp/vGjX2mfsZunUjApNzet
CDFQUejZKt5PK23FxLWy+vUuGdyeU5m2T1BEcjlU9ATBnKR4uPy1CI/HcKfSG3vrN/1gDNkv5wKA
ZVN9AyRfBJdb60EiIla0lKqjWhxUB4RRWwKc9h2mnhxjM6RSkGBQm6aTLujE9NFn1Btvbc+4ODWB
fu5c7q6uBsBsSEcMRFxbEcpjxvS2HYiWLkcvK+hG+10AsDiu+ta4kKxHL9A1UJSdhaPx/ijcEfCJ
KyEXxHen/p7rvN1YEzlKT0Bmbsiip878McHMf9U1cKyXI2/rJ8VFixmWzpA6AHkFCW9yM+z20gVV
DSEXvc7bwyOhIyh9UEWDOGffVo/sw0kirlNqaziwpklqEhdwvLznkiYBJ4Av+FyU7R0gRMzSXift
KqIkRL5YKjlT7cySJ+jNAX6nuHi5sT6YV9sHezcdJQoJ9YjAx6hQhL5PZpycd1WYx5wSNR7Ull6M
5RwgjuXU3imjeEBi6FhdutYdM00XZlI2vXSRcqPexhSFTxTqEYZouP3SN0aU4YMTcLhFLUprK1Ki
dlOC3uVLQSSNPQ+TfIxtChdtk1OujRH/1p5IoekhY3Hvx5d60O3HUOAcNXXUdLa+qRPkx3B9AkDP
vJ5gi0EM4H2Er4ehKHAvfCZnRO/OfkT1Kjrw884otCn/KEFDyfLVcjPrrBGearuCyozSctaiNxE6
2cp89P3jsvyBDuJUoj0kiF/1pxiu9Hlwegowd1JIxFK3VZ1FT8lu9XRMLyxwdapLkMXPkmSgksfv
rbV1TnN6neqcXiGruUf5Do2HyUQdUKx17W/rWhmZt4ofuaYfB/RDTMtL6diDTL3LETkADxsfXkUU
ES1V0KMl+Jgquxa5a9mc2o7M8YRX6b6GISUhKcwaDXIIpTCRVwKgFZ1itZn4Hnw24rgbip2GuqT8
mMgdLdjZq1l2Za66/Kwksp1+8TZrpioS/DMqF7fBEvLtbPEQSIMTjKUTFBiVAdfz6PclnXjwvviz
oaiJypUd4Lbq6YlRW/w8xDjuhCJU0gx540tPX9w/q+qnT8W+n9eWlXHPdfHxpPf05JgkCdylmVNw
fbesDoaL3SeIj46aLnRiq/RBqRvnjVMqucI8Vq29IV3pS9sIHI3hhke+Bkll+YyG7JbYXyTXS+tU
mbx+BKLNAlXejs1xyxp9aI9JB/Y9vMdPgsc+tidKlZkV2iwyz+HDdAy7gcHduHKo/uNiKSsekBDN
Cuv6RV8L/RFM5oPlBMjdI/hRpI2QhqUnTgM5Fb8DZCXdHkePY2rIn+l5SxQIHEsNEy7QDEbgPoFr
SojnlLwvUEjR2Jl6TPPP41hIXzMgiiScWC1mEClfp3mkvztCKZ3MCCU2t9pVto0tZJEvcOZXGPMq
44JfzvR4zKNc8zLfCPgtD/yT0bs27JN33wzx93e4JocVnQq9Kvuyx/O6AhoJoOY4vUtm6nc3VC7e
pPKZJ+BmJpYv1jrNzkwGGmGJ0JSVLh2DnjUx72GKzo59na8PKBXMPwMy7eocOyPnCXA8LcdZHpzN
wFR5FEGA/aYpgkQ8DC+KoNkam94Z8v0iV/6+ApgjvT7pg0V4V+cBtn0Ark/7Vx/n8X+bVMYdnV3I
FVKH/r9Po3KSxu+G1JpZgVO2caDN5D9pNf5AJRJz1KlU8vLGvpseD1VPALe4ecSbpSrXrxFyiTki
UQmQPrAPyZ3MIg6xViTNmVyPPfee7y0ANDQFPJmyBGAvSGfq2sQFYja79pOuD5QBbSZs8Tlh8xzk
rI8a5nrv2paNF4EVbwk2SqHubnj8LN/5X+2bXQDzRMKOxF5L8RDkMZrMZyer1T9GMyBQsRVctiNJ
S66b8Fr+wrNlK4sLKHDi7MuiP+KR/5bWUlstgTZtkSO7LjAik7Z2G0yi80HZPwc2wfXis786R9a/
NN3AqxrHFMQ7AnMmlbV3TEr6hfFLPjMCjWWdTZfUBlY+0PTfKOOtI790SjDUAqT4BDrFqlavI4s+
uwXDf7hxmK/1FoDv+aUrOU2SJZRwj4R3kWJ+xddNwINTcPddqoFM0sli2SKqZ+iOa4d7A5Quj6bb
ZBWMJxb5rzxudcpzGoplTwrS8P+oO2OO98rFJkRJRQBr2F1e5wri23wePrlp31XbrNkmfQv8tTuI
UumhgQ2GCZoGdkCzfspJ9Ep3cha7kYZrM+0abAfcwRj6kQx1yWPsBi0D+Kr29+1bjXTPPBZq6rAo
02QWKWxQiYiq1mxrn87UwHZ4HYGEwy0mvIpI8VKzBno1Kw529QNKp2u98cEmjZ9TQ0qHo3sBasIK
fWf7vxHe+J6KscTaa6i4gPGmvuXBN5aqyuqGFbLUjrTPDDexKh1M9MBkO7izqfjN6R4dRywibfva
trUJFmVoXF6ZVH+/qYYgpR0KdwDwFpvAvyh4KUZqD/6rDgV+28ib/kW7ZW+b99JNKgdyGtftnpY1
2mTqK4Pm/5Yq8hDPlyfpBfCzDKmnhVAmAHZDIp9N6m7slCEdhqGr3PFB92BeGBUVTbHcu/+yhzAx
okBcX3dZytwhdJMaDA+Sbj1UKCWUmlFExJcFOswXqOjDhmDOv6CWey7ExTosO0fwJurFgZLZJret
bCuNzo8r+QOslKUJ56nQ6ILaeU7/9FQr8Cg/BtYlaFY+V29T3uPw2XbmjhCpldm65BKa7wEV6VNl
7mh4gnRu2VVcuyhqUnKC9yp+yr4JOc0EVUg+xD880BZNZXG7fnoCPK0qki5ps5fCHFnPFS+aB/Ic
LMBD7Loin9ojjQ/2AXbo83X+uxmqqmhipBnhxRcEjD80jzSzS4YoC5g440DdL/3UZnxEEj++VIRr
puVp/nzSb00k2kCO/lp24Ad1mNLOYoB4vG4nLVy96M/XvQp+8X1CDQlmhF2B/G9XjIn/XtLMs/+1
x1rD8X5ptotQlvTwUWKFiVoCQkz1Ph0eWTRpbMDmUkSIspp7Kx56MxoqkPMkcTKZAMVftV4C+wli
4P26TEZlJ13+oK2Y5ANzvJqL+1wtsuXXDeBw6TwbBt3ShaYn8IhErA5PsL/sJTMnVwkY6+ac+4ax
F2FZSCF8FSQpNuwhGjAQirM3BW3ztapaTyeJMqD9c0YV6lpvVjh91XqjSDNKjTFotwUC8yt/zmjC
nXCk3IeC3ZIOjgFdkn2laADeeGUfVS+9BmRsvpFZrk/RF03Nl4T1ujQWMjrVsaeoGBirZHKVYwXe
UO4CbLwq838vDa6tLAO87lG/VLB641PvDbJGGGKT4/+ZPDeEtt69fHiJle2Mm1Qg7f7+SnSiRPpA
jSrkzD9XSKU88SZajgYHPyQHGo3spgTaB0+i72ZLDKxRHHFSTf+uAM8UBW5MR5NG1ZD+dNY/EPlb
pbxLvWPjhONmosW7Kdgdx0KdMCS1LCGoXOsbstTm4CS4Z9F0eBz+poUz6rT/OlY8Y/QNXqfsR6YV
M+7XrmbQSYrghcoJT59BPXSMrf2XJX2gaa/QSfeaHuAguboQlpTAJ/fHOiFGfUxIIMW7A4ktZCJE
1z4WNQJB+cjUC/bFZuIUOISOOyK8cCDF11stlOApIC9L8fuuAu5GDzG0/8bHPTpoSLPEf8z70uXM
7OS3rThp1gNUZ4mCp/rB4Baj8o2mcEe8i8Vye214ViwkDX6rv/oVgpVhbbXOg9tCoxTBtFgAeV2B
dNHZvIj4DdbyK3mRkhUyanqQozayIDuIVS5CU51/P9W+LFrzyNN9L1JY1mJ6olc2jGoINuzOsXQe
y0xnkC56Jje0H/H/Pp+W3krSJNVIW+oMVRmrr/eqTJJ42VdsvuENzK7at0R0pqZRxRZH7WEmeVL8
wbvxRUmRQTJd8Ot9DCA8ivAUCROS5rykW/JUW+tGK2iHPKMG4mrMWp/QBDBvE61l4At4sg6xSaRI
HeChR86BJUQT/KQRlEBttfevHzFN8psGrzmT63/kGt0agCB8bDZGFs6y1I0bO1v5A8RMvWTuCvyT
TuPyfZ3yXIaNanSbNNDPYIHzns82/8cjjG6xmjP7x8a+qKHZuXBnwUt/jMnWhIn51TvE2Uli/Qj0
YGwglGutdP+SUmgAKsSzT+Dc6dqVQQJwUICx3YHzQF/ImLqkWuFLlHnQH8pZ30pnWDl6aPlb1wZI
SQFCO/OIHZZUop9iwjjQXPLqhn7Rwb0rKtwuBxDiFJM+qqP90bDtYjoXcU/a0BM6LuEB5dEnrc1e
rCFM3DWrtXX/c7+FJLdYhDPCV311fz8dRYsa4rO6d5LlklfDmmw/gBO1Yalz5mTxgdln5ATvhiPZ
veQLigmP2fjIc2WJS+mdBQToeM0JmK2k+lKgrJ5DvR/HJOnS0Ptet1zQbHebll91WRiCVFqTwL1D
Fk0FtDso5S6k88ULJ011+aiX1/HAtJu4r4De9LIMTidCrnq6kjdt9VvoVDdKpyTckD0N12pzUgML
/AKJNbD6eNgZqrobWP1G6UP+KziR0Lm3B+Fgr7IGKsa8bpSox4oVypx7LRwNnBRXJAL+iq9lSBc6
Y11ZSWEgtoA5w2EaqHDqnTB9BCPH195o1Tkh+oHsAGJnyCHaG94eexkhRI65S07ojtw7xiadv2Sp
zlJwoDqc+44jme8D3eYSXIF+ud5o0erTHt8a2W2ZRdU0Dh62CzRw93WZ60e4gWiv6fhfWw9QMifA
vSEPKsEOII9/GtO/88ChO6vwDxJcjTC9h4tLI61IXo2TjLGRpYHaURPs7WkaqnGiC5B76VJ5brfd
7WFLRaXli9dJ/R1D4GbOiG2iJrqLoEXsSb/cIKseEaCs2tTWDcrOZ44NybvIpFgYlphKbNmJ0eFB
tpjZoAY2RItjmxBYDy45lbP+MSUoHN/w31aqPN98p1DXve0BqRotinPg+eWDD3fSzp5tZUk+1oS3
tvyIh/FqNfLB/MNNyYaKAeNqj8oADph2lyXSCeis+PhiQyUbL3pj3M9/yBmc5oagB9NEXjCjXHV5
0PLvf5yNCd7+12vI5VQtaW2Swxp6Lhp2l1tJhGmmQiyZItzpWXtCdlOgynxGNGfIUTqApyehl7Hp
Hpm3aiAQXHNOi+k4b0YqbABYxol8kHM581dwjDXmP4na+02sOzAzi/+occCa9zFGsD2kjhgJo4Vf
vpmPvrOYSzUXI2kQlVYiEAI2L1GekEuBPRS672LnSdQHqKCtwg7aRL6RaaVzkagTOVoPnymVTNk9
eFfse9nDXCvjlYLimNLu8g3DSsFwACV63snt+E/bZZ/GcXcJnWT5rSJMKLk1VtqbemjEuJzz4MvE
+GlxzNXV/MvCVOBZHfFZnDQ9rLIe5sI9HAor1XQCe3QamFyAy5HvVBNkg65Cp/NWiahWx6rdFXIW
POgS3xpBBckbzc8ns/f3yewlFGGWxqGljZBijlEJr5jQ3yvlxRFac0uauj3HIlxOliiU+5pRTjf5
fAC9XPAPORCUxUXDXAs7j58WIn2od9ZMxBquwy3KQualNblk8olE8ECaEMmKulsd6It/3+wBvcBH
b+OIrMhWGrZ0sdZoUHsD/bT50/zXYrl6xQkqiVmGTlK0afBNgXaf5SlZnKpZmCYYSqFMy+4rttKv
WrM9feiywDl6N1m9FLZYYAx4/lgiFue6FqDnz+2Gtgu1uDgdlByWIkbX/jJOzogWSK2NJ8PTV7wn
yRXn48SDu3E3YN1tr8Ho+/bzPEeDc01hVpYxWfHDegZId/XFg9q/LptMQiq6wChX1vS63RyaANYK
WeFBUlBzbrEb0zM+L4WXF4OxZR7h3j9CqDwSPAQyHulqkaoHDN0h898/5tAZY0GUtRNWSHDaknhF
kGIDkKy8Wckq84L18wIWRaj3Fb6zHShg4KrLE2OwPUMbt2ZQF6UyPeROiuI5kLFJy/uCek70DjRn
1izxcV8eejYkjEJCBz80W+24REfJ/Otx6Kw1Ys1OTi9XbT0d8d02c1gpkTyTr4bx8UtkIKvN8TPG
UuKoRcosuT7T/JQlQANxKJdTxs8xZyIRHO/lw9Z11c9fgCdQTU9l/ruxr9Ku8lArtVoqFIPYY0V4
haASLvkB5Ll6sSNl+i4IJMHxMG7cLN/rAdrAoiPygBv7f2dGF6CEzNSR8vQg+0+WDw+gv4Z6JsQ5
kuIHGWrKGM5i+jUVxScEcAMR6+lpeEF89nmZSGgl7OHua8I+xvXV3roLS4/xKAxPoFGGR8oT0iIw
ozO3WBONjG0tAiHHPlLgIc/AlqVlCgeqJj7UfLITDMTrqpgNqEwSr6Ui86cXqxQqI82PPEom2LUM
UdaKGrCp5Q33LhHwwaYunAZYqjxywzpIPHkxl6KXqqeB0FFq3gRdmEj0SOGj+JgK1tju6fYRGtML
AD92wImX+x0IcwZVSU42XiRN/bkC7sRXOnCb23KgwHHn4RCGB+AfxdoTlbhuMcNpHCCzB2FNVwEf
KVmff4jxCCwAD/ye7qL/FgQM3K/zk9HzKGx7HM1R476cXAMc/hzI2WkZET2Odrh4dUzaEBhP3Gq4
DPCcez/eN5DUGCYTmR78n+r4TDHgHQHCbYqJil3BW4JtaXRi04MIqejV9og7qe8712lWLfvXqJXz
VaN2f5GQHU4ceWc3nT569A1N6FclZmBKn9gmWsvX0vr2rCkN7TngE792ByO3DvffgRsgkqogITmm
Cgpkk2c3WX9M7UTmuECqoIXZqfuKFuzK2KjIh7K/lr37eZVENHmAWQjyysoYMlUKy6QRBPY+A8Ot
F2EWK5z4mjP+WweQRX+YXWLsSj26HGFkMbjhuoI2hvgl5TONjKqfzb3UWbb8hqDdRAFGgkR02NqD
VRBZEO6ZJE/HOduZa8LAtNLF5V0R6VpJzVkhv9WE8BnNVP7u4Ecg/ok1po4yYt03gN9KhQnA36xR
xaAHDG7FFV7XFfOU4UsUjzZwuwAWScdbzIPFpS6JJbTJC7W1qFbt5AV0hfZz95t3fpKvtRbTO/Bi
73jLUFBzAm/ASPZe67BoSHBG98dWItU7MgN90XBXX9dtjIG4nsoJR+pmcMbgKmWSiVpUZd1wJkyX
lzy7UB8sy2NvhvKEIrlv1f0/aBh9OP0wAb90EylNr9ZU7ItyAWINgnqUFerciIX9rV+1WCynrZSW
NSlT36Ey+XltmsUO2C6JoV3psvj8X3PLjA1/NIibuP7IbbuO/1R4MKJzXGUtAvQhVJvAUg6XaoUs
zVCCDRlf2DXlWdwYFqGiBZTN4UL7D/4df4xMsZDUF4PgfJfwbL46EVq1y+gH1kIlKULax5EVXQaZ
JJbLyUY3Ub3EiC8MtOEGJldAQTVFufmTmaCJAgGgScXa4g0WcWBdEhgZNztkqsAIAaEcQRMdfxcr
6xmRDDVd3kW7urRTsfRtPjv/E7jRlsQuDe0uCZXytZTkQ2H7Nb99cz2vb7v6fIRD7EZbiYDu+/IR
I1DApt1YMZ2yQ+6C34dHt1xpoHIz1dOcVVsHJewkM5ASizCirXggFtm/WPRLVvyrWHitBvRAL35L
+7X3y8R3VWrHKrPoVconDkcgW7NgRGMrQ9lZDCisPVF+p5BNNYwvhBJ8pEnQ73D+XUOvLNT0E41+
QfbKRh8un+3KOx2rHTj8coqL66WLTNXhmnHBOQtMabf8gkQdz4hHmCrSN7FDrVGBxAyxSdZOp1s5
A2lbd+8elTLAoMxN3k9lT/le9KIi7FhOKjUKbQqj5hNHQB+3TY7hUTRGRPTqrJ5tmkzD6YfN2DnR
T6xk1gQ33FkiW2GTB8wSbza2EOhky8bv3UCOqtbcTCuYNzyuImrQmI7yQh7mpwu+S7s6ZEmlLc3+
HC5J3ZtRzsPubE+mEWSMT5cEik8/57UsFUm5z4FPvBZzDW2JKRzrwCWyzLN3VrRb1Jaa6w/9bfBx
YUrePd7tM/ikTNEkZ+nOgRyLPWImG1+1BiI+ULN5pwFn1/J43rbb68ZGjdGeusmkO2Iymo1hGLGB
ZeWMF7BZu4B9gLFH/04v3cQ/aa6xEndYzPPPf4DNG+ZFsBGzL/uigCG9xIbzqA3b1OCoxlmEuIwb
pLXqczRbtauQOh5TuxwZaQTOq5On8qoyCCOkHh+YgBclf8FxKLwqjJNsaFySwWarqJWbHMX1Y5uv
T7benTJyu9Y8mXk1VaAUObFXev3kXTs+6rdngorkjLI/d8BDpcXTepQ8I53ODVoikt1HM9G3PnU3
hnWFmdUXyD4THaZuJPSE+Zt24X2ABTPK5OINWfzP5fRx+wY92DRKeiqVRkY6NRCXPLjXd1kDxDPS
kUS/0WgMwfcqp4LvegYXeXSPBQmen4DlmlJk2V3kl1slaXD3rpPQXcPo0XJ34SokzaEppFApEwOr
P4Nb0KwPrUjbso8EZm9+RPawBCbfy22PA8LL/tHnpUCrrM89wDZnRtEZlLuWo1QZ/Cb48UOt5Rt/
5G7n2PJggpbWLcYr8n5i02W6T6B9GNsulYSZVZx0XXOQRKsRnnDoYWg985kpI2SxRCZJuu8/9Ahm
i4mbnP84IDaQTBtcZtsbKNdnxSkcEoh0lpoO9Vs06ZOzwoePUqZaq97Wg7ZpUiXf8eKD+8Q6dq50
jhjvNbnH/YpfKrbZkv3j/vMPqsTcXgwvV8T7wNAKdviGhkqGTmnRUgtYV9DAbmMZNQ086vmAN1iJ
l5vXWBtWUBDASX2SBVGQi1aG6yKiikRp5ZWD0PDvA08RhDopN2rD63CsCCEqugqJIkkKSOIH6YpK
KrUUhoUYE4icSQMFZjvGQ83cf8XQ58rx/yEHMiirwe45W1oLV+qn3hnVkTt61kDE2O+FJYPiafHP
3UUrFItpTn5R5frrm03Fuqh8geuzEzjDEzOFuriDSt2Rmmbmscffw/M3PR5AmsAhzbejS5AAFQhn
gLP+rJTMg531GMEixZgG6DlVIwJy7EHbKpI3J4JfbgTr0l2/gwEs9B3uR6ow1UclmfZKx+1tz5jY
45Woew/F0ZjqerlCs6/bMtu2K6DFE/qFPpLPK/7Oe0EzEwiwWsXOdDV8t3hZqE7kTVu87onaDYFw
GOoH9oeaLhWHc/DSWNvOQ02jseCL6E5tDl4eF+S66JeZQqVoDsv8qdT6Ea0kCUhrPJMTnccstr5M
00JVyOCB98paLZfaps4YDiatvImfac7tvIe2aPioWxrRHWC/iFhzYJbdXJNemjsHnJ060bePheHZ
ll3rEQ8u/YcRuoWFBcv8MjbTUl3FrGwfaVb2RkYu4e8EcXk4OwJwh4maiTDpFXggxIBtMg2Pxq2S
KWT9LE3p997UgYs3J0l+HmzgdlIqnPCM02bZ9AH0kI0f42qn2h6fXBU27UKij1pCKANTzkyw18wy
2F0wYQTPkzA3nUCghpqTba1OOms2uKuZ1b/gmReduvuyWMYnbTRCtaaNzZ1ajvSbaElOWiJJzNhU
K2uvtnmxzFm4R6a3+K4I3mnw+leNsoVPTS0EFef2h1hAkPLcpydT6PDvOvuyTbF9M1RR22JEY6Vu
teeItfoICR1RlWc7xF2utp+2ghmNnT1wD9TzhF+FvGZDa6mESpAWOH8z1rytaQB0inXYQiejyxGh
/JVpdCqcYrDE8uNdRTVAvl7A4AzZYL+gm4eZGbkTPeqf2AU6xOulESjEPXekbGRIABgSGZEFtkmZ
kbgfLs9wAbl4frX3O7OANSFyNSXvAM+GOCOjYaNXg6t/cGNExuGY+mE3UMG8SIQ0UmoQPL/yCqfu
EcqMoNE63lK+8PS/Z1eVh0f565mYsW000Q/kgKnPjJM6sEYMnCQP+Y5iCL5UYw+0xZB4awHeqyaN
AOYY2Mlw02koCmB6+dNN0wo9wYV+dRI04Mw6CCrhGaJfuFUyw5zcgAdUhPavaNiwEODw8KWhv+p8
9FCrTpyiVs47c2JbJP0NY8Z+LHCKjJTEWPSmgUMRGgSv/ghx8SdE5xej4TxYgp+HFFG91d2wfshZ
OOBobhZ6nAcyEskdWMIc9GrWTo8xAwQ4y1fOhoQKek4A1F1YtqUbAtJeIRt/CXWcA6XygTLvcmP4
4/L8HSLJBrZ/mkqtfkENE8oZkr1Ui27xSqL3SxY1e3JD4qSeYaIgGHs9R9H+VXHKtkQ8cVLiz3dH
oEn+31Ro0BPvukKjL7tSqrEQYzAnA7Gv4lB7m3tMLR9DFKgnl1WZvEV3cUmATG7r294sJCpaAg9m
Nk/gNL0ptGwlfYAJawrSHW9lxpAXpa7aIoMi8PE6Qj+Ez88dh1hZsu/1OgtBGINnFiqfczxbni3h
GrlQTS6hj6PkKlNFacKZv6ZapKNColRHiGst2U0PUvJhrMF4G+cNRgRJta48DZN3D8qyZzey7Zn7
knb3euKWu1RqLo9hOqywQNlxyalHdpDlo8rjDf4CDkHLBmd6bc0D9uJkRgnEWzTllo94GI5zvPoN
KdI6bEsxA+djiKZrjU/O2n2J4RrNtu42HeBWwKZfEKr3nlpVRSr+jPOc2SMO/IxA9069NxHxpjjz
0R0z28X28A8pwrEyWk2k6RhhkpeK30UtO19F7EYgR5RNkxzKy8DVhT1Kgnz2Hf4hcQ39Yt4MYIXw
1L1qrKtbsT2Gz6AP6scLAtj+T24X1a2oglSlSxWG0Tj7l/+F4cpvh1Q4Fk//wmpaFuSee/5X1ofF
atRDb6frcG/MspuRd9E6iNeFqep7/dYfnZkHXA0glXKjxJM6kWAg5SoG4plqLBR40uDl2LPXKidL
1aPlltbVcDsx8AWg/oR7GfuL8R/NT9pz6WMoiCPAMWBiovnHQPJ5SXNKDHivAZySuDXjPeduLVeX
/ClecUGlLoSiUQHyjPgXsYm5KngLxwC2LULe+y5jkqpd8+19hxp6YMd5EAoke7zKUsBe8Y4AEUwj
PWxyzkBPJV8mDbkbRl7nL+wyXDg5hR/W9zDCUwlEQF3OzClZWzcIh5awBCqca+8tUZGyb17MnCfR
o4m7ZeOM1mTQaGMZfeaEn+pYOztqxrnGym8nDEHacUiF5CdCcD6jbOZ0UOK7JCnFBsi5WXubWxxw
Yf9SCqFb5FOgiaQEPyeynNPiEgA/aEAoEQKdOh2IPNNnZIpPITpeT9XXA1iTFsFpfx3jdN1Gnzy0
qQcOpokjC/7+TBPpE7NESur0igzTtOrtSzkZx1a7WYjUSzp3y7sI0C/QQ7jBZxLwRgvwsEYTflXg
t8yf2b+l8Dj+uXrz4RdoAr2Zm5OYSJwo1yUEqJ/qlIsfn1XWUu3eTgorShZawNAgBfqUYuN54JBv
vHrmsu1Fpw6Zjv5ol9XO/B+KgH1ytrlou1RPKa4mSeJ5VwgLKx2ldFfNiVC5jJYnj6WGcTevoSFa
t5bmS/McMy3uhOeobCG8be8gd7BSBdhrkwmtsXRzmERwY36ET7+ui1y/XNKws/aKdza3W3x7NxRO
gZNtWYLthDLauKZFYPlhO4JI46bsnY3rzmQnOPje2dp37zoUT+smEpu8BdBVkcDCOMv6TLfr6HUQ
Hr+YyNGQndOkS+Ftj+VPRWlvoKH/hVDyqTBd3ozUW9CPzspj6QVwVmb3oQBK6PCbIYdzhG4aEb4h
/QYf3eTPECTovnZx+m/iyh5kI7GtQbK22CBqUsy9vyLVz811oMRT17kqtz7ai3FjlGpHYkf7lmoj
bjRAMPlRxj3yCiBTGWGBIjMDBodJBM/aiaK3UsZf1jVj3jcFwIBuDQzsIeYVHk3FCrVYpkmJhdbB
522dZ5GRH/vpvpl4iddJPhwkl1ZeuslDVxJDyQJZF6ylFWABkzKAuuNw4PM4a+uqtkAanGGxeH2w
QSzWw4JtI3zagNIz2TEePYjYXtG9Oaee6Yb2Zl79z/4W2Fs7E6U6Sh23l603YjdketJRUS/YaPp2
juZEPg+SeSx2qqJIEssML6GNMM8VAcdSxxfwt4BfwDLX0c/2YRv+zAybX5pSBBlT/HWLcXh7KeHS
D4K36iOs21O4/GQHFjZBUdT6Ai/PfD+MiuxzP2cMZqjiEm79Bt851TA0mllqhLrJchjg/jiaRxE8
FKkGCCQ7j/ongWlm0Vui3oF8QyA6pHqUw7wqvmvarkPMH/ojfWCymnxXLEeypZA4rwOCoU5ScEYD
8uvV92PvoVN2ofNFP/MbfGwLxnHdTUcJV5+H5XzoqVyTOXoqy0hCuava/uRtZkpIETfbLEAyk6gu
MOhXXc7LfYi/HXPWJqHyZMqlFFO7N9YXH/2m3+yRQ4P/ztyN9pmEQU6laqnoKjuA/DRo9G12xGx/
LvRA2kqwhpi6kXAHZKPJRfT3euD8qIAbuLdis8QPKa4m0ziddSadNhrGlzYGbmgTv4rcnOOK7A1H
DwlkPWFDaufBGHIhcS3qTj9n5N+gXwaVaUjXAVJBhdvflkKcm/egg11NTaV1Aedyrh93mIlYdXto
wcAs4aA4kyOLsKlyhglz7e+BnYoiH7uIVgXpSqUH0pJbbodn50d/k59OyqfqNYmVw60UkQ3Iwhku
fo1y0U11yUPFt/zvmWbmwXjJzQihx3SFgpXbnXwsCOdS+rVmZcoGVajgFLa2XVLm+lwnrv7EBgku
A7XVVLly5y2QkRuA9jkgGkCXbGTUanzc3Cix6c5GaSr8p50NZq496cfXUoUCeeVeAbVI/CDIjR+Y
AyrbVlntW6aFJ7PMSSZOInGkD2msUnuQ5u2eHDC51xa18YIrfuvPWoS8UMA7OyuRqqP/o2k57iCq
0+fMCL2Q2doTg8vpBEM9YiCzcASuxyi4q7ReISWyE06IkF4ThmdtYvCO5Hfm1X64yDflduNPx3vb
Yld8UoUKOdROFeKOg0pNnURLXsLP5V8bcyKRDcZXZJOOtLbOuZpJ5Myu2c6VegVtCdM9OJYCF0kW
TYIpYw81XnejZU9gHxk1KECuCI5mALZ8fx2OWr3znGw3ZOC4mbblhGPnduiWiJHdUC37Jma5tiK7
9Dq/nNfUlV87LxNTPto8yj6iAzx1c8QUqNHrP0TYmzcqbEGerq0o32PkbqQs7JGqHbxfSqYUQTI1
HF0W9ldijxKimjh5lW/G8bVyflrX1VtI8cZ1Qz/XR/Tf0ijK8fQRQeSuNuW5XytpySBQkXvaytHq
cTDSsmsj/W3MXA5qjxkgo6vMiZtFlAnKW2SM73ZJF8dwluIS1SSdVAHNCXmaIskzi0gqHAZsi8OL
f5IWa+6eF7tte+I8B0mzwj3wkhLgjS5yxrZUBZhi3tJBvL7hWiJOCrGPmj5pT+JjRXWZjvdiEZEH
yTGoG5uG6r5A3auXJ+RWw8P2ymXFUCgVN00sjCrb9U+ISHfTqjVEc/eGP5wmZoJS34lcDhzglhBg
w7JvDMwja81A84ADv8QU2uzvMTaLDm6wCcnfYhxS8O4tCGwp/LXFThCTBkA9EKKMCAl2vuaQfn6O
Bdn4v1x9YZmsunXHejEkZOf+bBWe3MiwwCmKi3+A0JW7RAJKOMYYaIULB9Wu920i5uy5g6fT/rHq
w6JgOEwY1TAmWsaLuUyjOfBFWENMGGSLNCSoQ9EgDregcS8g8dXtLamH89MtAW6Hzj/j5PKouSQa
FUdu+3R5Tb8ajVq4U4Dy843McG/OZ8VPmKXHktp8lykN3cd6774yHuc9VDEnGfWRa4A48JyEuH4t
nZKDgfjfr0ZdWCB2vwzSo4fRA0iaTt1XMSzgV4Mp9e00hHUMnV+aBmLknmnDGJtWE5Utdg+6r62T
Xxj9J3CW1fLo4ISP0YZQnfGeTssxE+Dani+1wpkdEAOZ5WXsfk/yhHvf/ZSziQs7QA+5HTu1ibAS
jTlpvdSt/PrdUiE3ZtOBy1rg1jhl05QonmHVHr28NoHFGaWTQcsEza59CS1eTFfU8VS5Sq7Olypp
CMxdsZe6Wk4bBku+0gJSUqksn8BLduOOx6rRV3jK/CW+NbleBxcIIkCz7VyOuvHlvFyjUub1KkD0
EUb0SpZf8HZL7ri8Xq3beIYxY3HlpMrhKxbOp/vufxdCHUp/Sq6LHaxSbRRjks+4xenOp54XWRlC
dX/cFTys85SptsOHpNJlSiY5zvRwobZPJ3DdXIYohu516Jx3yzuTsrGCpmkihhH2v5JBNALa6gQt
Nr698S9Hz6b1CfQRA5Xg3WohukDZjrVNPv5BMZ5zLqaJUU5WVawXdBh2IjXhqQq28z5m1A/hwwnm
JuDcdWem9D/r/oXULdDLyyLCFZ3NCkc3Ewkstl56Qrd4KKAFWlO4bCRYFdUPdJ1YG5qav4pN0nfV
Ke86hEqjR9UqppVH6rhMmjpQFDY3JIKTSY18qldGgKpxUGWcTZCYcfZCLYhUUey4ozI9LDc8geBt
EDeUgvxtYEL0nQqyQP0CVFVCaTdq+WGQv1e3hc69thdmVPGvLNnkdCGbie/URP7NSXIkogL9Y915
0vAnyELOLFHC6UxazyeGsBV3uaDgfJIG7Rz9+7ek4DdVPSF/T7Mq1Wl4EzzfjueGGer2dS4kWkgJ
MhxifedF19rlA5E9xjXojKNJAtdaoxlcGCMqrnol/ttfmCiWbs3IHKPI/8ishgASL14ipnndH4wV
k9r3McstTmD4nKnmsRNSMfj+VW75bgXy8YDDeEfuxDEmHbaqTe0AgrKyHxhHp4NBIpnTS/y/OFRW
c0lvH5Zkb4jvLCfj6JYieWYTBhn5Q3NmiSHRAgkj/ws0QiO7pfT1oXJNfl5VCG9Cl0iWeRzUHfQ/
PjEjjz+TbuYSuQgveRsQzFbDyfHaDM0WLRIeEIaQmi6AXqb8RaNxo1gAKiekdtP+ImUyrbj/62Rf
uYRTpPUG12iooAe3ZKbUTPZf+XNaT3Q7SkfItZ+CO/xkyZPt0VshERB3Zqgpg7YnJ7HhgDITxF1a
Y8K0eOENhbpTs/4sMMNY/j/B33b8iThATv2HKWkgI8R4eTCBdf6665GTV0q3WwmMOfa79XaP0DfF
OsfColVRP2tPRPHKeRI/XMV36mrowyYJVnz+mmp8zEzbB9OXFXv17MGjn10nWVszkPKwGWthAkpX
CLeubykM0Uh+BFGfiMQHdjLh26J5Fh6GuSjpyZ63oDd7SzZ+jn7j4t5tV/wOoKc/i7FUxf4Gjp22
/P9/Z2P2/fc6b5JdDRjRZW0itfHxzuGrT+kJEZ9DmxwdX4bwVihnmTH9Hp2VsaKpGR0aAHhBy87k
eBmmNw0vPw/8mqRWKgAtOJvlJcKBGeR3hJYYu+mX5Q5aXkWNy4BwS+8JkY/TqJ7OETuPTdBAabpe
X84S/sDdjoUcROZqltvHuZw7ohVD2ImptcYYsy0jwzrLHPnzbQe7XqCX5b+6f8/KVFrSxXQNSLwZ
UOcqjDJtQqiKou73Lv+i0GTNxmE5htcy8KQkh7qlmyMWjbCHFZIAPTjiXbLXilPSlRJ9BC5N69Sk
UWna4heIsz5tG2+sh+/qPLF2Y0u6pWe7akGR+zG1yUsOTM5bNDKO0VrHXqW+hhy1be0mYfCt1azZ
pSRYvyo957EuxCAVM12jP6mkl9L/AJvf8DBbr486M0//hOQpjBMdQ7nAIyaGVBmYGzUovYPMXWWc
WGMUf9ttWyv3M6tB4VGMbJ3wZZV6lQAZXV188KRcnvTIlbUnxzPX9bQezVH4K1JhObAdISJuzFqf
n/AuDriYv1exdFDaEeZ6IFXBvg4xhakR0/Biro7zjlE9QsFQW6yWHwmMtrlSPJg1MNAMC0EbDYLE
WoOqPA7VsaEam1X3Uj9LTcG/DLrY4oy7Qes/KOfa4huQbtwsBNKwQICpCgrHzIU5t0XJRY1+7qwL
mNi+GnL7ObSFm1xzv0UV048rpWnzidXxOMzynluO/qdl594G7oAs/70dgpUkrr2vUIol76hQMOyc
XOibcqQT/bHYvEp3mSS6BuBNLMSwVcngO0SukLnA/QqU1TTn5lj8UljKe5U6yCclpaITIwtqdsmr
X0pftME3i87AXLLX7Daqqzxb9hwNwqmaeMLwv+GOaL126KeenDOwUlkFTu/H8GJEEk4AmZ7oUlLS
GoWoPjrCjSkceY6MxE/ghPoNlekoHoS1Oz8XYMMsKhn0UPu52heqSef/KMiJFFQjdYK2ivTEa6F6
R/CsOypQltIfIRtZSeXIPs01HWgDB5bTaKRpWgTy2SA8FopbpsZ50vxLWG/AEvRTu4HTf6/X5+2P
0xCaOCOyOpt2OiN/WsvnQXmH8wjO/fdykzcyR7DX4u6iFCBli0oFtGSn1Kv+1Ze9utAfjUSrhSo/
V4A1xYzxFzGJH1vK7YhwFw8MvS8yM0rNj8/9aaB9CjEktriXOvTduDStjTSkpVKCvFWvQyCRFOja
xYmAXg+95lsKK2npNoQQQPPmBIcCVzeplswp38OZ8QElcb8UGaslRNVIDGNqdo+XIFq5PhVtHRvt
5Zrlp55SDY5B7N/MVqlj75Qpyl7dloB6WnBUfu/jmpEv3mpm/MBcrVRqNKtTYlSwBVjkfjXjJIcz
u/Wl/XMmfbrIHbtTIpscFQPl0TNbRMLthZGvKrmDJ/9e0XClMDLV7TUZe7D9d9OHyGZNI6IYwf4I
D00hymsJtqjQUFbEPsPRXi2Bbd+G6E+sR1VAgnoOKNZ958X9JGZHk/qSwSjN6Ja2xv2LBX5ZqHAN
HyRGlN4iVSnWn99w7+j/5F/Y6ZjScvrwDMJlHalKodEv871vy+LGGomkokMG2HtdX8YUBQRJDMod
603sZB3eaE5r+E3pJd9Oqs7RyiQLfB5GlxpQkJ77zwCd5BEBfpQ8RocjHYNNohMltSZZQX4t+4ok
okTjfhN3I9NfBIsheDBohIbVbUikK80YNyZs6FVa8QZrs/cOW2j1suKkAkExXJuc5JzWwV44oTPU
k8AJvcR/qhQVSDN5N7xttZ498wNDMGy4JUmloOeP2qM7LSJwdhCM/kowGAkCXDR2j2RJZ9L/YscZ
PLkyfm+63HBQSorMPNrRpav/QgIcibW/GfCgladBXQ7yiPFI1wbe4oHd6zTKFt5izxEC7NXLbJvV
CQJjZwqfFJEpib2obiWAsSJbxKa/+O4hONKYeuXyAAwVo7CfjbJHA1TynWciIvJ0LfjHSTuaa9Ff
nbYdpaikNDDBMU9APfOLpKOJsJv4ZHkrW3OPLUXeI45ZXCo6HjrEVwZfJkkHKyg1gBhWkbRoqKMa
pJHhdiwRVL93QKlJY7JU8oAvwq8+IzNZ4GdZqDt7aCse5GAOEzo3cOhBKSE6zfAZCMt++MY+MUST
KOOa/5h6TR6lCOU7qKxJdrfhArn5nIDMzpVFCcvHIlxy4KtkNREL9iOU9jl8aSGSor4rse7dR9yi
4iX16oGOcs/wiT5cBBPu9aV2TBNtZ2FVBKcwwZSh64nxChSDKXfRqlH84RSjl6CS/ayORPNI1sG/
tUTNKaGFZqllOl+WI+fkx9pZ10UGyAlu9bxAAGUWSwytba++uyEQLdTwVkrjPnaYTU5K+aIvmm0W
WrTMtwaZPWBOjCYI+mK/rUsygOvC7qzTdhcyAL08MJ6luUKBeidwznOtBwHDvVqrbai1eqhaOXQd
Q6l1qVdeaOtssgE1ycedDFoPITzKCRTvIwNsnrSRFeFBFYUeWj/4dBAdVLTJVSwcfReB0Z8nbszC
+PIcJ6kaptz+VsIRa5cO6wNS9qRNwsVel6u8fONrzQn4DClWFHy912rzL/kna3mq8F29q8VQNorp
7yeeMByzGNsNK83Vo7n+DRbLq93aHnQdAIFJXRMQICKzNEbp8MQCT0egvNdbHlnumIg1l9N/goGi
3/ySND0uIZfkAG4bTWmfyDmblmhwbz/63JLosqcdSF4b8SGlXqjc9GmuD24JVTHIinpb28zjZ0Wt
vvfFZR2VS2g9uofIPw2Ra0N7d+Cf0Ke22VDOuq80Yh2fBH66OvuJw2Tzx13CEJSumbHSqBzWK8Zz
swVn4mJokQF7VslnXmwsaFQx88/wf5b6MU9X6b2xEouph26xWQCR2NX3sGUMh4hp82cXcmaSxqOs
m+FehJVN4sFGdAgRToRoOF4FLnBtDNSd3+vDsHn6F8S6j4uONFHukPHfX4QP3NpBAlewWDqTdXY6
hXqGWIeHU//U4f3mDh62qfQL66Jmf98GW/lP7lJBbrQC+OEGEiH0VRZR5Kq7xHqqqegVP1afgVuy
3UXmpKfHGMPv7fvx2Yl0hT4qDd+za64vHJIewtLjcVaWHKQIdAHYibFzrdTLgzgJpklmLtlF2q7K
V8l1W98/ksVD38F+y3eQUAHA/xZoCyBrbwfV6fjQ07cdHbewHz8aRg5xRmwyMRuwArO+M9o4/YPV
CqZ+BntFL9B7CPTH6khS1FTVtOafmOJ12nTnTdDgXOMly43Bmj9S0XhNTzCk+vrQlKsnSyZaimNv
4r8yZJ5t97UfIryi6Em1tQgUiUQKmhAYeWmxZdrLzrduuK1La5690nD0Rv93nUIe3H3ZtzZZ8j8o
099iZm9IkyoCRGCAjxeAboXdsnyqxZM8Jeg07MpCs4yhglY+t1jSQ2i7Lp+Go+WaHqqBIK4dffkp
Fco5dU3MOSNxVzfKZc48pY9gm9ZW3zJS9je2vGWLR4JzZjxcWCFU69cPG4tEo5OVXFAPbCf01u2F
WTxBssauE+F8WjirwTfHHZLIjO9qhbPbOB/Cj/Tj5Q//juXyytP58lCiq4va8KKqiU3Oh+MqWIws
98vtoCkktQG24Dvbk4jb3X+8cR3Sox1vPPjkIsZGglO5wM3ox8HBcfKSsVG882m0mkWBiczPS5KQ
+XNxrbmjTBioxb1fQoT2XqhNRt6wBokaUvHbudseZxNUMP6Eh62rdrvqvbv/ALm0h2EVfDUr61Mv
SXVa+Uito3OqLEGCNWgIqI0KJ234oEUG8qCkuPa7JZnPbQXKWybru7Ro2lVbRGGAANp36pErEawR
e1HJZeDluUt9EAqyGs9pns+X1zb2AMh/+FRfYxznhu8+PGjcOB+N0jTw+oRH9QHs/Blmxz2p9MWL
W2mMQORxP7sKRGyiGSpkhag1n6BCb25YTOnX0Oll9aQEG/56PXrdgRPpqOCia1IOrBMpEukj2CXu
ofCSYB0/x69ztG+k+xzeLQ91oFKD+sKvxc0fuV1hwCeLaVtEFIfAsvsJiMlXZmp2SHsTmATRQkUN
dC+CzVzuCaVg7Fk/7CMeyY3LdM0atjdGMkyQw5cXzrQjSoZ4nBXcmri40Sd82utey1S/vevIacOd
UCwu2Aw0OZE324S2Dfpp3PsROePXUdJMxRckoHbs7aMicXHarOnF7NLymM74eP8P71SChdH1os0z
4quwuqP0LVTdHf0Edl1Y/G6bLED9yN5sum3cCm6RJC3EGVOxvEJqErURw8QeLcHNhtJKeWFqry27
xM2SCti9ikoNZASMplNvXPPkLgegwGYz7s6zWeAaOZoE2mpLUCK3WLyVEoSGIQt0i8KHcqAWAUW9
GukR0qAt66pv00UnURaCePCw0vgc6oA5zk1UI303BxSWi9jA3xW3OKzmmJyhfn7DciuLaA8QiA/L
nISIyBSXamSmVRz6aeZoHtZnaZPXg2ymeQWSjJXDn1c7IO+tu94hhWkfC6QvJu8jgqME8Em8Px+o
BpfvKHO4rkzdWTU97RBgwTIuzm2RGrw6Hd1IOK1AS1wPguILnPogko4x2RltipuWPHccx7WPNfDT
wuFfAO+Xl4tqvhm8jIZY/kQapiAd5Q0LOa+MFakkjYVgr+/v0m7AF7aEBbUatuiGK17I8Ydb4Vkn
GfQxQlEXPFIJIvd5M9DU2euhpTO3aKvKSPMSD/KMFNjLsGrI3mK62DCgoCt++dLFRjGmPgNjxrp5
qdTLocfw7DAcaNNGQSqI5IUIUpc9WqAld0XCiCKVZPNIjwI6VEWLRIfYjk+K9IOZP/CJ7cL1VVgm
K/SQbI8kTlw/SmHVD8s3PoV6ISc712deFb1RX1C6AV/yOHTSxqXGhP5a6K4884wTrneDvZt7l2SE
yQyv8tOIBU858uKiB/M/+4Iv+KBNPPKLMd8BZvnAKPp4OCrzmGCqZuwoQszBYlNuhsyP/GdQuTyL
YsC4FsDlUY8TILG3jy1zOZinUzdEn4K3tyLoQr3jSLJCGRTRyJqQG1/vgI3HYHBcBfKt8Zg3vFA+
eeLr9DBiTQWMDGTrjJXvq3FVGy3NKc73WXz8l8f08+dx82IVCjn+GVqTiJjbh1EJr0r1JpQpWtiT
0eZIJwDyU+qPh+mm/DM0WKB0K/Ni/8ngRp0kbfKeBry7g5PHIDRYAN4jt0dw0/z/+u26FH8nmoWd
rv2nOUJ9bunra25qwwBP5HoJBpCHAyciiQbvugF+40wAWhdowS6PXi4xjTahEe5y9m0iUkZd39FF
5rXyOpDH9it0exnm15wL8Th1n4ABcw6bzpa5LNGS3aHHqdhSo4z1FR/M8tUS13mYhAN/kfSRbYD3
nyuhEWXyV26281VS0ER7ccPGfwG6uZBtkKw/j6SVcwl00P2iVKok1lMYx29wINaJFl4eUzrpFWx8
GnnpptaAu6YBNfT7ZaD8O3fLmuQbnxWYWflq74xJyTHpGZZsqjNncPB6eqFmrU2T5CAtFteEuxTe
uFoC0sc78T5ol8y7FK4x4TUHvfvlfRzlIqcraGJZEDoh2/oQqN4FgZOhXySg4bw0zrMu2WbRUDjJ
558ZVKF3z0CIZjKMw2daZ5YFEuN5SiaNADfPP1DGTTjTUALmkJaV0YWmqxXwfU+/O3vRrv+PiaOP
VR2LXn4REfsCJW1AR0LsgnaHdJyAf47E21tux9LtEO7hgiSTn+j2IWgQYIWs6fgXNrq/54Icen1L
f6F/EuHzMZBza4JsYPGklPQk8rlHz3Y6RF6YZIMo6CXzm6QyrogNxil6EXdUbFMPqcfpPnj1OLf5
isRypqoRY3a5t3s4gtbAFGtDs7ZheUQKgEusoJYhvE2f82HOx1B7BSHYzf1DNwQ8MnBvgfEQ5mR/
C8Sh1TGjuBR1tK1Bylq9tcKaPSvSrjsGiAJdeWLAnRWPHqivO/SNAj/fR3IxGkychds2JDhUXeGm
TPDenwZXbLEOZuXq2cE88SDOgYfF6mlQsvL49uLbV5Swl2cG+Gua63u+GaeXxLU5bbVmRepn7lTl
AkHOM4nedeQOP70jYIRg+gQ1OOBk3exe3PGf0z6H2lHMl3rDWlvEMk0ZzGPNjWrKI44x2ig+yRlO
EvqFp0nx3dlI2k++BFmryoVO5L0A+ebMC5wATFTab/vDwsXihf2LyUlPkkLziC2VjduH8hJSD7wf
mVjXHw12d6RLfO+/iOba84bnRSJK4k32LvyB+RxIPtOkfIg2F9CQqr19dsMzEXKUa8JZn3HiokgB
oRC/hx6XUP4ztICFaDVmQy0hUpTXqnW4eEf2zhiwaWU5Bkk56e8FzTNXZFAZC+ETllZWBrefvLVf
IwDO64e3I0lpo1C76FdFpJIA4ZkFEWZNALF3GGTBM7pD0F1hpfxjQ3U6iR3eFtErmEcCocsFtOJC
6G/VEBfkC8dsnbcXAkpcAkZZMitUkE0BjDXHBNJoZe5t6ql562U3kDCj+1Iftlpf4lLIlDa1MwFA
GhNUVz1DJGnXfCyORogTB2L8py/EMi8x6ycWs11BczCoa8S7FMtWCTnXe/mi4xwOMj5IWXQOw4AG
xzlIVtqCFMu1wbgMAQI5ElwbDn6vSliT82DgY//8VopdW9FP75yQJsYdj+gOwSxnT/Vq/RN8AqqB
JZBOwJriszxAFsDjmlYpqpkUOxO3gkihfhE8Q7kXM6mEgGrOfkDKSZW836NP6+t0AsxdFdwOBPBK
H+gnld3fnyy9BiDgS6lEuSDIy8nlvtI7si/PhIReLSCo8lI2OjB+hceMnJHwAfjfybrxDLSVEjYP
QNEoHBs56SJimYoFxtkezzLRDyeLTX1HcE1Bd4OgrPxTUeGwLqL6MW52Q9C23r130a1Nl2uQdrij
ItJ8L3OMS2OEOf1D67CjL+TK/QtO4RCrT7xBvg1l7/e9op6b1f3++KHAlbHh3s05N8MC8HhoGix1
CXdvIHYPUwz69ZOVoB0CXMAlzMPzY9A3LJZZCKcy0LD/Eu9N87Yf8Knqsd9VqrGG+5Don84Xst3r
hu4tUTlOe7jeVBjMhXsUIPlTIw3duOqf8zhbLuXFnYpGCA7SigEtFm7dYdV+GBbd8oZVzEYT+75t
oa1xhzTzz2Xy38fGpBPPReewJxjZ03LFg5IvITpJgSSrL447FIXxDd7cGnTKCA98+Td1KxV3NyBd
5cCs/IPXl/AJeVG5KbHH8ETLzFAuBcm9oTB8zh27m3MgrP1Rh2FTHmED02oRo3bG3BvehnPQCKz1
NhY16KNvwWLjUpJDeHurgUeiAHqRAa6O1pFEjmSJ2JFB1QT/TdcYo8RS9Xq+HA4edhkNISuGAK+6
5psJExV4m4TpWmWrFUzi5D0jKluuUeBD913oR7ER1n3PuYpjmt8vJFrTUD48pxMlbaeU1VrXqwQT
PuJm4ZJz5+ub9krzEtcalrSaHL1Twg+dzzIpBgNQm18AbttJYJLjCOA4hcJoiWvDGzk8JnBpkDNu
RICZMs2K7Y+uavPWkTQP+RPmAKIO8dcaajpNnnwlEJoZb7gpOsXR9Mzveh3a1FUyQ+2QCbb0+GR9
Lsi7TMFmhssFYXSuwYDwCcCTKlAR35LlWGfw5e3cZyQ2XgH8jTXYMGhxq10gpT2XLRlSkodxBWfC
B9/hovEK7M5X91CK4SaHYf7RTDRd14piqYPXNJ5TDqgZYkZooi0zZD8+PUPAIwxH3+9Bc14+irOE
VfbTl768ZaO0Z4dnR6MORBbVn97b4WaQgEzB3dJN5fkW5wlaoYLuOEc32CR0AAufQyko4AaAIiFr
TdW0HWQKllpsKDd5rMpANTtOy6534UEOK+JPRKuX11fzd/K7OMz2KD/oSc363YOppb+jcxd0pXgW
W/ZTdGQZ0t/Gr03BC/+iji51ZuoXxZ65qT/rBn+VVBRp+8WZb4KiuQ8BkxI+YnCGiADQ7ypr7iKs
JVkxv5jCNPaIrqr7CV8q3lff+mF9ZzLeaYvLg7ihYbuyEVzVhgY4LWsK0mAGqrTzC+H/A7OLZyLS
7Jw6kbZWMjxbt0nE1YL+CdvQ37pfz9j1xJocuvdQi/MAdpD/JhVvppqIy1Kn9BtbbQvMFXnds5l2
IDSuY1A3hzUjY0J62DJy+yJUDGp17PvG0dXIZw1fwhCmkw6LzjTS6ac67iIko/qJm6s2KB6Q7Qmd
M9xF7gUMvZ8CMU0GYON1UOxPagH234v03JjdFEPgfIboPBYT5JuHfRmjNRCElRGAgsoOWaW+nxHM
kMNPItYVrMhktlcZhA9HwxW6lQvMlhuEzZesMObjqhXkN4/O18Y/X229bOdpIEG4N0GdSkTEXfjZ
6EzE2c8Oc339Ljm+OLSs9c/E+wAXv/pj3ZqZ67S3sYZzHjQNR/C89DMnWgNd9G3OLVwoLo386L6w
s75lSaubi2SNYJe6kpzoSJDrBv0swlB8f8sfZ8i0w5kcnIt3+rhduFhrub5cH1Ype268jzk7Yc4k
Xsmp4pMiHjKXl1ofXnhVSDbjlEus7d7nuI4XvOxrsB7DIFwuRbbGmNPTLIb8Z5WLTio7lAxm1YVJ
XQnQmrESovpjlUyCl7Makl8OBsrL/CGrrH58/9EBGwI/etS+2UuFrtfM3JP1MqC0nV5qLafJRG/N
WyhYJiMwWOww6aKpUNcgDDuOzEA9ERYAY2KeLzgCWtFHzX4vL2LZUfwkwjtPOqpk+4RZfDFnIqp1
Cn9yW8cnpg4ypdPxs53q1TLOf+oPQeHygsizXGRp9NUxgZ4QVIAsYYF3LySb6xg0Eltvs/LIvyat
IwWCnEzzrlvbYo13nnIvKAyeVxeFym2fUrDJp6DhTh/M+0mJNxf8whCiGqxoee0ZErob2WX1Nvwe
xqaYhEF+ViBOxlHoeSP5T+eRXCXtO86m76Hql7xGAQPvSze9bv+Ukq1ChWpPP+rHi9gj9UlP+YUK
by811/uL95YBUV9PycMlarg59hA3hTzgqlv8NmJR4Eo5xdp7872ZuVB4n4k+J3SMfxvt32sZjcuo
QP71Ra/CsKwZr82l9+yAsLtiGCS+WB9JZjL2+U2JQqFNiPf3P1AaT44P0OIKzxkEOcDq7YURtPvC
6Kgc7EmQTbQ/Hq08J+3scFBQ+7aOXQCYnoQtZki5+weIJsHeQnjNic/XVjs0/eANdBx72CurBuiP
0aQJVwFbItaHnccQr7ab2YJfC3NUA+L6xS9LR+CiH0klptLEdDpFT4OiVDjAZQSGAHNof52QnHtv
266zQKMqWKzQCp3Dt0lWjGOws0d8AViw7TyKCDyrV7fX8ZtT0Wf+lWusS5FMZWv16vI74MmiMi26
m2015983YWPT7+oAyZuLodYT4LyRBqP80lm8uiJhc9O9Gt4Yf0DBzPgwAE1LmIL2+blvgPBFlyNj
cfH5S7dwOenglvsal2bFgoEPD1XFi7KQOzZq8Od7Vc6usBNxPFskfiO+fRsYQPg9iHjleCW9yr7b
CUGDWeOjJ1QiZGsqMYTpi8aFAsI8YXrCwdCsCQC3ImlSE11z7deQA5KDQPFO4Pt5jfKSTG4nCkyB
XrqAWIstHGf+ftvyCcjuRBCaydyXzEnwVZVF/28bhacaUrtfuViTHNPXnF+2/zwNLKXjUFJiaSNH
cZN8y7aEQIH4zA60eKK779R3D/PGqJT8sjYfeDFpm+fZv3ndwOoBeNkWIjWb0gE9CcIvxVsY0FaC
GkuOyvD1+Hmpv5sg2EemmZ5H7WJ8dwqbSiauAXbWQRW/L4QriWe3iMUyikaRewvErU9mA9yV73eU
3rMXCbYv73K3AMJaQhIVHb/11YaKvcBjlLRj5phyPUhqMEkqrWvr5j7vHP7vhvrqNeg2H5nifHZe
x53hCSfImqyQyVSb+IbrsoTwXrpodc7mjwLdaXY/Ii/lY3y27yP7Akhf0JJib4Zl1/MiC4dg/guc
sx0pgQuiz8b76I5mIU7h+fu5loSBaym9/iaYeovqxerOxAFpLzGvnioy/uzBCxnFGbkHY/Emyn2K
bBAf7Xz1d9RpsQUvjyb8YFDkrVs72i12A0UZPZNnig/usd7HdMe3CwUUCqGSYdK6M9B820CI4qf3
b0PL3phJOdMt2twKI224QB/xeb9Xhpc46aoLb9IIhRxOH4mhgaZedyXkFjYlie2JBSuIOqKO/KrF
ixLlTOcmlsWxsGoBBNJqWDVt6Ko4AK/L8AchcRWXnA9a38MJLjl6kaD8jSEl12kd50NeDfIfFA4M
3vQKRKjcc3fZ1ms9vAehLCU3TUHGsc0A45s6oPeUngxL4UhahepWM61YYchquk6ngh08NeAiVRqX
jY1Af9TZ1lsGf4vkumJo/rS/kcu7H2aDKSrREpApwx/L2Dp/aU+ptmXEV+fbot3eUscjIopsenAZ
uUZVoYKS2gOzlJuLyKO+OgfES7PA+JFDIsK4D2O0OqK5mVCrMLTczieNG/5npF+mbxvgENEwxmY2
6wFbeRi9vEiJIdy+IZk5Yzku291dv0sjC+nYf0u/uo/PQgq752swF1DTsuHNnVCRlYC87oKEFa8v
sKetSWujqHIua1EbsILYk3R0V1Oex3TFQ8FJe83Urc7+rffwDbO5N24z87/QjisptHfl0t4+Qw22
Qxn9CE9DSHRdExBq/2qc4dFHy2UNfBoXLkQDepD8/277iFz4Z/y0cQcKyBRTdhU7Ns+CBr5GQTUa
YFhbiBX7qu7iCwddc6mDJ1rFCD4+yvffEU+8dWpfEHLnKlftCJhgXb5z/U/OVOPw6NWlpqejZf7r
zzAd3CXOObEI6unwZIuOnxpi4sTfUmZdaW8A0+DWlSquvexUOWasfqptMHyzw9lAyqUITU88Xsyr
SGwPnsh5CIArfLBRaNSSZ7LXYKMfjxanckCcPIaYW/v4GlBJh4hS0ODFNkGtOVBwdkzptES/wJui
XJS1BCEA/aVfrhCdpI37KbknPqJZYCiTF8XdqDKs7V+s9VhMzlppr5iAVZHN/3c288UGTVUKVB2H
mVrScHPUOj/PvhcUWYPh8XKPZ/BC/B8h7PiEn4R//Zih4AhQ35tgn+B1jW9udEsZ2+VVARdx8j0Q
F2Kp8s3OIdQIrpgIY9g5QjIRWS60Xja76jrOOqIdumqoRlbmA1bvNGp7LnWP8fAeKH17oXQBCqeW
xdnqcywj7SxHT2+G+Lx+64Bufc6cEkTJpIA66lsTBJrk3JMdt1qeDA6rd8DcvssPq20jsPYFHqNe
FGz6u63Zsc45Qwp6f1UQfjaGOMTvSIXBoD7KnMTkA054MIIykH4E105yDQ/QZVXSccs35LOpcLW9
XLujvohwRrwXWdZUg9PjV1YwHEl+043DFTW7rdD/3QXU9OkkV0XtTcruVTk1km85TDAt/jgOVHlC
TwtSgtR3H7D0nvWtWKdAYT4i302dTja87fDo+e1guIrM5by/wQbkQezhMSaAjkquLNmZPSdxYWI2
FFkF8Tr+hCAqlTxqMtFT2dyXd9I4InZo5/U7Gx5LcEO+eTEMJC5g/Z0+Xtp7oSeHCVcvLHpOR5+R
b867xqCjnZbKUbjNJaa6+kJ1K1bqljz/TH447fY6p0/Uc6A+NwOGkq7/9bGREOCFGQLExhhcv4vg
T9bqLea5Za1d4rCnTDV5CttI9qEBFhGxBWguwWdfYJmoHWoi9/FB0deIIMjii0ny0Tr1lHLl1/No
RPZB2iF3wK+Lk5rub7EKvfgMmQiiWvj3WpA3U1j+73QqKqIi8DlMB8t/HkMIWlpjrKFvZIR8oviJ
64pmu+b2DaSAiXGLPh0IaJ1/vLJXyZ6GKNI5V/j0GO7axgoNdNdMdoLSEEC3wrS5cKKRnzIGXIYm
DGdyjzYFmG3QH95qMVmmUkqg0X4Jqq0q4GNMIJBZk/vwAjoU1XpEV8rgWzUlq5DPETpPTy35TJwO
Ekfo+66p2RGk/Q8rNm4ziCs741xA+eQ0jBovg/G+dzVvUrFDtRD+uxNXjS9gFHm5i0BrSIqiQ7yF
AEJOKgRQYfKZy4rqApNMNHSkZ71hIw8VwQwKwQ4ODdjMNSFRgYw4B1CSNHL0UrJWYRJ72JheUODk
uf0w9A1RHS7xN25ip+b8B3I265eKIqmPcFQxtfdifl6oaaNUGm21dxivdLTXkY16/WnQXeCP0Hf2
jS8mp6pllGtzgyKBFzHIWWe5HI6CCEtd2cMX2mO2tLR1bZ7nHPhz784Q9rCeQzg+GG0ye6SUNl62
KNqX+qgNl1UsIFJIOfkfjN7PDLEJ9TKT9Itgk6vjMEuHp4WMOQOpZTPBwHKW/FxzmquTdckorkiV
0bB6Qf9Zp8ddwPb5GXXiz4BCnyXS+1TP80pWr39kV4xDRok4kzC1Ag2i9K16juvfWTEgmBD7+Ahd
pDEvqJoypQI+dIyYUolfFGFTik86NW760lHvEl9n2VnrMPGBG4NdBptLqLTOIGza9jUd12DUI22S
Ayx9dF48MdlXNR8r4Xe/Ba1tUt4rIyOSAVVEfTeR9Cuy+y1U2NGqPWX+5XfHAEh/m9IuGr+ldhCp
q2A3+APc4ot8xoyCPc7gSXBbAXUyO3tKWJ0D1w4ZaEeW/5TKveDwjNtkqDvZc5nK+fAqvlgLjgDq
3scxTP4bhq8DZZccCGWamqqcFTgTAWN48H6U9/k9weixSPXF0dBLHSQcoKR/WngkWVxJOficOWfr
euDwKSOFAwWT+EUL6UAW+FDL9vx9HCZljeJ7630LdLqKIV/vgDu9dkBZYgttj24N1Pq3l0wQxYAu
ZkJk70ApkmsSBEcq94cflGrfu/jI6dSX76c436+2cpo9RG01SMzS8PZzQrsagtrdJ/fYRZXkDkUo
0V0bG0KYrvdMpaVnZfs8IhJlpBRIIR84WvA5rvzNLbynPGoZR1exOkBWE3kSjqcJKhBHO+X30gtu
r+orcYyEaQjm3lSBQt2ucpyLYHBcxcZPYN51Pw6e+/elmEOfGTj3vh8G2+S9LfNPAIhrLrJFTR+r
x9TCQ4fmqp2Ye44lfV772mJA4GZjKZiWNjfmOAYYZWkH6jSRzc8tjyDqpXDfFczGbPvw89/LuEpH
KER5/Hs+blpftQ+MhSR/J1VSiqmBCIHoelGX9KnCtZMzG4IGlO9JSHhxD0KF9UFEdHI2M1l881/e
xM0dMhpj3K65HwtN0JK9pnQit0EhPTbK5kLQJsAymY0lQTjazRfiglnqMi9dA4V/yKky0Z07EErH
ZpVdpZPJF1x4G+0pRiU+y5Q5W0njHdA2O7UVfHDa6EUvuTJLJVzgXXnxR/hqHFj547p2svARpsAt
dQe4Hw5I+JbEsiqufL+TQHG3tNJm3rhufcX0pS7Xwtp0tCFP6rVYHyVuJlWcqQjZpNCv+9U8iLQN
V2kXDb2KOaQ2XQzlwi9JsGoNKkWI+0sU5sCGAQ1pWnjVjbjNhkrTnseQQed73N/wVW0+bemGZ8+h
L0hfMiBs8b13I9peFJIDQF9CBo7+EDL3uN9jGZGj8Pe3kkUS167HWVo33jNzM3ksJg6TIjfG8ILn
NnYWnm0XgI1gbtQGGdP1bPivZfe9C+XrFetArGp7MUx1LkeBm7lOFlE1l6dB2geY3Dqo7b5puz4j
aTglhPRXqMDflIzMo+vkm5t6srHQ32Z1MqC+AjgsCUg1vldx1PRw3GQKux6sQ86TmPAMLQjT9d2Q
CzejgJa2Q77O61AJ9sNcrKUMkMD8GYbZkPkuRB5BNdglHJTqx3wplXC7DofCU6bBtImXCIEPL8QU
4opBsNfN/B18WGUt2aXUdsHwuYOIFaidebe83KOl++LHspe2sgPn8Hvb7BLcQkTVvjYGuPOiVj8M
Sxko/KySY7/q4fTwfJfacheWU563npQcPy9M0AhYX2nb248zZxjr/iG3MPGd9j6QnkwwcOCtFWlp
GWw0iNNWD8UzHV4bon64mfWywVNWmvcwThRnEQoc48U1c62CpGHow/SfdIqVmgr+AoXAR7t+6Sfr
hyg04I233IkdAhUFG5VqgctPHylSwZa7ipVucKbtyfEVlLmKJAV5Iyq21mO5tZkgkGEI51Obde/+
9KOyYEC5QDpidBEao+/ioAIajhguF/hHOwcsXnO3oSJX0FQ9QnCXclm6/LQv4FiYQ21X1ts6HXRK
mcU73CYi2imBX6c7i2c9BFAl6IdyK7FeqKK0EwNqXK3NbkXowTwJpms02LxofWYV4m7geB1wWd5e
TjwLABXZFfF7DPR0wjMZyED++HSC/OIiRgDvEDYABF4EbVTN2ktzL7KMe1VRLF9/PsqzM9uQhSlh
//YXjtgaUBDBZ8+lESGgKUpJqW6GFZcuC1On1m8UrCNufSKo/LCcTUYvy04etGdGk7LBdq70PLCn
EVSbn8jpxLYr/0piI5BNCL8nAdfPQd+o0C+UcUQNiN/pAr5SSr1BluQPZGgiEX58QryfwuUQOrD2
tZuVnmWIs8kd78/+Yfs+9AW1lPcafGtOon+H0zw7yAJfGwD2+JdSPPqYhtDQLrGcSzJNe65QW1av
WJM6Ck6ambWzFtE2bJMZT/rKjbiI6nd8NEFRwGGFAunuDiykXLLoQkVLrr4IDJSnsalEezXyCDDl
m0pYrVL6P2JLLjTZon4/fZ4mE+sRB9hZdaxj9LN2cxe560I9kSMHXhJT4S6i8C+sArkwWoBWe8Th
G2JgE+9qI+g+vAlcV/WmsTg44TflbD8+ljDSSD1Is3VWVRGDfjWCo5zG4bihceKfF3VlVhFjAmCE
UyE1oJY7pF46o3+AXLzuG+/uoNUaHsc5vw+SL4RbCFjy+GzAOkangtyE3ekZyjALh+bT70JCP2JZ
0NgFkwm45U1Z9op0n0XezN4RESt7CfskbEj14jCl0uIh4C8EXlGa/M9cHqV5hev65cKtRiiaQpGw
jBKFtIlfRORLaIOJV6/TPEhpI3gd6DhCUDW/2MsOzzpN7JCUVQzy5fsTSXQwTB/NXpRq9ejH+QrZ
DyiTEP2nOZvezwP6lDM/rzTYhMAKFSbNdl+FsveRe42coDuWCOlp9dFkCEJVKPaAXYEEnkwD8nAu
cnuzCc/5hlbjOG4MZl+2Lbg7gJ9eZ7Kl44E+Baa8lTfZdMb8bUclt7AyQXtze/7ARcf6mMzG0V3m
ElAUbdbSDLWKPCqMIJ0PSVZOuGgVuQc5M5MtZGATZjT/4+jtZHAzlXASryz1HI/XTJTr/y8yg8fv
4ko2xiCqgquZqsqS9ji9RbN/hgRlk6+ECeAkltlJK0UvhWWyIWDumXa5/El8bgqFxFpydl24frml
dQd+VbdC8H41520j/RL4uEzeVu4IrxXwd+Mx6AXtK4cVnTNPLd1Z5kW+mCnuloH+N5n5RmI+W8XG
2RWcLeMZh24vJZqt0VaCvzHoMJ/yWdpnu8UeQXiR/9t79Z9ubolXOYWbyTvKtcf0W+1u5m8edA50
JbXdQrK+SLSgIn5IyUuEcszKr7nWPW9FzgQ01GQ132O9vYK+Kl1xUVopQ2LSAVeWaLMHxRtWmVxZ
V139dPxYjt7XQ/dxvcyB0lIGYbpuAAlbitSycYZVscbB6W3ZAeCZ9q0Motnj7Mnj1SH6kYQBCC4T
NUlJVkT3VDEn3+OFRiTTuBVxmVHNoAh586iBv3piuUP3UTj39AfEEzR7HDy/TPSswn1rULc7DJAM
a907fCqWgWzpj0kbvJ5tEZ1rBTQ+1xxgEm/8n9DkpDZu5oEq5HExlnBiN0TDLWc4GnSgowTTHVCM
qi7Dw+sntMezZZpxaqQR9XjhIahdcT1655PJnBUcJNYzSWxCcj+JEtAjIjXJXhUSW8LWaAhjWyLA
gEA5oY5J1Ql1HsP9kAZ1Kauz+4xa9eYlo0apbnqbL7Qb/NfjQCpmxAJSpwLZyPzFClxUGfb3Okni
Lr8AWD3XOhZN7NMu5D2n+SAIayIx1LwoTJq4UNFoX0SeZOkD0CB2HexH1eMH4Hjp4Tvfdl7Vd0Vw
lAEt5cZ4IJktblYf82mwKLnVV7N7ABUXRDJpWMPU5Le7kgllMB/pt/73AS7EjkIV/mY2LHGcJ9Ac
wBqMBrOWJCzzKhedZIdRm77lJcGebtxA8ylilJsHmubyfpK86F5A/gs0/Ix6/gmFIdLTes62Btwr
veG4dzWvnuvFZqg2XaqVP2XmKpZYM7p35zfhHgWOlCQIBQQU80/PSuZFp9nltsrawG8tPoGBfhHf
M9w/vyCbppQNX3w5Djm7vLKXNStPV542xYvUa4SyfQML9c7U49/DoZ6F0je5LRTJ1cC8820BJ+uW
FGWo9+A3YsQg8ui4J7k7SQ2CXtm+GeFXDM1ccTTQ8NYhlTdbPeLRM5dUcR9wfciTe70/t0vxnRFY
YAkb9inkA0nfYy++pKyKiO/nZ31b3dljOcAXZqQdHIcGZONvfGLTqvIbtx3wobgx6uRP8yIePrAt
eDndM+C1VXCyM4v57g==
`protect end_protected

