

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZqI7Lq/aGyAcoaejBEIk07VX9jYIkvdeTPQu9dSbDEADopcPNa+0k8THWemULZmXocovtHBV2sQ+
UG9Mr3L0hg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R4vPs+jPUBq40hDi8U6b9avbUk2Eb50U4A+mDDli/Y0olyqpMjS2bHK8VDjTVAFuQ+H3qih0cQYm
+ik1m47VLNMfNDfRLbftE2okRK8Kx81MRcEafr+7z29VxyL2KSwmOKbcDCEkIT1VX5y+96x7q9/g
O5zX1cVuj6hrFncQjBI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RHGRLed4zRtfx3HaMZFysMR3Ua1JohlSUQn/uIq0QNaCK2P96ztDgqQoqe6ZQ11betfsHTRFzq/1
66ClFz6QxXME/fh2KrrXSgUZxYxwfstEZlyOThrSfu+qzCsdk0R654q7wyvVT8+Lni3RuXc5nFXx
raCVZl6qLm50r3EadUq562wDBW7iVkrMp3OgccKyJyw39sT1Jc+0IkzHuHqjKA44tfGTOOSTHNUj
YgsyeZCJS72pabS90ZfprHyjsELB7Bxw/M9/XLEV7l1LP+SCDJFvOP5dNLZDBmwYIJ5OoU7247Tk
wYu3m6ZFZNnTwWGI9SAZJyiXILRa8hVZPL9TSA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OU7rNiePgxinwm/ruLBNeniAmTTLdwPhOZ1i35IGtDWXtaPoMnsPLRF6vnJo1xeYUES1MIlBqaG4
FUeyfrnBl3ofk5rfTbxL16dBcEtA8Z/duJARcLCIBD/J+xf2VlSqIo8dG9Ww8/L9pBTHpNAObSOU
o17xArTTrLfHWXZRGfRwuRpGlTLTYOMvS1AGhQcPbXjHrlijOoz3XigDVsnyGbHfkSgOlGBCnyDS
TPebi8IC8YIl88ieW+lqTL6jl+3DZ55iTfCJKbFt/HrE1Uou1l+60xI/9h9XhrNzE5ANic5eFmyC
tdncsHEBtx+UfZhyFrHV8z72yZoLCX2rOJ+IJA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GUoHfgebfwQKNkw122kR1rRfB4ZFf7/0xjFIvV3auOQ9RcZO2jgecvvtUAn3nocoMNPW1jFFZW0u
xgkVDSrwVJrMR/obpu7gqo1n1FD2E5BpOJV2Gwso9aZGhgTdfd0mINfCxPi4lxUYuTw1vd+iNkBH
peC7j2xzDHSu6o2S58c=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lW3oa+bS7VSdBch0q4Lk4kIel2MxeXNlqo+JkBKYCThE5vtBv3Mob32tRj6s2h8BAos9XGsKRu0r
zWpu3cgAnv8lYIL4/UPBP9T+caGqWHHoGULrLn4zuybUvPzfGPj+ANXGfPXBomTO48UgPFWBnBA2
3vlOjCiOyKLMQAUrg8RqpfdYfcnwHxk8ebrE+lZJf6NCQtrqGu/EnH7PYFH/8MSQa6yey02fLQ2J
HenzdGNam7fu3z20gETHgePuewowRrJu5bEZOzlor2RrSnb0hcSbcO4/KSA9EcbmjzBMjE5uRYAM
1y+0t4rNGr+0XAjpp8m6B8lGF+m1jIGYMJ55eQ==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AYjoOGO5c2rCxRUY5RbgjfKwpMKJQrCDGPu9wzqv2ZhoT9Trod7xJlCnzNNU4kNJPTgmDf05Bkoo
EvR1hgWeTmTgCGdy7Qci0Z0L3pdxnOg9i69qsJO1qAW46sOYPeZHpvATo3irsreTIyOEcblYRdLh
Raj2T02eEhljrx1UdWXHwIq6kJGwbPaiMRXRJewJ75w53lF3nNUwTYgttUbm/hKuK4MTBvyDWlHF
UReBw5kEbERTaRF91+HNJUeoBgfLIgVhtPzX3Yzqy4fl1PxZ0BzAGNRQWfLI4TBSyl64znmxdzaS
+wcpSJ3OHZL4sBSIwGqpZ8UuNr53DWWwkd5lqw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F93W5rP9wRsskpVAtvm9VhlFJY5TOuivcFKT2bVYmeqxn925TMU0N0nDRJZmC+O7NbtC0kbL9Hfv
iPaQAjkvtWKCEafU216A83pjNwYVINq3GbStXAtCrvf3KbYJMQPnr6FzKWLa0RlmEqf2z1LRIJMY
cR3LKzziLGgP+oQLz6W3siXeoyqxsbDm+dasSbu2YxzGAvkTos4kX2slGrQzxYSQogS6j/MzVgIk
Vhsm3BYDbtVT5TsiHGfRfi137tS2Q9o11KN44GT+JYigwORe+GyKi5xjI6kGPl1N1DK12TlRGsgC
Wq2YWMn2ABYXE2F8mkwPOJqSaaAR0S5MMCjkaQ==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EO2KlFB8vWgjeXvua8SEZL2APl0WfdPtqoF/0VTjBDZhkKh8T7GBS9tSSrCin7kHRBUGF6hOUPK2
V0JQtp4yW7c3oVbMN2ePIV7UdtkAszA2lMqOqeKJbWn0TfxRWL5adG+jGlhhYEbaT6tkCGPbbtbk
y5Kew5kT3RyGP8Rb0tim3cGvqi2BdBxqdc5Sb+Vyj0havZUyZo1AsjuLnNukDIYIrPCtqOY22MTp
VlNOr/u23OIMx+xx7Z4aOvZacPCxfg662ljyHetf5a0wu31WI6zf/69lkXq1iWJtHgEJn2iDpIWs
bSWDEtGgKAFHGKVAoc0vIGP3aPG6DIsqRyQ90Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967968)
`protect data_block
VpVJ8QYMIqiYZKvsHUHVSlwOpQe8mSP2Q4HFrgvYIsAw5HUkI5bHK3ZU3V+uaCVmPiEg7MkukIYK
ua+ZnYQWKmhGRjqQu4PKE+MtsiIIckRWGY3VG1tJf3ps3XXGtq7GHDqZp8lQMa3i1afghxTreuyB
nc1oFop4f9BQHiOPNXfKcq3DbeDx67/Uf4QRz2hHwIfRpPmMmeBBY1Tl9FzZ8FYMf9h+4h1PtWNZ
fvQLmFF7olDfYovGCirrEW80vlbnkXuH9xK6IPJUT9tRrcAzgr2TFxIazvBHPssbuCO6N4FLtjDm
r4+C8kdTW8iRJVUqJ+JeXb7+KuwxBXS7/YfHJsni1xBc3drF+eejGUYYo8dMmiw00b8r/3r3iiut
us8y8SOcJFdySqV/tmIcm6cQ0AFQA4EDUvr5GEyngun8T3A1OmGXKMFFeDmiiryQGMKBBglfPIyS
oH2Cn2cX/8zx3LpBmRSnEDh0ViH9RC7/2Fr2byD6Ea7cjXCZobl1XovDyA3dcO1wBV5TkpDU6Ba2
HEz1Fk/TFtrHsqhRHO87C5cZQhjaHQCWgrTl9HB7lQfoz7ZaVnW3GbQ3GWEy1SMsyTsS3ztLNNQa
TsVJFBCPG7XWfy3e2RDqrecwULQVK68Ieufnkn9F0CVnssmcRafVe868qqAeS0uJwB64mSNAv40i
1xSN9K/wXDjFXxwKd99alm4Z37cUFUdNNn3S0+JG6Oto43RxcAqsFEojJbTRTYPoiSJHp8VsCGIa
PviQMRrkEIlJsuJjbVkPBdfVazz0wE8jhMcMEX9291J+u5Kc5M+CxCuzJZpgx9RGUlyo9F+s6YYJ
CjT8KtBnJHt8OPotjnmCioRoBdX4uhHb3NYkfhZb9tvVhBy5OtpKmtgr1AtcdWGgUcnfFj/81gXA
zh3qQGd0cO0yKbIXFoVe5Rr4DcYbq76GaU7AT0uDpW4PpxoOZy1yVNgIuLp/ovStiDGal7X4KW6G
X7S09N/2TKOBj+sV0Q9FBi5L8KK055fVkEm8zJEvButppZLykHaQtndnTR6hWurl5MVVfmAgxE00
HiepR1Gr1GI/Q4u85BKl1+NIYW77bQlYxw/cxeicUU3cSKcGs/Nt1QzVnpHaY1AAKOoVBSK5QpUL
ujz36Nqbm9lMlA304A+RnaF1u8Ta4WbQubDLtStlAuVBpjh1TKw+rB0pZRefA/gSL2Vcn1DcExZ7
mDYTNCQR/xAghoVpuO7JQGVx0EcaXLqJHi+lnNU0nc8czhGuHUsYbqXvCvhte9ZY5KYVbiIzRVl/
PXGr6LDEwqfQH0+BRFczLi7phncBjlhAKWgUwUExTB0Wp2aF7BQLLuvoZX97LxFkNPkNodqWdYDb
VGva/LKuDQDa3vIN7nrziWP6swa6TYx+bbwC8Kf2+uYsy4kPChQ8fl22PhqNd+Carwv4Z6XZGQjP
vC/tgx3SoriyQScw9MjZ80FpSwRYSkuey15eWoBRBtoOJKv7CIcz+NSLEoaLZmMfODjA39c8PRMR
LOmbFnHzDzZKyrRq2Wy+Xr079XnrrLKLbDiZYRJnDVre+fXDUVxPrAhdxaOa6cCT/tdAjmMW2yKT
eCP1kgeNk69UOKFprWYO7xEpXgxZIwPYDUS59OnRGT6cWzwU2hpihYuHtigEBAnj5LXzhLZpY/cH
Hc9MZfM7xiIrmdSDAIRX8df4v4HVf5yiiLilwtPUInrYkHvejVow3oliqxMh9V63+NEGkark6gRm
NgWoYIXPQcZNJF4YPA46FeOVaGM8aqNRICvuJvgHXIumsaG+tg7BFzAH/8KMwzLi3LNY5cgIsDvT
4qy5IGlik2Cu6JiBdY4sAzqrGDeYSfhkI40lPdEmEmnx2CGVjRLMgTYL7nXw7QREBQlxHS85YJNX
2ph2vYy0DtwAQx20uyzf3PNKa7HZNSzc7s4bbJK6eA4hkirUTHbTODE34OqAUPrkBLo+qHCiElEF
RZFXXKJJ7fmve2zvCksQijtfm1zDX0aA3cXhDvLi0v9UGZVOuarE4f72TOzyYRzq7o+43+i9yIc3
Ohl6dMAxx56MLYFzhOLtOiekNTDhGLP/Px7jizxuiuQAN9p4EyEQDbTC4LdI9PXKaVkN7DLxEikX
lGgMFwxDbeZ2rEX34V635O4V8Oqz3HgRIIwrlky8NKxs4cYYNgyxYrNrnmUzOXm06iYQInsEWDyB
UhaapiQGt5B2a68S5AwF6BVzkxSEBvsel6Y4lc+bOLYF26tQ/0m+MshUYH9zmd8BpNAneDxRxTtq
BwwokA5VUrn9DKRdfrnik6MhBbJ+oAikM7vFA7z2FOizyRbR3LVttCT84mMZ9bRUtdQ1Q+98CE1+
3I/Hdb74nNF9yI78PdFDGAV1P8qQUez7B+1cK7Ps/EHBnKiq3Fj2vnH3d4CjhZSZ8XeNBRUt2ngJ
vEZZupdvPB2gBwAlYZUnxWE3GGNpzHXWLBKsAAHArzRunjx4Y33mR80aosgHs8TJzIG9R1fKaRQz
EeZg/saQCfL0xH8MPwjk9CQmUtBLj//JsVgippV4b05rUa7v6diLTOCapF8KfY+PcxtnUp9VQgWy
PO962zZzqvQoYlk9pwvS/WXZN3G7cKgglY9G/RRrKArkG+SYOe0pvWJ+iTg0oaPfKszamAARtDoJ
vZLqLcsGRc3H3Y1m6Ubi7a9Sqebufb5OnaC07hlTGDrK3Y731R6nxau0qMokHsBsu0F9FqnWOL6+
jD6jHUVqWxm5Q/iQq7uDPAaeoSgPB4coyldCjwa/EMFLi4dZILWSJbo770J9VIB5SC3/cC0rCPV0
dDjwcvygzVVkN2OKXjwuk+qv+FzmS6ShV72A6UnYGWPt8jJvmFJagTkDvfRmZtpz7HeVHc55KARg
xY+wG/fpzyyO1RPjL4CXQdjvwJdRFmOxTW7uXg8gO7PRecc7+B/ZrwHEOisoFfGv4h2aBYx88SPV
PnXt/MedVxhMQ8RkT2OIQyEYjSjSw/aRs9lgAiSqPxIAfbnbv7N+afV6fzWfloLDR5+KJtyfL038
gVvcHuFJDjE8EBpidiuIA8nRgD96MTj8gvLnnPQCTMoaMJXYun4ngw/jgp00m7sX4SZNtoJg+uRg
OQjrY/tKIuB/HWzimE36lJ8FY4tkG1zyvt2wMd7RZhg2bgo579dEsxnuCgJTFD7tGzGRKcZmELEL
lt80hwmURswmYleDdsWv7dw14xRPaadcuE0VytvhryfpmhbZhMxMmVizS2Vowkjyqy5mLmxFgYi4
yZGlGQApHI6xHvy3BsI2ElxcuBSu40GO8YAMKvtY+dl90CXO7DZ+InySkuvxmB7Hw/HfIu7W3zAs
9HPHM+kHjLrlQpczVhbdFQXRIzCtlpi90UlZesQQP7HwIJK0rKQZGMl5NlMdj7FKCOQsGeIUUylK
TQ0/xDiWLg6Z6tg2NxRcalPgGftdIuK7mzoO3PtgvTHqsxe5FP4B4zlOlIFviaFKOof0TRyMaIvL
qwQARLMjuR8an7GbIESSsUyk9jBo2+RIEGhmivFIT2pO3/BoTwzxCKvZlJsa7I2OUWsuaUMzZyoP
OisQy05rmxnluJQVLGlgraEi14rjomV4Im/SVQ5CzeM0vsfPGkVREQadWoSmMIOPrzMmASZPCpyz
uiPNp+kpAanUSCx/sk3bZ9dSnOwcNSDARRuqLrbPvxdf7xKaZjOJ9ccZMGNss2xB16sTntsFqKNK
GTT9XGJxEU8wPnBsyAtbo7K0+oKjq1SWWaGHZQQEmy9e4WC1qMFEKN76NNmx2hyZXU+KID5T+S1S
uK8ahWVU/9YcST/rJsqmTF+LMuuXr9YX9pRtZ31m/yU/PppoxTOxJrFSXnuPGwr5K5ZyBAPD2r18
XXfPtwtEbSr4oh3JTxA17LFrMTHaLp1D1kD+sFj+srdYlX3m/o8saX0A1IcUePQPibjupBW0XmEM
hfwl21RxzE2ro+Nsa5CdTufynZmF28RD6qgZm82uynS39ChIlPHmbi7aMus8ZWbXx5ZjQub9kve+
F+FeS2qiJuKnyj6CeM85XqVSYxkbe6EMg7UjfeoSOBaioogfbln6I5TsYtpIt04T575wckpmCoDk
ZDcdYFbspGa1Ihl1KQJIxIZ9jlq4QHoRIu4J4VrbS5wnk43u9P0I8YR9el/ASDNQx0RvC95KacMQ
BNMuRlNz3liNdhYfoYaaOsQ2lIo54mxFpqd3JFgVfAq+bzArV+1K9YnFfyxOh3uO+jYqDbE2OSFh
+5nP4LSQuis1CxgDZUFZOymi0kcpvb8BIOCid7v4vcfJnFc97lA0OUikyV7MR/eAmZlBzpxFKUIH
gmlWC1gVZF3aCUfgJZN0xJ6hzMD4I7habHmwiEYpO7jRoHg2pNk924CQI6qEKq22DlB7GZvadFT8
43ouO7ttaiuKwjH0jMTQUDcWKNgL5Kg1dNGhz0DDRZmHNxdKsgx+YqxiJ/LRPwFOD95fS1IFHAJg
3dRt21rIu1qn6E/Tn14ALGNkaeKSwXsVlIYW8/L2gEnrVBrTJTasjG+WAMARviVGRCrncXIx/bAd
uv73udBTwjzwAGpVkBNcQbx/TdtVcXrAeeTD2RmxXZyTH0xFxh4qS2EdI2+yh5ki/9VogUPlozIC
2m2VU/zrA7m9Za066eWUAcIGt5T2W8DJNWlmgBBc+7Kx6DPgAWZalosCcLgUVLPIuJ4z4bgr9W9X
2Xdr37GI9Eua+BaYn96TrrVN+GQjux9mTbJA6IqZ8AEfTZuWgdvIfh1ISskkBPz82lvp+eegEBhD
1c8fLJD2gWgwLOyoKj2x6eI5HqdX7JawGPreYNhVFRKI27yNcm/MXJzhb+WOQgmyGga44rrWrr7+
m2boFCWjd/tp9RkCc2g7AW5WqokuXU4qIIkjdKdcL+EflxLmml8/4gv1oB3GaCMd6AZchxdrNWnz
UrUrPWkCbtfpYvGRd7FY8Z/iu021sbvyYskbCGwFX/VNBlYOQm+FZ1F7NELaafXKT2z5mT/gDIbe
krwIE1VVktGafSTnhODJY12wnoaYYK7pqROIiPrtubtbzMIvK/ZMfKkM3WBgg9ObjNj44TtHK2Wi
mC0YMk0e1l1FJ+jBw1bRMqYHBCLmjEzZ6CWauokExFPsVjjtbS3720Fus+LpUPRWir/PlnfV3HUV
p9CFMi9dF8IddS/qQkxxrnlFcM/0wsyTYcrgxBoCYcV5/q4D1W3iBPSzCGXsJ3fxme6v7pfEghW+
BXVJhw7mnXY2dR9Vu1xN3N218qGnwHJl3uCwa9D+jyCF1Zku7FJ94V6aSm0pI+dvWS3tpNvpb16O
9OZin7yXShZi2xi05ZLK4SobtKFDSZ+1uoQ0lnLS0Ikrcc5QpkaR1zJaEdcXEYdASRPqlDr/lN65
KcYAB/jMmJ+XW/3Gkn4SHX6nXm8Zac7dn4/6TBCjaEFPwTZ9ox4Vit+nMt6SEZi/lEk6r30LQvEs
gYPgxnZtDobqN9bRpPiZmxldQmGv8LLqM0CygaC7WgwPpvi5OLYuXxPwfvjLXfiv5Lk0YIMQ3xs+
5QKv9xsipOQAd/dOP+TYnOWNUJyIIefwY2Q2SLm/QEhpUm5Owp7olQNFexhMWNsNl6dm1/gm7v/O
FyQXFiZMo/8h1YyrgdJTtdEq0QKeKEKVu8BwLbOxb2q8uwtvK1jtyl3ssGn4Xay9uIImZXCXwH98
MrDUaAFV6GEKG2NxqIbpbQvV/IptvdEviCp58dEZsL3IBFe9yfdHPtlOmFHc2XEjCtyiCtrKb6J1
ARJ9LwvjPJh+m+c6VBva5zAjomgUXd6cQHbLuJFb3pnArr6iVVd9Etwtr3d6lpbcasx/Th+xQ0Ft
1rYogIZfh530g4B4nLTWhlYPwcUVk57aBqLbTd9L3xV/6ISQrIq6324PMulzki2uvL0JscvlQ6Ka
ya2aHh72bpF+pVG9hjqiCo3ud8MyTuGbf8n6xT5Lx68yTl7E6rehYev3EIWoaT8XSN4ttw5RvXgG
h0rdUKB/F3VhOEDzOsN07ywcctUvI6xdkh6NzKamwibsjIJElDDW3m0iS07O0OQsu+5NFGRfPc62
W1BG+dBqeBIH5oDMgHL0Qkhoai+CJFCCFtAvU5QNRHMq62KswoGthXOAzkpETvDzJ/vONk1TW5Qk
c6V9yfKOMPpDSYKmqvXwmp1cGJoHrwFNMLAEba4g3VE/b8OdcgLW3vODUSm9MCIqcl8PXvK7dzMi
m4xHDb2Fm8JwsW23DkAjUTCGUl7FgcWIm4bjvaXCtTEIsRzXiQXvVYS22y2Xn1c/XTJ9f82aC/12
mcIWKpeDQ7CJAKEGuhMKMFJQPwJK/Rhpkl4W0RaD4iz93fkJki3R8xhrf36qNEnWYEGzY93YCgKc
Vh3Tuywtyu14gCS6GJXaGVEpIab1y6mw5H2iDLvBbJd0zadX1xzuBEajX0ytW3jpZncDgDOmCdv2
GW35/gr2XHM9qGsufYvQRb+ZTPpm1Kng5oWUx9UuokI2WtctQCLFOnvqV7hda84H7ZoQoICCbOHx
4dlnQV2+Ws/X8NOcEt0nbbOEoe1/3ljRzqABZ79Q3nqn7QcYYz7FlJLc6ltPhYpPi7ELAzfktUuP
cl2g3nwl3u5ALcmsAdImJ83fyjL+D5xZBz81s0E8LNB1xkCmgVLoJPHEta3lraDSZ3bvlRIjO1rl
eU/K+255+t5/xwafJJID4Z4ky6fXf5J0a7+VZCBzR5D5aon+YC2GLIOGQfLOs2Uv/HL2yl8WbsV8
K1pMe3ZbfLAkGbzqrr74DEHfviQGz5pGUReY7BwLKv9Zt2R4X6ypLQNnANfHe1rQ4sk4IbIv8Mx9
hYzIYGaqKJPwUVs7U89oaTnOb2bZDk0MNeHElEt5I/gpCHlbRBcc77XkCRTHzZWG7H+59rLSOPoT
GdZAJVJFqIBFOMi24YdoeGxl9RWu9y6//Rrq25WLjKTGSolsz0ro5YGAzER8//b1Vgev4H5YBNAS
v32wrkrciOZw9XT6dlfrBAEiW3TR8DOz8p8jNfxyUceRZYtqwHTP494+UMmBsHRed4TKn6SctuIq
Q8Jq0pMSIa4KDsEN0js/3/8fXDgNELzWW9GgJAB+cv+fIGMgyPXpkgoRpEh2k/EO/etdQFg+5TUg
8EPKV72esWf5QMYs5VyzZ7Q3/zHspCVEt606cL1/jpXUpkSjjSRzTDASGQRbHiN6Zau7V0NP7A62
Teeu1K7GClok+r0Sq8sQfr6/5pV+WSTJsiViZ4JKocRV9NVaTOjX3P8Q6UD6/iYj7gB2aiDCuSEU
8f0JgD+LnLaHD4Jb+hrhXsgNOB7bo/ZU0epHPrfcEA24dgIF52RAw5b2BiEl7bxfk1aF0DkvF0CK
nhFLrLQLnBQDg0wQQ4TT0TrmMSG4ZpOb3y0MCxqWCQ2E8W1mwNk29OZBNax1m9U/X4322eDtjOf4
2bwA/Iibo7lGwLnuRIDRX2Dah5OgLF0zbuS1P69ESpsUJ1RIWryUbOuyV8c2ZpDHyyFwz6iw0hgF
25BC+9lcDfHEkjvDe2TG8zdUbaY8U4pasED8Yk3Oi3UORFxvk8rRQJEJ64ryN54ySyhevFFjwb5k
I/hWFKnurHEUxAek8PzfC5KURKJKRWPOiktV85zWLYjZTsKqDJRmUcHShI2y+0ArXd+H67qIKNm/
zOOkzTggR0rfcmOruZ2HRr+vGwEFf8ZbIRxdc0YHyrTd58QIjSmvQvy2lVNvvEuerN1IstpDaE9s
VxZqqpzlV1ZlEVJFOcog/UqRMyiaO6cVBTYO/zGaF72WKop4delueIVRpq4RDauXe3xZ8ettT+xb
ZwSnHRfJXWitBXpIOiZGRzffzt/78Ybpo1TcJy6WDvF7aLNCoWHLf2viRlFkBnzoI6zs0hdRtGy1
8EaEeEHSd8ty3ZWi0qKzVxHMDqoXB6BtSQTjfmwu0oafJ+G9lJVKrptnXS6BADceRf+1QsCZAFE4
AJn4THyR9NV74zgtqxw4xo6/vmF3UqyDP+fVY+HtHCSLEzo0e7SlNa1ja1Phc8Dg0nhsm2epy98V
O7Pjn55F3HLhY3WsP9K+p4Z6kb3NNbivJO4oKjEuPdiA+llIE4jF8fWDNRvN2+xCmfHxjyD0qalV
0xWsQqzJlyEStT72N1yhYPvfnsKV16u+nfbEMWioMzQE5r+NZsIfrIBcIDjgqXJhiZfBgdiMS1BD
Gs0crVeMp+eb+r9xOFk4LW7Gbpw4dC+beSIY+pIKqWvSu0bqxArUgkySBWGBQ41R7+A3ID40jNsp
xHJZdqsZUqfEkRwrrA29BhyWZ0kDVu7blMreNE7PlKVuOQDqCni783cWVhg2sADNiMfXz7SjY8yO
5ILd2+X4CEAzWCMlIER4eq0VrTOtZ34iPqlvep7lM4COPPutPjYpddbvXNNFdDCyvRbZuSxulOQd
Fzih/7XgBQZMFpHeHsuxu7932T+zO+IZ6wPQzj6ysc/SdRHUm+dFNUdxW3LyMLMocm45gns8FCvN
B2KeFNywyP3bl1OY6cOW/91jlZL0s0rO7esYGhoYQ9v1zpcqpNJ4IfIQVSaOaGk5Jb2WYyxH7A5j
qbTjXPoqLZUeQm+NR93IOc1ay02lStQOVBNwP2FkmgKoJamragrOSbpbqJ2/7twu8fhVIKLwrdp0
WmOpHyMwRaBnoT3h6LfdExkaMDpzFtbbIAuVR/PRh/MulCZmU7cjdAKesH7sCu7idKH0RcRIk1Sp
q2ZE2Rwt+aVVX47slaEpv0JYR87AGWz4mcMzkV90q6fVtGRKl6nv9QALYE63FQzdn85D29HoCu8J
INymz/uUVqERuFb8dp71Cm72XiwkrLpH1EcHa9iwrbHJ4P1YIwCYdGpWXu2fa/jfTjhxi98DgOCG
nnoFX3t4OTpCme8KAELim8E/STY3JvdPJbB8YhjBw1dwdf5EcdtayojXc0mcirLJxIYGnB3pVM6h
B/RD5nAWnrXhCn21cIUh7LG/ZF08DuLtkuFWLD6j2Br6/HEWak4BCgbpnTquiVNiTDHlX1POvSi+
YoGHRoqQcTritP+Ycx7Pm4Uq0TtY1JOLwjreT9wO/9OhNhE+Iat2+npU1rIS6ii0QTjXCMMSAh6+
+yFgQfWEeokKo3MLGcRlOsIj1C6PDeQEpVi2BgQo1Y3XPaXjg7gNn8sQP7sqoTKxUWhCaHMXCE+L
cRcGjozll9YaSK4oJKlREHsZfmDSRl3qoA+N8cY8IP9lCYTjBVdR4XbaIXtadydwZPvwYwwEC8bF
S+1Na4yQBmcOExbpdqlRBnSQT1c2ykyksmKWeIssR2VumVOhElRqSTttX8AqPZ6a5CHT/ZRx9JCp
M5oxvWnmcQnthA12AxRSnRy6H5+G5tlgYzhnTfvczmWlgODGyZ36KiT/HI70EVuhWkpUOGbmM0H6
xvSfOglXyeKMOUOBCz7il5dc5oNue0ayOCgRVTO/PlXIu2EtR9W1mizLTOBARkB+kGkjwE/Jh7op
QP/HKvHcue4GuO2iduCWr3RnrOOkMphJVpUxYWCIoultrjMAWgHIqvT3UqSm015Ivy8x/sEr9iF0
kyF8GW314yQ8Tv2PlvVJLsr4iRetkC+dMPjh+MRmaVsL3VSvnoyFiERH6i240cuqFkyBhI3GgXtj
VAUIwa2EIcbu/i6qkClX+LxhlQUTpNcALX4818p5Ohs23ljORZCxIsEyE64kVtePQWKwsGseJSHW
SN8bUU0UDxFyYYEHMyievP2agqOmUEGNmBMEECQZ6jzUOxTuvxHMixARdg+Xs1nMw0I+ZOwuDa7H
V+8IfE9l31QMs7UBduTuTiYrZFsp0rBCK2lolCQmrQLklP8N7I2AbOxrR7bymMEjacGNs+UeQDzz
oPRlu71dQUuWRMKu/Ajj1gtKdlHNlDrLEYRnvNQrfClpekGHvN37Tte3Qhl7FaEdDXkgDowRjrEA
tW8TUmH5ZlBSwQDUrCBGNgcuTUvGxR6mPpHm5CShPti1WhG2twKcPm9Pr+jVdylts6FQzgfvFytA
djoEaHijliPN/NLmQfVUhQjEytEX49G17NgbLOF1SR6781mrOzj9uicqPq0BoiqM0dPeGyfcg7gx
SgObmzh3EX9MdPL4Pw8kgV6jBIu4iqDbTGTpk72GUuKYMq9kcLZmjoDR0UPCblz0P8Muk2xaE5gT
HgmuEp6JaG2FhSYlnrHlCEntHINWjPOXKyM8SoCj1FCh0McbQEBzkwGCnLlc4nXzvMwyX72MilpZ
Lv1yuc401RlHpXWiLfvobQgdqSHWHcX+Hy0f1RUBF7cWSMaahWznFG6KZ99e+/Lmez4MxGcog3d5
P7J+aCcfREc3/ZnK1ll04Q/IJDozdL5Rhd/5j3KtMRFTSsJDyy1lOwQO7f5ZpScMJcqhn3RUU32D
E0NnL5mQgz/q5xqoryWNtv8Bg/0L2CZBWsizLhOF1yjM1XHRt6pxNzW/JdYshxhwnGuUAEPzQEtb
tQP5Thmeyu9VhmK+OVxdt9nkG3+sCkc2AoUPiUhKgEP+mE1rEZTYzGiLOkA+j4/Dr+5fq+WOdHRh
zkw8L4jZ1vPFI0A9EeciFiE4Ob9Q+TbhiNSGV1qr6EhUZTML7e4Oqm6PiNKS15qucmzLk6rtejzv
ci2FqLEXxjbIoY280BzFB5PfOYbnhOYn/pEKam7Q9DW7SFVOd9NavqrjUP+M5tPkP2PNMqYONt5Y
BLMxmqp0aPh5l+Qa8+blOj36b2Mlrbmkr/Oema/oTDJU+jkd8VfnICZFOTgnCVurtEYH1Jensvls
67OY96QUB3flrfHqpWlu5euykr/UG/eR65HsDpXW3MtdIP0KyLpQ8RvGKGk7OCybUNdc6DOYJLvd
PcBr8QEo2ToZnFQcvUtm/n2MHf67E/3ZlZZ/cnmdOIYto9djFejZ7O278fA71keDgvES6cton+3i
Dc8iuFjnoRgR0VeRERXAP8J+zjdNAVXLZq2jDBgf0MXtPmn9AqyaN/r7wLqQvuLPoe1IU4CH7ROb
N5lKhVc/4ZparQq9KD/J62QWelVjpABdaw5/UN2R+DKmr6HrEuwXf0LaqvMUc9SjCbK0ljZdTI6o
wyoCUzcedsY0UfHy4410/Tenhw/uqdO7X9+iQhl1FkUgCZfxGlj+2Gih9UQ1n6JDt6uYiuNE8/uB
2YurG7W0Gl6WhyvILKbgqkI2SlPjgUH1gl5TK+r5QjSrKhzZM387b/8jBAmybH1KKmnk2FAAXaCD
8PFbidJAK0l9pFSse6pzIZwamCePDbJ1Hl/hctzrJQ4kSCq0mz/ebv+bVWXiL9RYcvEWkVNyN40d
7Jb+H9duCSD/K5cWiWEn2EB7oE6q26GBL+CUbCOl6mncHyZ0N/XFAOrNzjX9RZzKVmi6R82Xe+hW
AOABf1f6aif62iaB1Kq5R/zI6FZuNJXX7ct6asAoO2UKeR8YcqaWhPcCXW6aWJHhqxWIqvvLh9HR
qN+sX2i0tu2Os53+1TCFukc3lS3mJNHrHaWIuQe6Zst4t7wjvDAHi7/3ANhIJKWPidakuMMBoJhL
fTrZKiQzkpjcYYATBXt6vVnS3r3F9fq3W4/bJF2pFIg5fW9oGW8x8VATuaE0E+KE7Qauwt555tI9
jzdV9jB3AJ5N2/k1IGYckyYfPVEI9Kj1XFGFYJNlud3KrA15dPALl6Fg65chd0FAelfmjvYaf8PZ
8HWOw/y8xddQSxFfzeaiWyKcDI4BhbdWkNZQrd7URMmMApxVKYpiS2JcCcwcuRyx4hpVDRE/cU6U
3sSjy1RRBw04hgbnM+IuwQX7oOGsivHjTKohdwZdsSPaA8xR2iZlbIUzCSQfPgnEWcVjSTYwt7l7
gibO5dG14SJdkECKdY7/hQVroN6fmbfpAYEwW9D6O1oCDu1MYmOhdBuvKlts6j+BPmQaWtJ6L8yL
rMKoKPUwKdmEjcXytmkFMuFunyVZTqASjIuR6fzvTVW1cd5AoNUbWCuvhlvyjdfdeQafvY2LOZIM
PTUxX6Y6bq7qLwTmkQ6ug5G4RacrAcR1vCiLVs7MIiH4+eCYdv0pLd5NWFRQK7LULYuj7Up+Mdqu
Ou6EWOJB+nYPGlcvKyrJOpL9sZLsri0G/p7NePbBIwLV67geKxTRF7RfwypEtP1VwvD3pYa01Vm6
4jcFDQWLW5iHe9wrBKfifYyAA1zsAlUGvgKrN0BX24jJTAselcjxaDe4PBsiyJ4PEFyrSWPvm87Q
4s+VETGAze54kAcC4mSh0H9qFZHc/UTo0P1rFBcnpH3aRSux1zp4Tdk07THRSlYau+JMWUgTz0EZ
Of0KQPc6KHlow94SGhS4H1pkiLkM8+rQijwmf28lwqmSM68eBUUjyyxXDAK5UYGu+QO7T/FqdTFO
Pjz8oj+HwFs5XB9debPJMNfu7Ozic4w4BJFhwG/5SPCxB0XA4Eb45ItPYojXxCJyKLi4VR1tTrs+
d5y2gKZSrWQ/sGcOWJWjVqaf8ecI0joy+5iiBptPdwLo1GCNf/G4kTPe1TnzcM/0Eb/Zsy4iLjHa
iZ1yFRKIheu7IXlIwmnGszisvy+V8c5brQWsgLQ2akpgHJkTfimQsATiibKnR/II4JiWbVPXG7c2
RhV8tsfwPjSnlsSxVdOlRmue7qbv6JbrnVXL113t2mpCRxNK64OrwDDsWqiL702bWaLBMjtW4qrP
LDTRi5etFRaVJZoG1OuRk2e/NHjLDOibufwsEFS/m8bpvBSdjvL8b/SfajKFzP4Eu4P3no/iUL19
C5yWxWRzxSkbEqRMToPkPc/Ad9wJFfqAj4MERvVx5Jyui9pJ/v0vOu9wxW/IqL5NO6vqkBqIsxDE
Naociyhbl8XumoxmmiAyrC4rzgEaAP2fjCeAOfwa4TqeaVFvDJ5NMluzJEuuy3IE79AAhy58YAKO
P3FFBTGA9BkOqnNxfYJ6v5FWttVYzxTg1sW1GkpNa6D3Kug0EgWAnPXYkIh8kW2O7nXj1ajAaPAy
OEQZMj/c0MBvJhOM1qA7OG39SrIFW3mCkbny+O/slkc8zGMMF2aqvmqZUMWGXSXSM8t30DeQcdHc
PfzbSpTPmLb4K6Uf3ZOPY7l73Gp7JPweZhd7hPmaSkMqXLiRP8GGZLd4M6cU4xn+bi/RDZylcToO
rx9K/kpw/6bRmQ/LMj6d5hNS9M9Vra+jm+ADludJ+rthvf4kvS/ESYpYBJQCSRimlfDUQj2GgpFq
7B0eykoPhg7I6DX/t45P1l45Ikhgy73hxYLX7aoF3kxFMkrbtSqc+rqB+hRdaFEeX/wxb/+oKJHY
qrtgH/2bB+uHSZsqpCPHZjZKyd3RnOjGmAsu6KMqJ/3UDOAHGThcK9PMGy5rsQ8RuWaNtXjWm4hu
aVSdtLhRdljkrpSsSZZstOHJbqlNu1jYi4hIwz+bfEOUDEZ/UnSaOl9ZPl6XI9AsBxOAKmoIbuau
nmPvr8LyekQYm7CRcJkrv1zZspgLXyttieHWJDWvB9evXNDG3+Qyh8JOVlhgggbe/sXnRc4Z3w9y
NL7RvjMhjqLMxRzRrENLKmeEaKR6MnFHLnG0fKvfmxIxm7ty0NBB9wW1IXjuIbsj9GymvTSTygyt
VOO++rEBxZCs+bsy3C2T4qs5hRnIWYO4YkxL9hMnSgF50vCmzgBcM0YJzhdm1CvDwPgiwmxosneY
3WJVid1nHnkkr9L+bjFA9UA9kWOc3O/EOp+qbvutaxprfWYf5k8VrEGLnGBZUSJ9BmLICSSmQsNR
jcWoBLkro00EnINJ+7on7OgZYgg5BvTxXJKVCNU8TQvikrIi9McLhK+Zf5ie1vwSHoIc+SVe50PQ
xSJkcyqOFXe6WUm2+3Y1nW0WkSgjl0Ysw8iJOEHerb0sDF8Uwyc7scoOYQzbEEmswUw2Rao0VX8s
XcbNW1OjvkqYV6b7ntWgHVWHn1k2SphDk7WYqrdGlHaSnzWq2shglBY1dGcxlpaRGrN9ScarC68j
eVc3Je6uL0r93V/12bU0Qn5ajc2EnzIDELqa/oavHFMkUo5OtLl7KBTdyQm/zQrxH6abVC4dZ3S7
f5f19X6PCakQRSXKXE484THY/DDuvQvCdm7F96YFAMMFWb6LEA/7FgT0xyLJXOnIR9NjYCCgWEZJ
RTMNpaMokmZ+Zpl70aApP3XwleYvHyo4TxdEWVx3Og5albzJo8BdArOI+rgRMIzWMyv3COPalwQS
Q6ByKGLP2MGT/fKocY1iSUEIri1twpwzgdsi3CfRbiS728gn3NcRIwbZB2PA5CRDtX1/yqJJkwVG
mQig0XIEmX0rlAPMLj8fT3oT0nifJCreOdKCmtWWgkV5NX1SCIbPoEY7ewqf+50PNv3VxgPeI9va
meIpxwyLjDolFtpm0cP6BbXwY1dFIVwfCUPJNxwq2erdRvbfMXsMdjer9utGU7NvfkRR8DjzoDWr
rvoyv/X99doBCWRp3sJ7xCgsqjVh5abaAPjrR8ED0rPotYR9u5nW+DRHQ3dueAh6H8Ql8+uDdlY8
kj/XmOxl306jP4ZUEqHFa5aV3dzUNHtv9hdoMIybA/6eEkS4VeeFIPZaV/Braku+okVbu5H7qmOI
plJ2DTVpljyV+F1En1vJK+QDLtzNdMaLoolFoVOvehy47pIJGpFu9KyRsf6yZfgiXWyTdP7QX12R
5yYWjdOSxkZnGC6ypU8UVqV/NBgc9M7mrs4ldqKYJ8jALPjpYyksx8yOc3ObxltFjoB/2WpnC1oZ
DrKrx3CAOEBY34Pn0iPiP4U1Ux174/ZM5ou1Y94wuMyvXj6oTGwEEIJy6fVRebhOifg4mQGk9JzY
vY/OYYFPCcH3PjT0DBE7Hha0UxUQx4y+iF4VS98O236gQZDJkZNjFpK9q4ShksgTfJ5j3xZ7q/pw
dnAy4fVqZxrRDxO9sQVRcJIn2H89qa+jDoAR8WAlE+uHRGfZCU0y0WpN6RVKS3ZQagSEWHOOztGk
zc68ocGXHrKqVaLDGV94hpukVijk3S1knIVGw84iWReg3u+IRJ6/e5Vc464oTW2yAbx7JjlAvo1g
5n73yCdcTAcrRCs5BHAGSaCzin435U7ZRZqYETgSKVy82dxJ9wU2em42MFtbyK5BGHQX7PvVSf9h
vlCmehUk139snpYA230Sxn+L1MZhoAjZmuV2OMyxErmf7XEK5c/ggoLKIQBiudJEKuccD58hDXpI
3zoIC1Y+RmzmnEtV2Qj4K///iEGaw1BoR0As0YXyvE3IEr/UOXYfbHD9D5/i/WWzBFcEyBHF25y1
PgkY0O4uEcRqWGCqh0Gn2DWycxKWkGNNNaRB0xZZt3w7pq3B4/nvx3mfvXCvw5nZiaReyJvSPNg5
3sMo4/kJz/+O0VFl6F4nxZDxadXdoqmdUDlUiFmW46FwiNlRH+UHLJLxhXvkrNu+CXjdvktS1/OC
6V0Yi/nTTDXzecs8AIWdhGxpYNgqPxoLgAzw5jfWczQdmtxlq3ZfoTZxyGNXOmuChxq8lBKsViRq
nF0NsLEAQpDA76MOpIfYuLUO/OFzQPJccQIFys2Hd2xQozw1uMndcsM+bX1t5D/3I+Fr9Isd9y3q
rgmUZmOKtLL0Od+GcfszmwH66lwOTn8D+0aEwYeIfRVSKYCSkceC4f+ZK0/16to0u3iI6YukaoJx
CROFwisqNONx3moI0NcVeUSMi6U8HGxjjdy009Vc4t+Y832gyE27HdokxahIMk8YGyVANdsaozWE
6lppm1bbZ53JEVAyOr+5om5LhQr8M0fSFHznz33xM6cqOwdbrlyOeyMxAOM7ZEhzr9AoW8hoFoDA
dQfppLo3P2lJGrcSjpBhTBZNDdYdicot7W6/ScAigFqwAPwfhrboQH9dgPi47uawWTdu8X6MeSli
hCOat8bDkBN3A032paErL7aAaPisuZ3aaCQl820GsxkLI6WYdbzu/BhNB7cE5zYE8FrVgfBwtG9S
hbJeyTVP+HJgFSQhtT766QdTwHUxG+73zalK5g6rBGKSEd6IvAo/pPUW9pqqVG77HFQFxcXDxKTa
U23dAv6ORTQgUAI77dTrgWsdoi7SOXLgQYADYRxJbkPcabY9pxdJMJ/gf1EdgNy7ZjWfjgoQDVdg
8j0OtUhnzY4ZxFIz4vOQAOf3MoxHGA+kljG5xGgROv6dnrvABtWIwHUKVk8QJ0iZwkfCy93mQvMr
xBM5Z7sUM9S3vNC6y/s9LwZT8NLrvS4aCdD/GL+yGpMScnbJEZZ1WZIhLUrYfX8rrq0JZqBM8X3u
RdYH0cyYMffIPfLWEcQvyAjDbU7DVvCcoxA+3NUSg3/iMfymyhcwl85fXGnoemBYZYovesGYuW5T
QRN/4ZT4No4xT24z8DmPLc8/Kmif7PVEgaEnTjJxfBSP0/wcGUgnUjgKMOf6Fy7BwwYPka7j+usM
MfFPgKDKs97tqhnvwasLF+XSnT0vSmNdR6A5m9SJISabyc5skfQb9YCIhSGzWVnaR4fFXHUmmMZs
z4vpUVYoTqE0M8vSGAivykmSExxszMZaRptmNbusN9AbaXLOpvDCwNkGB2eWki/HjBPSNut5+OK0
3hkZTwjFwQS+dMcBqj1WJkvAAYGHSO8LGjJ4T2VJYin3nccB/oDMFZuqOhKBEq6e5aKKC/DudxiM
BzQksg2I8tqob8ypdWiFEhK+5t9PXQC4vdXHapwk6KxI7bLCNrQDTIgyghfauxu2REPyIltpY1RW
yasqrqcVYbm3dJJBwsz8k3G3xXiRSjdCShhlEa83f6mHh0Yr7xCqyuVCGIPsH45r/j7pwbmvqH4w
lQ9Udj4k7ECV06KUNbydmmOj8YYsN9Lt3Z1HIvQDKr2gzm9yRuevpsw+8H2qHDMjnQfcEOekBp7B
gUW16To8ea3IHvdc9uMa8lRckJzc2dteSgJFTyASYWtOx5tChNHLcMZD+opwQwkB2SUdBYsp7nED
E7yhFGeFty84iHBB2gxT3li3HmLxo0XRyM1IrovuoRevmi6LPznmLA9Oul1pVjdpvWnkhse5SW8N
8VJlulkMctQY1+tFOMeqW7BkeTFR4BlACJ6Sm+iNQCsjtQ3HFDNT5HzHwqTJW48WG4I4Rcwux5Kg
nwl5AiztCXbEe560wzviEpQNZjMrG+TamDiJDEYqgLQe/QG+8NQvoOPPgi88lddWbxlZGzMTsLVo
mYxaYQXNftRLaDHS6rY0Jq+sVwGNciHaUWUDTvOUlMIsef+S4BnXh+K1vYvuFGbQgV0B8wp5E3U0
+530Vt5PJrxmBQ0wjKIOSsLntAxr2yqDQjKgIgRHUQX3wf0mHGT5I80K4V3QogM6nm8+dibtL3cT
F6XnwGfEZKGDs0rNN8cPDGSvtf4EJave4cGm616bWaEtLqMHO5rBC3wFdn12YOKTb0RiWcMTgrSL
EfqwD2KKi4lqZ23S+TsIqKblkrQ0rQr3qtL6Dd5TY7oeV0PpQ3bQ34KeXsEqafu4hohVC9uCellS
d+4vEwtyQonfZiq0Mw0pRFX0+66kU+c8wjnLkew47oNjO1gg6jhabE+NxQdfVIFarD1WIIi50qF7
jt9Zsn1njvDQ3KQyRTyR/sik1vSFlOqtPZJYunGZiSYR+/VhX5xC0cr9YCoLIyuZepJRkc0eKZ9R
v+bC5UZyYXKwjWxa46grfCO6ihL6qeM1YZkhfDY6c25aTD23888+OKuz5/wxn+6257JFBgjgX+b5
HFXXnHk0vSeszF+kcOVlGFlNHmPSJlxoCYTPugwkK9mxul0otgvI+itqDNoTYqrJkE47lFtyImJO
mgvO7tXpQ7+q4X1RivtoNuIRRB8vEiQZoOZWTUqssM99fxOfNKDMeGMQ7sT1eovW1nHq8DzLyN9/
V5zykEBm/5PSyV7VEkYZ+9Jf/ktFPDyOUfEoqM5T2j9eGj9cKkPMv/qyrAZ77+LVp4MRhUOtKAdS
W+9i9WZ6sOv4SY8aDP2EPf/LK4R5LTEoglVz6Cyv2RyrTVMsmAlxbIO3Df4UHtYsSzdM2zDlMI34
Y9213y1l3TPpEjtGZ5+QlCGbPi8eVv2rVjwE+WZaQJFFy6WGa+thGMOmMHEjiV05AR9cavq86su0
ymqpNJrsVbN6EqnXS+zC4Ay6EkbgbQGqWZr8SlRpzTawgdqpX8JZdOsJyUfJTsAKjqZlG1Vbe+fK
yllCmLyX7MMWuCpjElvky8ci4gKiuNKYCp/mH1+2Lhc4xYI+t2zpioKWNZUzA7bmU+DVtaSF2Z8K
Ks51FstNB/3rvHFFsldwKG6Cim9oW6iIW82ujsNW9La6PpufsPfR9+oGJtCBpNSvu8DFCoj8bDYs
V6V+wMY/AhV5S0vLKviHmbvQGe98kM5EqLq0MvOeIqFdRkWxSAnA/cGVlyPWTK9jljCJ6/unuiNh
iKEY2FhhZg1qTGtfwo0dl/svXE+HJEW4Mjoxb97QFqrzOds0qdhNTbgRgUP7TrvjsaoVy/A4Hqdr
U1l4Rc7boEjhf4t4NrC2LzcF/Ifb0kwV2Xf7M3xDpBCHxJkyVxRh+6Kx0bGhsMAdtr64pjHd4KFH
14GCHEhFsmPuNfE4I/STdjFP15js/O8HiwMe9/A8g4sobCe7ZFhScRnttPzUhs12WdpoOs3sZBXU
7JRQ7iX+eORceD3cHB5TfDFfjVBv4QLc5VbH3ir0MLrA/BlukBR95mvbztXeB2NFmYhU1Tl7npHc
FtQmNDf313ikB6mjEvJ38J4z4Lx/RZY4ixT4LTafgcFjObMzEgHmsccGAY1yGCQLk4wHdTv13r2i
MLhmiAWFlQYe+iQZSKvvWFBK+s2UAelznVF+0PPeXZUY995Rko536TLoDr0E3NzK35gBClr5hMNX
LecFa4Iv60TSt06C1FA982ccA77TDGEncswhQGXF4gTEMFX47cW7XA3QCkNb+0u8cfvFjApvzvQx
D/hcbnUR7R+5J3dDAQCYu9Dri89k1MO8v+U2oA/n3VjidVI/+eUIupou888L6IL6ZTbg8Rdfz3DP
k4Bpow9y21sdtRgxaQxYwTQ+/ZWVHITNmwb78H95HFIaTMDDx9U/NLytmFjfaxqcki/J+q6oZpmH
dk8qFtiWtPyD+pKQvS7cntYmYmkjRg+XTOMyt91fYRWVxfbXy2+UnUqrRi3iWbvSzbk/wwKFZaDl
I89bXdwLtuBIjjrMfZHcmea7jBRLbF07E0Z7zmeeLRcAqJOuizpXjanBVQ52RfHfrUgZlGYJu+VK
aNZZSiKmXMswuBb4abwxysAw6Y1zYnVGibSCNmsdGUzAt1RGgu70crLJzO3w57xyroQW94Ba5p4/
CkPEM+Y5es+wfgxXaCyIu0yS26YvoKZ/nt/FnJan88p1bBRiN/1IglmBwucOZTd+bGQvNj1Guhly
OgqzTN68viHOJSPEpYD7jMWdKDy0FPuAWK8jmTgTjip56A9/YSu6tJVl5YNa2YY626fVkmNUFzUm
KwMoY+0psJ/+9G551JhgS7sG0mr00EsTwhbp7P0FawtFUoJyR1HqSS1J/gNVmSK9NlEI0hjglgBH
xJm+B9BxPLwiZpTIw8yfk7esfotfff9ZAf36WcEGMqd25UAp2XiHPcUd8Sj5u8sk3P2bczoLYfDM
m+Jp9wOCQKy2A2VTjLPTr3ho26EosjIMLp0mB87NfK86tMjmcyrN3pDkDQ6A7DhtVIbGPWBQROgS
xh9FJP9UpgSNB1hyaQJWI8DOtAsb12ddkY6Ir26ZJDdv7OFRbKYOXXIquyi1JOjzIxXAiCgGNFdV
USWPlpn6WKK5GAKXHbHtHALXYXQUraaPCf8h/pNVc1A8d03E1GlR5gB2EScxMAgus6MeYd1mzZ7H
bkDFmez5SOcSCQMa1U/QtqPkhUSLLVMUZugcIq/l9M8exU15QkAwBib3rKt16turtIQxjFjtQIW3
u9QELtZ+bJc8VMoyetouxvvsUjJlAhjjDoE3SGLxj2rSv7Lmtm1oc6/7ALGigJ4MInjo1j8cLW2m
Q6WRuhrzysDt7pvS/Pk2RxdJs6cH9g91y5LXCkynszlyuTlquFVDKdC7NBJWPYcOO433Cjf+Kfkl
rniUmwojb6hp4P1elu0Ztj9JvaJzPBl3cTkDI3MZTDmARJprSMyhjayC3+e6tWhNUZxxi4nGEwRK
+ViZIc1TmrzJy0Wiy8RrZ8ic/X8uVH5y5jrEf67VOak4r4oOVJousIRXnoB5CR033c8btnnNcDQE
2bLQnYY50nHFVVWt6TV9FO8fZtGNSb++ArlzPe/53l4w5CAqpx+HLnVs2rby1/hJOtv2rNSn43qT
pqKNqiwQSr7+5J5SCTrhyvRwn0POOvUeOwppOHcB42wgQLYtBMoZTT6YV8YaZL5AoapaX0WSkOSW
6t05D04thkJVQ9JkrfjmNC2+TNyuYnPrdL9OQcW2OhirTuoeuzOKVjJUNJoI/H8CUHKWv81gbewX
NAw8MZf4PS+vdLcH2IYSUMlj9LXOuI14/ukDSkuIxfkO4ROJzHmgTOKBOAxWoOVm1NaoI2Ao+UVb
ZlYcVwQ1uttAPn/3L2PtnN2hjC5WuNdesZUxw+mfKf10M2XRuYe+n8zpjGCmeTbd5lWLtn8Iu1AA
VLENdwpJ9KZEpoamzHCTCIyGItwz2t1yT6oyAzjDPkke6Z3gSkmfUYPmpN+B4obeY8htYA54w9Mq
AqI3MMedUX2LgfnpAHlPrU+mjXS7pAWGOi06XCHp2eS1mWamnjKBikThpaqtSvQCYC9NDs49hZP4
9sxrMI21um6Sj1WzeM/TQoATn5xH0JX8AmpF8ZRoot8/yF4Enpc7iTCbUFQLj39hdG2jSZYNioVJ
v5R26Cm0b1VoKg9eG93kpBwyVBBg+ZR3jXkNv5CI8clk03hh1gF8zkKrcCUYX1nAAzBRsvFEX4ZD
jcaaSCLFIcgVH4bmES389/0h9wX0ryjVVacr9AcaU1TitHMTvtne6E5hUbKYseVm7K/jHiJq3nPv
vKO01/Eu/FbufWuU12q2CIVXMBtCnNLOvh04wGFDw8llWc8g7A0zOf9padvdjNVwJEDruyviK4Hw
TpeGq8gNkjiU5K7x6GK2yoOu+rKYQQWA6OmXLvDaqLosQU+lj2k5+YKcZzlR3DhLmhx0Jp+zwoBe
XntpVSA/gpn8MgDr/TDvJgE7M8ho/ZYK+sJhP4ZB85VO5Bo2ewJkcAncxqLgK10Z4wVHZ1L+r/x/
0bxYN2FlMDSzAiSmBuDXC5xhikmu8ey8pvybZ3pCLyIQmgEJr8/Wxj0D20E9fVDquzfMZSjc3Yb2
7TkGmSHhLGHPViKYOI+YGMrQIpqjHUlOQ8v+W4kGPNiWV0rVd0KVolQDgB45cosiwcw5GcXXtuJQ
676qUEXArBs4VcrUo2X0HldhMMyBs1t4N4V7iLnhRiC3L6284ObFPxk0OkwECpQQ1Is4eWpPwlRQ
GrPbAihneEGLEFgWhS0QnF3aJnFiThLQMxRsI6Pqeeekn0Y8la16jxr25sHGnL0jupUCvYi/ifCO
kBQhHFchchpHs5jERsC3khPTHQycEjkR5L2dPEhbq9iBQygf4rLqOvuXNjI1zi0xhuL3eyjwEhBp
uzipd4QO73bKm4wP22k03x5sFjtSbOI7y3HzT693kSPGp6yXyMYTtr4E+38vYWKqJ1laPAPpVPiV
LNfrBDTtOuKR+SSriK1iw/lcJDgPM+De38EgtTUuLklzmL/RpdnJ15pA+yGzn+hipM8mAyjeGoNS
BDCCMD3uw2XY8nht8wPqainS3uywJU/hghtz2VUJEzhl73Z07l/o5EASkZkm82JaIlHR/yVuXtho
6c7u8qn+9kwA5wNnBXI/u7DzcNSFQzBekkPKmQHi2T3E7/jPoPpComxy1I4P6or9rw1SHRcaaYXx
VfLvHUsrbXMGxyYWNb39JHlbtF8xzEkO4so1GXHQ4FZlF5eybIhj0kGHhjdSk/bgMVDv9WsBwx5s
hQWdZ/C1i8DF3j4pqSZxwmFLT4IQbR4Db1aoh+QG0PUgPDXafxXmuBFQDmek0h4+u43GOqSVUDQd
bYtMxV/kA56IZ7ynimTEOSCfa2d3FnbgIF2ThE8adJIB3Bf8zxG4lSISXtBpAuVKMReTBdT67/3O
r/zbwUs5nQNbo0CE2HtxfU3Zb0bvOxbkgc3uS1fg5YZpt3NnTBoxXF6jN3GXbPLIWA0yHv3MUbwo
ARoa7+ieive55hbODzSKGWwMQklZeGlhxxxrHNeVd0P3Vc+ngUCdZC95glzmf8TgbiWXFREf9Qno
AqNaUl2Chx+qfAcpuqjALW6u498Sni61vmKu1ruwSCVdOg5hy8Cq7ZAG4GcZ4bjTHExCNHSCQM32
yc2HiFLiA0JqL6bYSap7nQ45byONykqyLj4VRQIe/+LEQyLANcqZQzHTdefkAlH2RexW8vyA6vqW
q5hf0SkEzsNh7jDVEx5i9orzAhHAp5xLC5DBJc4RnlN1uk/htFTH65MwVbY6caOep7TyxzNKgM9w
5dYw/sEjfSnBigvtxaoOF6z4PmrRgO4gAGFOx7YkleoiuCcfHRqm1P2S/NbJhUXeA1HKeOOi57ti
R2i2GCe0OHA07n1CJxUNHVyYm7xGXVICnfQivJGypmka9ioWBH6b37EElLesZF0FyLK6aL1IufZ4
DvKgyBNtlduz35wAdLN2B+j0h0nlhFxGH/OfJIGFsKmI8DlaE/9k7ABeX/BgnQ+9cgAWuWxEoNNz
wbKfc3Ut2lZSnI36caHbTRnCs17Jpl4mqYV+t8AVpGI7emip5AhVd6NWes1rXmCyl3Oek96IH7KJ
wwcsWDR5Hx+iTdgMOS9jrc2hi26pgqRKn7vD5pZOZDPDwG7eICs9Mxc2sbhqtK5wpE3hwKB2fNIY
JnK6ooFgwRHvzq9IJBTFhpur3YB05yj5l1RtBpN7bFNabT4S5vGM0iUPA6XWG3DTwgvvuKYNjMou
Kv0DuvjUWBKHWoAA0dr2cZoaOhlexvVarqJ5qRDhcQF1KTh387TRBqUby/KvB02RdMvcyHgbDHzB
W6YAaYa2xqIoogtC1z5X3Oi2eMSb7gv6bWlo2ll1AZ7qqTlnPd66U+JJ2VNirBSaBH3EOhYkbWcY
LYrw84hluTdg3R+iMGnjbErh7Dr0QSD2urcY1SUhh0auhiuCzHLqQWjvcrBSuG6RNbrUkdAnUvr1
uUn8rJaPuimsxOJMs1BBtauzsDjTKinEjkfukhAJJGTI3k7j617fYGXzyqAPHvM1bf+pypD2ohUz
bZDeQeKg8KZWkOVbkyeHS2H0tJAoYjkHU40170T3sE8hhx0KfFIg20aHl5m8f0JP+ElED3vXcuvJ
dAfDD54m/KYw25LFEsZZgp8iePCp57FNyslVa9xh8b1XZQSo/j6km3tUITEFEYpshMqATUs58fvX
30jejJrfeg/AJ3ymZqTLXA+EyTmdm8i1vxHPwEwk6TVrr+o8IkzfLs9G85XopOgpUOvfM4iEV8+O
aqDFacHzeghhsc/hL7nBzQqRGCpI3aI/wFFVKEg604qEFvOl4bEj8cxv0Oq4MDQ0VAvUAJTA+AUe
56gpiPbsPh69fV380ZlC0fqgwPHk6ioeTvuOueXQjeCIkWp3pr0YvPa5lC1t7cm0I/EO14taGHzA
Np1BpYG+p/X2f/V2zMUFfwsPdBZ0/WX93wYP7/PrL3qkTr/YyMf5EEiAtpm25JJnKGlvfdvrJ4ww
wajGaeqrTNmBPU/fIhXAdolPKYKmxuCKQap+jV68jJFH//ARzdoK4ehskf2A6GsI8Pj38KNduiRD
0P+eCbrtb2fxf5w0L3zu2imTGoLMRqfqt15MHRL8tlHaDpcSVb5z+aCTQdh/YjyeHt1CCNhOaHK4
ne2YttTIuh5dI7+goZ3zRremlvKyAiVXlnKnnULnrMREVVmXmVNo2WkS2HQz/UwoGdLpXwZLljAM
ylClUq1Ew/Yv14unZf28fnxl86xiHE+SjXZJGGUJAyUkxiJA3VGuOHC2W+bd2m9vHn976ZaoQQn0
JBgpwZaSqYj7xp2Avf4+scq65Ow815Io1VFxVo+fIWm+rQzCg9YxhSM9/gyg/E94k3wSCU9Wme3z
jPltpfUnUMTB8tOHRyKm2PraERhpeKy910/r5HLHJKTxSNcBcn0Jj1m5ABf4nDmjLJ3/lJvGYwN1
Z0RsWmnDk35z/NPHTOB++qQWJQsbJO2+1tOTpmWOTCpDDknc0JCQGSYl9+g4IaNjVKYu/ZoOXGZc
8q+8iFCOof4yefI7wHMUuOusA+hdag9O5YxXGvCpQArFQzy7P1mcjaCKJPwa3FLlZNW3GYhnbrdh
TbCtse8xPvlQHLjsIEEPxX8iw8SDhykqy/dQ4jsjiXczzYmbcy4y976e7i4Msq66Fq65eL3IoMMJ
75suVehUUHto192scc1TGXNF5dRYdXTd0805IaxsFKHE8EDMNkqGObTGMBubXsYu83Nqg9pT09kq
TM4XZHX87izhppr8iVFyiOL2cm7MGOWH8ObFn4V3rVvU8aIpMbyAGjxmIFaMbXHNUwPCstDA/WT4
zdamdpF38z5Vq9d3PaMEH16P81oGK5+x94azZk1RfzBz5XHecTsrZkVn4hTbCj7YacPXg0Daf2d9
xOK4tcTkEUXdGW4IRhL994YvDtZyY0iuxM1fgFKJJ7EhNoVSNIlA7uNhtfvg2HlKdMfU2RF+m10A
yL+1tvgQxJUa7hNEYk5y+kPF+yi2NYb3RntKg3De8f5Vc1GzxHXuUFgdgNG5Cb3NBzEANLPTn+ch
1qE/XCUKrg4Or16T5HszM5d3pPhOy6XBBsfAABFDD3NLHmdB1tMJSXgFXjDxZGzmXWdinFFRcw0r
wEzunKqyOfTPWRuj4jjKUMmEbktEYPJNZG7ZBkDsp8mFx+SPTGMB5TLbw6kcFA89vRIT5ToAhYA6
WEwiQjq5Ydl0gdUA2//yxlPcsVIX0W0sTZS6DRNAHpCGpWcTcQWB28cVhD8hwxw+MTirKLPFj0Oq
obxhcg5x+IWPeVPUB4yxhDGqU+lhTGyR7X56AnWLtl2csqB5OWvWNrfaceeOt8lBpR83jFsRjYmi
w70u/g9yCwjzt9/RDK6B9Uf02K7fORm1U/p3bSOpcI5+NZ73nAWO3CG9JscZWLn9XGhMub98iIyY
67Tx8XSQlNy/x6CsCJExoa3gYtR3TBYsRzVh+jBbZy1zgij1FMbSGb6BD+zXXGKh3LsozFW1Wu9V
9qr3S3Eo6XfETfWGLDZytkoBSXw3ChM/zyiAxa3ehs7YlTn1gY91ULvdYBaAAwN8cN4YVb6b+5lV
RCifQarMaNj1paorkUL0VEiYf1j7FYTcOp1OfWovyFz80uRT1RgWYHeotVCdzBu6TEs9HB/A1NSp
enzV1zP0dL6ZZgvykag71fwDHKGaute2pYljkLeLRyl7ggnFIL6Gyj7NzHQFdHqXtyeDCHD2oLNY
kyCWFWup8dDNnlKWAS+iz9TIyuJvVErpKrFo7a1Tg+4cardnRqxlERdnMuTE++PiYpEfcNz8UUU1
TsqXZ0QZJtZOgAVT5s0irBUJrfY9rPZO1fSLObcjgD8TUCsz2J8wvSGWh4+2PlLaBsMMUDpoViwZ
bvfoPKVzaEwW/aG1UIe7TL2W5b13/S9uY97qKGgzW64ORz7v7BBcTXjOQgenkgGQJk+MKsyyPQTF
+QDreehUZ3KD//2eWdza0jykXLdzzYPUWOw8uLByX6rXJlsrRd8FKBYyGoVS0SRnC9MSU1XZjOxd
c7o1CCI81FF02/Kftul3zY6DTVvAIlZoukeqAaa5APafuvELpvyz4kzCTTsq0yf4xf5u4ixIcrt0
KP+EvvGfXSgj4VOe1Bd7MiQ7n0ZQyt8yfgevtQ2C5yfIYiClNrebvalJxHphZpueD3JWYWmEnedb
3aRLzauaZbLVYewBp0NERRvzcU5K6t8XTQ3yhjJcOevg656glZoeqOgLyOcp9wWunKnmTP1SXCfG
NDaBV5tA65m8VFizdO9nq5uvbmIYm6S3i/ui0DfMZ0cuycidMFd/52BDNbgEY3ZWRxYc4y09GYr0
iyQFA4hHE2wY771V1RuPwO+0HNRqdmrbrStwwlpinyTGv9MgJ7idVRMnL/q6gq5WVItN+LiWj4vJ
WP7jRESRD5mFQqIe4qa8w3Rh9Ea9AxLuvfHEeHPSMBDfIP69WgDQfXDhkoFrezJK/T1StVJAI/Ga
mf7G1g0YLPTQTCv1DQKsV12ucuFGYbdnW8wSDIoUTDtuFOIzmW0Bq4cpoVH7IoTxksgnD2YGlOAx
6/iz4ceaLUSyK7Bc2Mz90EFopWIEYYPaH9Vt+aYfa87yldUCtB0M4Nt/zqnOJJrniJTlLafwimSk
zleye7q+iRPcc0GZkRB+stOsqWdbBGT4Mvl8nkypnIQgKDcZO040bgdXEgFRBQXOz2SLCD6KK/V/
hnn9qS/WJH0coIxMsw6DG2W+hvLYjTnG8VEZQ/XAN8hWFznYSYvg1I0oV0LUV4NG+w/FzYNS6d4K
XoEvT/W/JRqzc/lPNhuLOao5jiWMFpRBR25w/O3sUBUaizWaTWavvKYiO8mwIcaP/ansDiWsi9HL
uQjUTRtMAlMPHFnedimu8QTxK16gh6WnoorXIH/ltWRKRFsZXI7wnX43fgJLknb6Ys0AYRP8igW/
kZfRY3N1X37Eid8rq/ZcSc25YLhAgmk05+ZfZ288bmCS9IPGcX8p2/T8HfOfv0tMBch6xKy0OT4k
WDjiL8AqtKc13HnLz/Xwo6GiJ+cYTJZ1SpFS0iQsuA86eprCu0WPD3fLrSk60kcp2zpbae9P3t4E
SVuf6GLxfdBcR/SRO+3FQFysKg7cbkWkNuh1+N7XnNg/0+e5xCH2TGK7iXVHeztFrVQY+x6EzdHk
dsLDUSRNr4Lf91ch1Yi2UqNEhzgbkQ8Aedq0Xp7ZOdrOzPlJRJ+VLQSL1BwxUq4S3pR9qGmaXWEu
ingnzVEGei7aIddkWE8A91uHLSISd3hXS8KEC3crU7uQ4yJ6upLXLzZmaxr7izQOmVgeU8C/F93P
xBfhPuqdNrQ66eT+E2Ww2R/XoUhOI2f8/sfznlkYuRdyoCYHFyUT5cKjG2MePRVT65C6/y1559zS
/VupXg75UC4E807U/H4XX7zRodzBliRQvYUJc5liQT38b8WQGKExU2FqSzCJi6qDkkt3bNeS43B0
FJxD3rEbdVUBHGYK5PUjoE6IFXquyLKM4cmw3r3H3Y8KGZRgJGBlRqpqA9PWPsa8CMvaRHlR7htx
gpxVT5mu2A1Y64JVTi7ZR74S+59svr723ohXRkdg18ZKC+fIQDx2tGXwnBuRjxKSsG9RcNd97uDl
bK8W+pYzFljFjeobEcDwebUQ/oGaGasuIBNfSiXOYnxzJ+Y3DpvjSoK6SriwTpqdYIk7MITITYoX
p2ykMxWTDNlVGBZGX9P3kHE/NSo/A/QtbQ8Lvz54pGBQt2MaXt39TYSPnnZ3zL9VDhk8Asjvj8ew
pncN57nwkZGYT6R1XhIefnOJEJ6dXnacdECggKS08Z3rgOK9ZzRXE8KFFAbGYwXRCyTPpRmjP72A
rcEiAiLGXYCoLkZGFnJ2+lwZMybZLT2xms4ihCIdJeCylEYpI6ceevxDimT3TknrMh4lQkX71HEz
m6yTvOQmNv8v3uMuDHimmqFIyYbnzbImYcA5BO/6WNqAYU5zyzmQBgzu2D6uJYIf/bfactw0H1TM
I2qMyED7CU12CPPB/CtW0nLPYx2BJTtw93JEZesWI6RO9Nd5zRwl/dLEi8xBnxwshV3rEYXx/6of
+WIfJZvGClI8Ai1aHXInrtDJZ0TACmL0MA7VBNIudRWBf6jly+Y8Ozt6hgKbuYK0+KDJEA3SNMRM
jQmgBbt7o3SCJKLktFPgtX8iGW7DczNGGejI9PLUsJAU5vmFaw3ezBsMmPBpvxD1SWdiwTvmLE6k
B/+dte9A8hooYqNmlXd1jD/AQlLFOWbuJL9bIi2Qq0BQIJjTHIYk0qNUtj3CGWTandv1cmFCwEUB
ol3Ux3PTZp4XzE2clonPSOF4s/aWkoMxpvzu18Y5BCu1uhbgM4hOKL1JOvH7ZPDVJ9JryjgbeTog
4/8JSerzUig2GpP/9Ys9Fxy+9/F/ltfJTin7br79VPDiEh+ft+AUZMtXWYk6bq/f/4P0mBn/kUE6
DAb9qPR/bYEnAwVnZrITe00OkoXlZhdLRIE+7VP0sdv6vsc5LrYL8KTVX/I28/LMZqsvzmbEUvy7
fCuFCEmQHV9NB4VWo9V8IRCe9SkZjnP6dcworFZcGrzdDstGWfVy04w3/XxaGs5HW5GpPeKlaHOk
OsRzmCTOqJZBoKJRIh/zLRF7XRbR5dbdiGMmLFwgEXI9UtdfnvYx1E2QysDJ1zELoTgMKoGQeqFz
TOyYAT1Hxz3qXxS0vMM2hWrT7XJg1i0PLVWkBxujq6wjEc5K1bAzH10g2MGNxbMmJ+WONIiwFER9
9bFReOFA5ZOjTkv+XpGnu+20koNmDQajff50JILSVeIGOaASHT6KmP+w37ZN6DxJR1O+CicJlFEc
YG1+RWDSeu5euTY3P6wFFBLZEiPBYscEu/WOvtFJg6nqjO8eoqZKLw3OqH6TmuaJ2c3iDyT9XMLJ
gHIXydE4YyN9pzkUvh4ym7roNOMwElqTraQQz6M9byh3PD3n9LMFEbL28S6dt+46eivQlRcgIUJO
kO+FIcVsmxMrTMiFJhWO1icgiqYmojaOrqkiPYY1fRMgg2VljYhm2UgNQin4MMGNHhAx757czLAa
gHQylRdJnpKA016w9qDf/jeu8Dlf78MmLwBWjCRMbgtqVWtXm+gbag9T02TtzL51e7Lp64dgxLsf
WwyjJJgxG1540kUlbNiTmA3lbiCOc2ljBiteUA6G9aRdaLQKqtJ5IkFCVl8HaUJXXy3wtaAV9omN
86+qf9rkmjoT55FzxpLeUTnXMibbLd3bEbnqbhx0mQRua9sJESKlbBA/e49GjTgpu50ujJ/kuND7
E5fKBc1d0HFfpIuBhj9lj9uE4bI7i70oh/hSPtEntIgE8Nfs3KUUuCrBWioc1MC7l3uUOZO/J6wK
kjgD9+zNGhcGhwuQGF3djrbKhU5i5rzAczfmGbklZFO/ppYmB1xWGf0GvJofcSQruPU8x9ZkSG7y
xonY3ODpCQJB/nzSNvR9o3qhd2Wfu1/Qlxm10Gq4Tp5oczUnDa8LJBNn+tHbz86S9tUAuLW7R90G
bHPKYg6JmnbgRr8LmQ7UVsT6yuqqKdE+JXkLaFohjmlk0o/vQpKTl4ILzGYSC0HWjMP+Zxq8FLoe
r8dKQ7TQ71ofaMmxvmbtcWbUu74rCwz5XMPtj659BpIAR2hBDGYPG6AOEY/oJ54rtkS6Vlgt9exA
GcswNgd2a0n0Shoyr1VqtUjpTd629Lr7fqqyIfQjWeWC8rZaTIeEZVQcvEGfr08olPAJ5rwhWn5k
rM3PygpS85BQzyhiqUzuI7v7hyQ0xtUJkZQrvxse5EBhRfYwvcR0ts5CocDB7QczZ7vdNH2f6BRc
jx3f1TiF6l3Rw3sVWueL1hamhxZhHoKEwMi/oehPOgYDI4lN8+fU8em6HPJDNulWYFYJsnRhRNGn
JUJmICaDiTS1oiVsz0eWrdgbubXo/64tyTQHcWXH+WaLPzQQ4d9xy6f6OwiIQ0V/TzpfYoRDvK39
uD9ARi+vr3smPrXnDH4R8J/mr/LA1OC+YbLObv1EqdDN36UWYx4pc8XQC9RwBQ4HZ4Kl9ljn3p7u
RosGTFhOeEQms5FcdKoEYNqMaEudivFMEEkXySG3skTLQ8yvvq9Cm5hsWt000ksDDi+c+q/hJgnk
dft+p0wFmvFAv4kjVYswcCGNICp09Zbeo+lxcz48wju6NevjEBZLbyoK/okc0rMNg7rzRC4EVxi0
28rAFk/Fs3PURDuNP24PqL7k5JOwQ+kCQjWmGgAl0QvrJ77LmcDIe21yIyOpY+wyutzd/Lum7jrL
53l1u2BqkwSRyuYLhE+99Ht5CVYGR3vZFSDU0zMsfqNMe7FF+Hc3Jn5Fcd48OIz+cgvbikscw7Py
IrEBcEOb0YpXs3o9x/pZauYsc78UyNXedDIbM5Z8ramuw8yaykIS8mafwT7BDhG84ik7LTgH/Ior
3iEpYGzmge5usy/6+LQ4kHL1T8rVhVBY0CYHvNRuY6n1T6aVuGGiCEbEWMPBaU6int/bbpF8ildq
GwHIeVmZEKx/NI0/zFgE/rBMzASwWfgsNWx/uadKbtOW5NAiwkDQoBjhFgRluM4grMw4LynMK4W3
kVvOkMSPoGOcq3qp+3wue1cqURVsRcp+boA2E3whBObswHjC8qf9QYMWGPN/umoUDb057Fox3nWh
WiWlaqc/zW28rwn1rkYz9WmIqsAgzP2CebwnygfdIb7CK75Gy446EgRvssuzlIpmdRUiAu3gFVs7
He5GUr9FieGLGJwdCSfusfclRQH3dMX3t/08Gy6Lf7kwQyN8t7IO6GAN5V3PgQQNkJyY3qyaOtrp
GHd5BJ8vUl92jbK4Volo6dbVbxd1/C5fPIIHniaY+ujkfNcchgRxM2nhURNoGK4vxrKBib9Xug14
3bZwL7qsuZqHEQuqTq3/pqYUFP04CuIY9blmQpAEKQ75zCBw1sxHI5jO4FpTDCr0CgMnUoy88mvV
8I8e3VrW5Ru7CQLPagNpHm2M/RFb+/O+7TNzLighM0Fa3B05IB9IlvBefQ9oQsO/Ojkq/3eBkU+U
mw2P3OV/4TckkeI+CeaQ+5Z3DPIidqOws3072r3Wy/5g7W1Ul34ppXZ3VKpOP1uFxp27O8xRyK1t
YNm0qwkdDN9HT8h8ZjAFDTe1fswYBxN4W1Y7ovDO6NHj3ioYu94U/v7JjS3TqdD/NnKnCvGQSg8A
hRfNjgEM7BFa1OHwP7kAbERydKb86/8S9stzZSPOj+e5o8V3tKef/ZD3qwmDDMCKmlI7jU+uegUG
6gp5hgI+KaMoY3tNb3QOKG0fKyuQTmhsMqCUICn5THQrNTCKJB06L7xzVGj/f7d0W7GysK8KbIgA
E4xEyzBKQG/kdECYcTvVpBIfIlbCnJxokzAXahsfqCxvhM+rJmxoEiK6A2zIfM9M4AsbWXFIbjCC
4T/TQgglEwf6aROtkQXXZG3MtH5QJX8thL5jS5B39EZIwpKb8jNTbhERBUVM5C3cm7ClBJMKOe2G
hI1nNXBlMO0F/RzJp8B/xQ/VCnyvNwwUXE8Snvju0BG0UvKsKXJ71r56cHdPtQzJjSWh0TIpG/54
5RT0cVTB172W+1ZlWOeLSrtl1vkSbxMb828TPyrgwro2W7hS43PWzneShe+cRdkbW80+hYJBIiD7
LJ3guura2YdrEEXI+Rs2i/4R+3mL4e5iV7rXLc0/g0M38d7CIcgsDdc1pV4s6lCF3wDirpccgHiC
ws1UfPHMJd2kQcST++5g+MfHcJDVsfF3nWOhIe2+SF0/W82CzyyucJfM9ZtVzOCh6dH8rt1aWrFG
CriA6qhmKb5n3PO+yrLJBNleP/J4SL51bSfhDNxjPf4frJghU6nVwskATU+DCQqDhoCLm6DOUltJ
G75eAao67UrcslJ2SFluWm1NiFoZS4YOL7flV6KGBYPGtGZ23QbJgofJQCeKztmhNQ7SpqrEUuV5
PbncZcDgKnDNvhxxquOpBZwACSxnSRn8E/3KwytQ0Z/Y8BoW5Wqqf6aFvrmeXEe+1jsEQFS/z/CO
rcx97CrUMhvVoB0Idh10lHjFJXpElVtTuz1GPI6JJD1cCtMc2RkDabuhbUU8cRZFhPzl5/iNXcxi
rvSGOz6OcIBabega+Sm528kxvS9IVrrpZlUIa70eY6AdMnkIXplGSbu2s1FeX6gt7l1AKRAFtI8b
PXKbQUQGbSdUkLZY/8DV67AMaTdL7r3SmHiaebjGxIsGi3ar8S0qfYjhy1tgmaLGBKklgVcaH5Wi
OPT+GOnQg0WDzWu/TsxvFP1QLQ2w6ilLyVYiDoGAOM8gTvNNWtNdtbgPfo+aOf7hbfjColtqDXFa
4TWHh0dFjdui9R2XHFIg/xWKxJFPE2VIIjSquuAVfQbUnUbiG9UO1dl7WX1KuGmqOWMtBPPxh+aG
WwqY52n59iAe5+8nzmr2+TBzCNwLTftakknVGIflAUrqTtLAfw0zlDw0VjxYST5MzbrC67C9GKI5
PpBUngYMYYkodC/2jsfGACDTwElrHbG9y7Dh9fwjJpxnd6Y45OD6NcKrqUtfSLHkm+ah4OXZSPiN
z6nyEHffX37axtOAmkUIUv3R2OdWBGh2QHLbDZSuzfDpw/1WYSR1aicON/hW6l5FOcRKnhf7+pBV
/17iaQMypAZtJUywF7jGosOqlY4bpAyaoo3YC+sY4AtlCXDo1g4CxD6+hAR42wZE0D/Nsk1wWtFY
/urAfY8Fr+taq/+72EbP5y4ymFODsZTBsQsI6iqMsclWADVhjUDkx+UxfEPQyqQMrjgQvogSAbIh
tCYu5uied6R3cK+/ZsoF5usXiuoO5sNH1o/ciiQ7u6/l31kqdKs/j4eFy/NFMdWjciUaP7Rwh64t
LFuwhKPqHJOqD+nMj7AwJV+6Xh4fqa5xljvXuUI7lkrdKCKkkNwX/vAcjI96WNAAOhODelMf0UEP
/Imnm0CHzgUD1YloASjx9oCoRRzDf7aeumPmb1F4UFGtjWBJIzkL1eL3ToAMCO98X6r29D4K+loM
kfcYrOamjv9V0shJGV69sfFnhrgkK+eq0cTKiYikZrEwmoqJ5seXiOM/HD/UxzfSXCCugsB5trPn
/GiQgTAXj+pV5JAqkqd7mkQjAeFuKl0TGvvVgES2TSPCRXWHQ9dxWwK4eJXuORAcOahIM/l1I8Qw
yBdqFmn7R1uvTsTEUvlkZUv2HcdiQnDHmtPHWSSPl8mxQQT2qceAZL+n6oDG+8ylrqdNIhGvSYzz
lYZ2ycGaqGLsMWqzhx3E0dcY863g7iuBIrG2aw6TQ73mPArJq7HqqoEG6eFnAYtM4DG45jJEkyJG
sjxeAZv0p1ZoCWNqBZqU58YNt26O7esmk9Pcq2lyV6UNCZp5eE2o2WgdsJsQvPF0kAktM2CowiAf
+6CAxssuXf3XlXL/xtAAEPigjKteD0vJwEDtUhu63X9WqIfWyl2d4jd2zoa1sPy+hbYtOgvFwvqg
64eV10pHDGL20CbWQ43sDk6Fi5g/qSADXCiDOooCvRbbYRSGTxUW3a9dEPtoZMFl43dkN4tsCIaF
c3lFQnUYcmW3gN/iDF/3BEo4Go2qgCsHduKGJHmpfCYR5WS6GLkskzO3Y3/OOk14GWJ54BmfLxDu
olTyG2+hrR8KmQbECNoocAFROIwotbPUSDKl0KiSFH4Ris4h8ViCZzYWnTKlJm/YtP83ETPo2HeN
DzRHRDPRdLtUafe1duwztfbbFZSbPK/lFlYqClxmqlQM5RPT8tELYfpdUbAac5BQ+W+VcXKUb/yf
MfaI0n/QMlEr6CVj3dXrr1lz+Hh27zYCI79E4Pw8j8lDBQ1lxmI6aA6Q10XCvX+4LwkqWDZjaNpL
Ndilh6OtdnqWImu6Jj+Nento5ezDvx6Q1E/XXJB5943Bo5bz768sW6/buydPuIPQkd2HLEcUNI4P
wpS3ChcKjMk9CXkeTAW6WF7wnhoSmlj2ehtXXxtwVchS5CHPZkmHs0/bLW1DZkDF0xq5SeGJ6ZmK
zXEdvMYtStrIZEI3PfhmIYtxskkZKV1800RJfFlcIbDl+aSm0QFQeOi3eBQ2fIpkFDojcY7ssgRt
wQESms2Ug/GNGHCiyef8x9GVlGuWI+r8tfldOGVfkcmx9J9i4uOawe6lQY9PBAdyTnnZmTY1X+wK
jBKDQfemluntUYOie4ycLe+8Z7fZqzVa6AVDqA+dYDWqW9SMHVLIrNLNfU/VCVL+AZWF8tKypUTS
JAWmS6U8MfxnOJe+b0wFGubow5RM8GUYx9dfnjQbXC4YkZD7amEhWZ2or+NOXT0l+mZXX9yNsN4S
9fs8csfSkHDvdMrw7QdjdHeBqFizz6DPaCSdA/S0Ub47Kl/Ughd1ZjzwjNTwjTXXqx+VQ8OySX2F
hdSFGlnb9RwWRINh6deTWybUy12dkAEPDawkxQGo1BeEKcjuWQuoxwbFfwpkTUVHbYuGGBokexuj
fef6uhiX2SPHLOoBNw3uvvr8wwL/K50Qzhmr/DZ2Gm/Q+lW6lU+/BhRXaofbjA1UGfTzDEhPh2le
GpUayiau/K35hdIgvjOkJptwvXzBawdck2k92rJw5IvhPvoNrAb3r0faNYfH7Gidfstn/35cTVuv
wlHzSdVzqXxlcnN8tgITB7FLdNu9Zz67FMgxFKmucxlFTIHAZXOjVifMqTPbM2UAkij80e/EIoHl
FmlJFrXhoJAl4jdN0v9lupJt5Ew6qCuSqN1nVfm46jOW4E4xS1fRPLebq5Q58rPO4TvwQeXnxjVm
jVrCBbZ1R+d901YuznFa94eIgK++JS434H2XYE3shoJzDGxvjb8DBGC0DUUa2LUtFq2O09LtVW9y
dgVVaOBFTiI71K4sKoDBhBDWGxeILhNjOyYogPHMfeE8c2FeNSqtdgHEExNNcTiw2zvVUQxikcrV
DKqWyoII6Jgdu472RyGZ2AdLkwnQHg/RDhZxAch2Z34nIy94LpGCyNgsttWTNSCtWKd9fuGG9Vn9
PIx4Mijy1OAsRSpU+Yu4LTnR64FAep2enu49iu4rbLv86A0Au4GsPoax6YHSB4Qtz5df0YqckQbV
t0z3rxMJVlvwiONFSzzPtZ0uXyz0W7mNg7rL0OoAqzqptF37OtVwSzX/Qh6Q15yud7b0CD3sf/LX
FOOQSZ/UNOLzOvTKPYdIKPRljPjzxDV69ptZrrjKkqZO0MDCokja+tbB4Z2AIPjyAE6h/iANJwzT
NrDwElq3fCs6xSw0itPsMkT5Tava2xg6tcpuQ2HVNr8m9jkMXr/LqS8/glzbvlnE/f9PEdDDHc4G
/H5QoL9Q4hN9IBn765usSmvUKeQEthV1TkmgdHU8enl+cqQF8zMhjJSKOPFGCMyIaoGpJcSlRynH
9GFUcsCNmE1W/VhmMKsc5vSTefPSRlxqQMKBq9cRah2HGfas6TFhaEiebU9I2t+OCv5x6jlYTjgu
DbPwuY8bFsuYPksXfkY5vlTvMgh6lF3d4d7ryyDqZl/HIGeRUxuzbeJ3MB3BhT+38CjvzSm9gpr9
6vdSZzU7VBy0NYFry6tdl4AqjIl2eskW51ADwnBJIXTrP3beTC5mfvpmSErpew65+cIyWx4D8E1A
ek53OCX3a23JX8QDCqteLXG9gETuIAbKoZGBuvGELq7rmepWoYbvI7lZuB4XVYSvys/zVjgZkeKc
jN9+gH8EbTpgKEVMW8V+7ugDZGHEi4xcfXGFUhgqJKTLZRwzcoITweAz6ExvAflPxQtQSUnCUv73
IqN/GNahfJXi0SqAfCGtL0NYMzfxI9M05+fPLtMq3lTKumslDJZZNc480ZnzkwBMdxBhmZ5FH0mH
U5dlA5OTGO6LGffVNPDgGuhm2k9d8wQ7PlPK0/X9lZjbUBvua3+5S0HnEtg1BlLTUx1i12tKJylv
8Y1Sd8FNrBVFoV4oqQH7BwNHTUANFNrIWfda5b/++SsLC5vt6IiteXM/I/GuAF7qIsipFtCaKTG/
31ASclfBwPxN0NkNvYsulO6wu1NpY/7iI5KAHP/g4wv8gn2A0JFIwofYKu679IpXEsN4cSsx6eAv
tMblm6L5UoSJBCt3AUSc1cVVi9UjqIDCGAJ7psoOZrkhOHnNaqXjkrLMq1YJz+51RtrFUSrF0hVG
btFMGFbJshX0S5Vj/JdgJdGsrW51BVHKaYf/TZkQa2sDf8mrhpx2QORBgd1vpmM5HEM9xsl6SpIJ
RP99UPeucmkC4OflamA6pMLrwdO0gGDjKeTTWnUk/qQPG98fBpXGkzCjD/ojr7mfhbmxQPALPnxv
twnTyNQ9HtQ5yjO4rOuyPpYlG6rksBoHvDqCdkZBTnDDTY2E0tBBstD8H6bTXmyyNUD7T1l7OWBM
9G/fe3P7Dwqri8Tvs9DxMJRVxK+2is8rtQdKXi6MqC2NT3IEb1L2q3xlqinAJgQC2NjDhvphDmc0
h4PjQ4RqgQGop7H8TcCblt0EEEeBbUVw5VtTyz83U8fx9SIYu5JQu+e/Dl9oBUntQdcqPvM+LLad
4xnFE/pzhi0pzJGaAsNws/+XIrPz1mCHZBFk7XzfJC7ndY9lLSAypbsJoeVe8CASBYcYFDqLLLi3
kMr1owvNUohU0Uai6Gy0vSFOZf1K1Ew54trvOdDh1ZAoSSf70uctbEbSOqySPpoobTKuGuVCg+b3
h2QO8ii/pCv4Vc5gZ3X3sS7ALLenEtxn7MAutfyPD18Ano0KPWZFatv5x9U4yVr80ruYuBpZn0lJ
5vEWH4cKAjXXxlLMzxDQj/pyL00ut0OUOeUln4VYCpf04E4ebJcF0UXP3ZxnzrdmpuPrQlxWAfuf
qv8rH0IFs7GcsxKZRRDcoUBb1kGi/+ebf8svCcaP8q3lWDCmGiC2Y+fEaeOG9dM4nMIVFkjXOVex
PnH1N4o0CS9HE0dRHHq1olD3OjmmUdyYILLRVZ08yLlXatMpDtDmY1LX1kZeJm0jflq4/s2shyCp
USg5OkKHkABxu15KkyEmfM+zdVTo0GCZhdSY3g12Tcp9zry+JrVPkA8EjOGDxrBW3IfAIN5Loi4s
jRDVaGDsDD86BsT816KajqpnmJfC8vtwYQnvt+GYsP1OznMZgTkkYg8Dn8m4Rr1KkS2HlMzXdWoE
buKE9Moi2dfXQKBi4tdks4r1y5Aot9k9QS/h2VK73eTZmFwJryCU0AY3CQR8zQh8Fmf+Ib/UKzi+
8Ihxexau90lGGwKjl/aNgRtGHbxuyKXkKr9ts80iHpRfDVeXyu8CF9djFGEK8EAC3V300FB+Pe5B
qWfXEc3x393rTBBvrN8AsGQkKX0GnT+n4TQ6IksUYOC/xwdKGOoo+R1MjHb3stb1jMK0OlDEXp9a
8osu8Ru0hD3RV3R8Jhule9MWWilWAG0rIthNEKoR8k+IhsL/VBoERaUGZUwVXIP3XAjJSAzEWrPL
PCluN8E9fPBM3yqrLpTIsFLbcwKsQg47ztIdcdXmeqTvoIjsEBFQg5rNurk7uEQl3+4zWD0EEJ0z
sw1j3nDdO8ydoZfiNrCYbnBBSLojCZod4/cAf3F99VlipTc4tUb8eAS9d7USzIJb/hcfs0WsrIRf
qZYy5VbaNhzU/4r2zRQZpUGFIhgsXosFEaPzVppghJwd0zfkXIpckRJLW1W9ZZY/8UuMfcRAQS7k
OkGG1YcDYM0DQN2qjiiMLiqH/QR2ILWbtpk2BGectGULVC6QtJIQbZjmGlqyWmt/5NxCJdwh1Bo4
ibWKaPhaR16SjcAPsM/IX0sH8QF5s6RitTwTKPMsGwy3MTfiN7oY6T+ff3r4pwCRrNkovoSNU5I2
JE+Z40tkTkx5wYNbcoMPnaDyGc12iHGJKFzSXMzvJ8FaBzHfjK39nANe7W1DMsxhkm1Xw/VrYmYH
md2S/200KgjrVFZvVhPLP2gt0bat0a5P9R4A5TnklnFTE7QMMKJHrADBd+PrAh0bjChyfkL0bU6a
P+3ya5x5gDpA5bVc7bJ8Xbl2PD+xsrrodi/yZyAhq1aW98ZFZy681VX6iQZDL5dWWHaR5+P2WNJE
iMzLt578vzc/XTkpN3OOEg0h3wApZeHA6YYq6SP67IoEe0sjEmOkBkhMk1MUXv1kVNWujOgmZ/qY
MFUpIBpQevIQGrmeeHxlYA5gnjwF4ZnrKc3gMXSFkhdLHlBtVuZt2Hy/VFdb8FoVkwppDR9tkKQw
1GgO/r+X8c2+D+ZL70zcM9ED6V7GYtsC//gRNDa+y/ZjW1YE96nrLXyjnGk13eIa6C+3jrqi3hWT
tdarl4HdJUty4QsbMj3XywZPlD+1PHzYuHkRnBa4PEnAe3QBwnA7CZbUpBl8HBfc3ox2u9Ak8eye
Jtpl9/sp+3KUNjad7cxKKTRZR1sWPp3jYZI4j/4vrflodYhBCjhZQ8MMFSe/EdyA+te+dWUg7Fsb
X6qAc+1m6vjTzk1HLu9breTjjNgV79TredGRdBCc5pAIbcqiqJFHMYnLSAQVt2X2QgoOnITiCxDX
S+PK5PMZKtmdB/JaeuYr5yC10c9PYMqYsOwP/vSy2EAG9Sts6aWW+8aJ4yZMgKXiLJEWEHFxpcDK
Z7dQB26oTGtYySU1dHyFNNlwkpztNe2cmqnvtC5nxBEqlshGLtONFVp0emKRmTl4xVD9nmtyVW/Q
HRkrsboskDmScn5cml93YqQcxCCSIyvmwbE4Hcu14V00e10on+78Vq2lSZoMz29TyQIAyknQowOJ
j+N0SImQfH2s+QoFdpFDGr1XVZ11qCH21VeA/4n0yxJC3aCB0R2bFMjMbSf83TBqWYczeFjsBWJ7
y7+2eCOa+BDDWchMWLriEIjMhpeF+R0nEfNVtpqxsj0csVnRkE3sh0Gzlz9Z6jWUDwHt3HX/hqR0
ul98ehZrcsyH9TiWjzCYW5o11SWp+G2code31Z/NS8A6GPq8R8cP2snOz5u3ERQ4ylha82xK7GhN
0xyQqf9xBoLkhPTLmRRaIUS8qZV3E2OkKQOTG42usLexHabtS6kD61yZ4qJNrmhYW2BjKESVGdTV
g+Es70I7Wlf1sbdtl8jWdpW0bNX04bMKBBYAcvV04VkzizfhhOCMKWtq2TuyQVRPnp5V4dOJNlUA
zuazFFxQtHvIyxTSUfX+Uvxtbhn/QCNQ7eVCCONDDAgj1E23Z0K23i4G5HN4ggQoPFgB7rxHBLFL
9LkR1aCdhmWioxsJlzO27NELyWkjSNlvG8Kx6KiHC3xD0BYwXVoeY1IuNMNKCOFpJI0QNT3CqY34
PA53wSdUNQI4poqEQ4I9vGCEXMm8ecHiGLP2E19JT5Iwp4eL3o/C6kULU+oEVATVDVmbgYlXpCtU
9YLseWbPi9UY2sdLFs0IoNof25Fqhvc9WFunfB3ketm8o0JoQBjeL1Uzeg+/ZfqSRBWlTR8uusWh
Dvf5QArUMhAFQJzd08RMUIrLAI4wWZdmtTXyJDRRaafGxavEcURS9nDLnzM+DP89SoSGKyKjMWlE
9JFL+XEkPO2NFXHu/vzEc4o1kFb1mtuYvE09ify7nPr/dFjno4oHc6esp77IJ7fF0TM5fqYlQyrD
zZK1mLlpxQF7U7hKUpOou6XRSajrNGqSOpLVOJJdOHsgfUZjVfnV0NxiUOlZZo1LlBuFLykAxhRL
B5bDhyQHxeeMOSSAPYSMx9AXSGytgYl3bmvF/nYC9wfyCBopEQuztRfnjfW1XgfUxTQc9fRUuBJk
0fy18HuiftzuYNxHBo4hfVm3L/sWsWP8xK8nBJsVRq3bGi4Bs2sm8dQKvB37K3rplWYc0MI8C8Ka
glYizk2g4FjSrpDWFYjr+XGFiaxP+FYf98Gm/Pv7MNsNLeWOC/q+31zgi2Imp9opAOP9HSz4rFjB
cX9vxdt9Uxo10kqD+R36ebSU51t9kC3k57JD4VMHm+ilkst0Hxp8ggAk0lrmhPIPTkAhPmzCoCPH
ZywpBiudDg1ugiy9YjbM0qbK1QhpgdAH/Ux9rJnup/UF1nmTpH/sM7itFRbfHo1GMcfWnq/fGGDV
D/pBjNDeTtcQWPmPvy9gsNrlMsJJLyo5UnlCxF7e/zT46MMvx0aRTKzNlSuKLl6mznVxPHekCxhV
+OllY26kOxRaZpWKptE9Qa59D5DZzKyJtpC8KcgEL0QrXUbTfFtEa/5dPI4q+j8Xpwrv9U27V7gu
F1JWzRVXra2KNnLClSSRxoh17zieRJFoPckKcQbeHaxMEOdJJ/JgPCKR3imKRJZkrQY2vGYjJRCy
8f5iJ/lFo8dzl03O9v5ZlwJ3o9pZHgNw3T9x2R6VY+lFEazadHj0UdWfWezqpdpA9y+fyq6sK4AC
4V64vE+TZScTjo6QsQYeXuZOnI2aA5j2awcymHqIgfIpWb2ffu4G2u9bY0xLzhCUwXrtlVbC9LPR
KiUX3KV1K8unmJ7ZunJgSCNPz/C/QVdAwPx+OMUa0M2FUaCYavUHpRT9SAZUJIRztGLyqy29ucqV
pltXbwSpB0IAAR5pZMuTUmN7G5hk9Bj+ZzylDnKMwTX6yHtgyJ12pTn6YZIlt5+cZ02Tf94n+JKs
TKFYPIuZD7d5tIwrhe1WWPuHNppHWUWt2DaNX1E/nUnPvnzwY/WNmr+loCNd892AMOXU0h64rrLg
zCDwm2N42dc0Y3t3hlcepjMX8eCeYLO4HcVo0Ti1rFCbtM9Mtt4VBofTdXfLI3DrOPtUPm/zM18t
Ysjwg2WUR6aJgyS0W/1NT/yEFEEft9graXdUqM0+8IuDD15mlDNdVQtjecSKZaW0vu2TVJTuqd+J
JqXTPwMNpPinqbSqCgwyS/pwJFb/h8+5tLMIMcYZC1lPTweWA5nvM2Ru7ijR+Gmusykm9hqNKfRS
x6zati7rgJvT+KG5fWVBR5etQ6WbTPFvlNED7fQNzOl7seSK3FzEZixmO+Jc9bWM4TKyGk7P6xyH
0Ly+s+/yw2d89S6SZDEW7kOMm9lS2h6Kr7hXas+JLSO9qaiu8p8SFTv5JW+4ZkOQ4tAlJIjjEBf2
ku66kPPRTHx4IuHcS/QV06rcC/4dmY9huU3vWP67wnKNHMNu5YEHZ5xWj+3+W+n0omDt4ssfIsXU
wJzPfk7OdySgkXEV2P+moJj7RobcgJeNJ716KBeRZqaWdSJe10cq3cx5IhJsECdG/BCviD61FSpG
69VwrVHI1By1eLQVqWHzyb7dp7QfpD5hB+JN9mZ1iD/hj8b8JAqt0CAmHzmcCaH+0IuaVGWT7RUL
MzI8ckD8969j1GYUft4ykNVb1qh73g8ZwmbLtC2mnPEmqMVp1ZQYqyECmWDSh6jyBYlS4KMTJE2L
xbG3sqO16jrajCTVBMfgGg3Wkex54raY7dxC1WzKHudwSFHT2UOxTanzB5eUU0YpOkd19/57KUBZ
q5Z/kOLo80FgfKxfpv7a/9Ww7yjcNFNAGB6Rdh4n9XpN6iIzr9hyin3ItZDntNV7zwU1A4xCJ8CU
mP5OQdhZrN4s3/mZcUHX3xvH0g0Mn0ODX68cQvkK5TxeQUsPj56Z2MOAWEMGoB14PKL0CSRpTvi+
YnpTdrvo8+QQ97xcHl1442pCat8ZyxxMCHmHZumC6rhmbHZSTPiyZ6mBzFoCgmyVHBydoT6BCfuK
oiYm60/X3DHR9AgGtX95TIrKibPmKxxaJZ/lbftCjlpAYn6VXbbw+oM4RicYqFnTGqKWtrU5CPQU
aLnOBn747hWwCNwCza8SMDfT9yPJpGIkFJHy9pgZD8Fdm48nyRbJElfzQPOoD/KZci4sz8AVII5R
dPuZp4ZWs5m8DTDj2/JlN8ZeHxOvh71JzKxU90JbVPIqSWi8srkDrfs2yfZ0qAVeAJf+rhT1qkLB
L8MQ67WF8KOhvgFihadpMqud/0ZPCot6ysGvmFmtVnS5Ms9vsuk4u8dDN/YNvO15oBqDFvvgVj0/
7g0a9K0B7ZOD+1hCKk1Ni2gcZrO8z7aL0ghhipe1fPRhisvmD2F/mzQDRYJHtXS9gSpAmMKBkk0w
4MXriwaoMl2eCDyWBh7fiGLvSGXRX2ZC//xNFAcQWVMS2aSRJYIQWy8H7+BBakL2HSFioBzVxA82
FpupzhPL+HPPjYWm9HnsN9MYl3tNkxO7TURmLww2A/udmX4AYloAaP3s1IGlldDVzxyY79t2p2ZS
uN/q2kWnGPQ3tL1CdUOHxX+JTuGQhmIzloC2rWmtzaqt2kDzcxVWO1Ep3wPm6HNmBZMcvs7Jx1iL
T35CKBA/VMuBGYakxcoevEsJaufgkZgfqlt6jbi5w4lrZlOqvCxbcPk5R+/PzwCjzq8f6IH50Qo7
OoQviSJIYjcz4zRTRSDCSxTtPFpcNi/dDhsbL/J1UoM3pZe0gJKHji6slJngXIlGYMy5Znnar7VW
EEPHPF2MeiQ1ZcDt8wLbyPrvGSGJpyDzmI4w6xFcAVovmPmwXfAWyp44NCHeekRe1XKdJ7dbU2n7
6pyKJuowVKhx6iOZDutATl7tl1+4HY8H+AewUgfdTn/eZrQtuS96+gCn7DbN/9nWPtCs/QxB/Mtd
0uFnZ4BHjZVTDWwkppCYLSJa6Lu23Fp3z9e6ZCGPONk/NQ0GR1K7Hc/B+v8G5SfJiw/x4hDYlp7d
hyQHJYQTqOuZhdBoLVNsNYQ+ag7xRhJotVX3oV1zhzmnKYTgaXMuulbN5M8V7Ovgxq2azGaLCQdu
qrrouiytd4mvqXkVNm4UoZ4tbPsMHJ0YdIiEkdCJo1l3elRmFu1k7tcWDUNpx12x/1KBkxGqwuha
HuG9WdzSuNYLtQEvxgh/hQf78JGLjl+W+FYJSE/nfar0xKT2bQ3RAQLt2IHK2h7mnm68EZiuUI85
Si+3uml5xICZPrgZ3AZ5zhNTJiiLVnfHmFJvjLDerIL1aFljEyDmmvUlzNR4yTK/IETh9xKY1jlp
7n32ZXDcAoT4+cwviCNc+lpWKwr7wojQwycPClmEoip0wxkszgHkisKDDVTZTm8kB9R3b9VFnrNZ
Fj22nlc86sDPovM7LFvOh2sm9jXVCu/zfaqk7D1wRCcfN7H4ou//4hasAl1t8NhnM0vbG6IlrjyD
E+AthmEi+rAyreTkXpFtLZSS0QkdOZWsnHUEts4Ka3q0IKo52oz2pJo4HxyHNHu0Pv2r6um1+T14
+msajEwl98GAq7/pIJ2FOnPM5DFuQB5mcT8hBcy2uRY8A4rF9vPG2hz0OkZ+UVnABQMzek3mzOOG
Vf5XlYW8XIEBcO0FbJGBmXfaW+8sBmMorWIrBptrvaNIjkacEcN5Cfzh1zcIrzipg3/F707rsSyO
jTi/HBFbL+YuWbi7ocHfb8Ov2PV3nKNNj1MrsZNSmYIyg5xkrMvq/luMW/Vm8Oqry0LywY+ax+wP
uGP1klRgCCEwPfJP4RpnDQVdZj+iuuNyoGitqXUL01/+A+e+8dfdeeym8QFeYT+ZYrsaz3jsGOnh
HR2hDblwtJ+OTFDWmeu559T44hXadTp86kRvS/UIm29tVwLFid660UUasQkW61et0YEnhAPZN9te
VLDvSsGFhmeUiCjIFEi4VP+xDQrLIzJsEddl/In0N/1YaOUZ8ccQtl+6JmCXq7V6yYXg9R5iFeQv
pmN04JTSlJMx3Xsy3yalVeJK76yuSJBOoj5HwITUzFJeOts0uM1b4ltAXTr6T6f8f+EJERT8XWAu
9Dt03pWtBFiGErWEZ72gHuUEadcE8A4A1Ku2h/NDitfXm+dT+rtm5KviVIBZaxe+LIwnI4T1QZhf
2hoUCEiwOxEzgpc6h68og4Nms//LDVse6/YgCM2BPiDNkFcPbsbZCVn5X6Tv+QNCgDAhnhYNNp6O
WrvjH3h91UGBXYMknKGNOnxkRLLQ6Dp207lK6PR3VyHxWBDhi5cNzzm8qiuWHC6MyL4YH5MfJgMA
uSutH80/Z2J9WHte2NfwyUkuN3QY0kQqVQIvBsEfmpApDcf0eStKQCEcQVkFtIfJtg3ZBcee1Y6r
GPd0JgSA0uPNIwWSQIymZkzE3roScvAWUIxGPqCTyZac8SN5ZB7k4icUe/z+8feaPi67HONh7/7q
d+O7w2TuYN5goj2dVSIQs3OWkA/VcfDyisCgp3l6Nqg3+cZYgOMaEcwiDLv3jMi6ySEr2a1GCAvU
6Yi2q4hjSJGzHkpGXC2mVd1EAVND5UOGEUMSjYOue3idg5K+PYKA4OauCrTG2k2mqrzTsHd2pBcP
kKpuyUnRnJ69gqn1VWAZPMgaxMg/TcsU0h2r6mruoWoED2sTFA8c7bBEm/MRT4YvpJMq2U42es6x
DPtnQQ5pLlzomrTzwxV+zoE9YeO8KRP8l7oxryWtbpXkmnQ+p3kGKUHoID8rKo5PKPoINzqiaVra
yiLFo9BTZfbDtbD+cGqkzBEozIJ/ICiCBp/48hxkbmpgTUU0CN6yVTvm+nFKw6dnJYmb6KTk1ZMW
/vstX4ZmXrOCGSX/uMVE8MTUXR0o5EmZHXbmIekKmQT9ilR4P7prkTMr/MODf5hR8kw72EhjRfUT
L5q8ryr1YxsrSFqgNjYyhRhkwhLOkSmLZKv/FRS/ylH6W+Wd5GF01hZL7qpSo+JK3vHJYwAQTyMJ
brkmBZm9XAzkaB/VKsDpDYN8zFD4FuUX7Mb5F6VqMjQBdof4qiwqxcXaMRCzljJcktAxUV4IZW3t
b2y+tuOrPDUG2mBwIIQvD2nMl1rySYpmVgxrkfX0T2kn5FJgot1yLTPwqJXMdZIK5MxWn7Pdgas6
xc6khJIhNnc7HxsK59ak2wE8Ytv37gCAkA0k8JFeCo75OPj4CJVSgAcpXXLw3qMDi4kdAMHrHR66
GxD79p/4U4dwdpv8or01VuiS/VAEpkwOs5Q5jl8retQFKm2VSLEBAq8uBnDeOa1Q2pup7vY2dfEK
MQr8Ti0kaegwO1ShFffnemhm+SonpoFgW+9B6wkh0X1gVCJXXvxFblCrydRCOWvbN7vdilD1NFCy
aNcxLLrPgXWAGHHBAUFgidFc/czXoJnp8+Djn52I6h4s4VLap/z18+5sb9dMUTPd98YEMQlSWHEz
BTNqSVRtfpNAFgIxTPjpVSTxrTX0lfjcgClWzKnVJgEk0m2lzDY9pZpwVd6YxgYwVUvtiZEv4jil
bFPyLV3fN251WVUV3rbgyUea3ijHpOCdVEkp+U75gb51mafO3R4yqfSrXX6EGqQWF/GmUxLG3oVj
HYt6Dfpg/g/UYqjAjuUdknSuojz9fjWw8I1wOvukxFLvOvfUsTz7ONr4DmMe4YsP4rq2MDM19Qx/
RA9WhCTYSZdriynTJvcTMzY6Dr9e7Soe2ayypSiLvDiQ4vLsA51IBdxQ/JzQKa63psi+/MyeFciM
DeC6bHjpS3J0v6Mb6W1fKk9rliWeTE/M+Lj53z7ZkDROIhwdfWbYMazvOxV9gdyYyFEtDCCKvK6f
XSIEdJwQNhK31lM1C0K5OAiOHNMagKl1xzvsgNck2WFGsBbCnzRKh+MrLwDgye33pG8EFS6a7aQW
bEVhKKoCjkCNJOOsHtA+eRz5vVDUZi4pbcmjkdtOrTQY5+Ox2bRDmIfKShiS9zPq4n2l7ZlPnMY5
qtWeZmQQD6MP1zwlU8JbhVYD5Wom9sCuW6Z50Mq+jbpL6cK85O2+yMRaVfZ8xXF91ry21DnvlQu8
Fav5mCNHni1DdH/OryltHny4R7F67GxTzk6PJK6vyaEPXUKR2hvZ8tXbWKIx8GWmaqsoNplRij/v
hL21RXnD0M4oL1ToYPwN8xPsY5sNgBqoGFC8v2xLWMpfFUi/ry2ZupYT6pnafu5ooWmVBrh81fXG
vJ1tASamcqoOPZ1/yg4sSR0XvMP4oW2LWIqoxcd9X9ve0lihR1RReIKdrXOtJrVV5ojJZi3a+G8k
PJBY/0OPLbmWJjnZQatQp3D6tA5KTgONt9AoorqakhAM0e1SDIJh7RenpujePrrmITf0KOo/4NTa
DulfwTyUFsZu1uwuVT7kAxkI7ti/bNZbbEt8yVX8afNqCjLvnFFMl45AKi34/i1xsPm3cYY6Eyac
XlD5Fp2A7vPhw863VIv5ouroSY8AZBfKFhG2Fa1Og+Zlgcf65W0tWz19oTY6Tpm1PqEDrK/Fv2XP
zUyKQ6P8YUpt7lHL5JqxqhGHQUnRk6JPItNmo+HpvaDfJU2zERGiMQriQAAadHrqM3UolVfFhQve
62lEqeh+bh5YB0i+qc52eUeDmB038/R1QkTHnw43vE1AVdRzVRswJcrioFNqugm9hotvqPIKeGgZ
Z68gg6Sy7/eHIj3jfVxIyuIdENS/W0BzXsaTaebE/otbKLAUZv4JnTuJk/qwpHTswI+rzgjl52n1
05sAlu0Qv29ZibdMaYjtT7pnCyKmPiy9EuZ+2AwoJ495+vzuTSW46/zpd9bM4Ba9yzcoMxIRc1HY
qseLcWeGt4x0aqP0vHeF8sisQIGCiUO9AOK0NwvVaq/EaQTzuZe+iZk0b5lx5Mp8EAiC2MkdB/dG
0HrQOThtx84Ypy3dyIQoaCNZzK2kvXEDy2OKcUUJ0tT72SLaJ9SR1gXBn1+oXihlg6TA7bt5KRqa
lTCt+fjwKJbWCbrIV6wPU0Xk5mVJ2C+Fw6YUJyPyloYMBTxqZWXXbtrIjieG0Qut1Stc80krL6Qb
J25vfU/KePuXO2lfOBgeOna0po7gzdArkuk41MceVDyFAEHs1nbZpT1qhnh1xORvjDjcDVPimnBk
ATacCthM5C3yZ7lU9N2Kt/yGEBJrNomBoZJZzlW+cREZizt57oofgKEH9Bu6XFcp9v5oamNTj0GM
Sz5RCJyULFeGJOX8NvTsmvvQ2O621O00DB15xvXo3mkQejkSAcQBux1c1nNPdgaawVyP4VQ1bQBQ
Vofvtx5kk/0SVJc1AHG0xqoecUStvRgSdwzE9M/NQfP8AgTAf/jJU58f+D4Zlgqpymrmejveula7
yaRTX6P226UprwqnNbkDuFcm7NqO4J1H/CQPOfqiOLZz2cqiJZgn7yYNZ42nK2UH7UFga2oYhL2t
HKyXQw5ZmN5LGFEcXBzV5fBVt9Ya4vwaqyjbfcHef2IeMpJ3SubXZhvOh1RkjwjO7fmLGny+8/dA
zFBY9qBa3/KAHWKrsW1Vwsixt7Lh4JJei+29+CW7CsjAKjp5kUSkSlF6b1os2ztRdT9x52rhuioL
Ls5Fnn6vwIYycqh3kWgcU7Z/CWbUS13WYf223WBQBYQY4AMTmSnFqHeBFaLJYj5BeyQiym0YyBRB
LoUF7ZoQm1xEQDE3eotENts7V+gOOmfaftnZjsE1xOTNaaHJKlJvhTKOWjM//5s5xtHMr+4K1YMD
AZnTq3YjuMu2Ii9FkeGq7Mh3vkJEnpnBT/BVq4E4+xHS52wwtPtGSYcg5mIOFnE3yWTZ7mDxuUMh
OhozahSUlCRJMQ01wtbsu75FJ46+Zk9jHdMNQXkD1g9BORRRSiRdbjyRth4LR4VSC5rPYdyL/72j
HDHL2EKX3klcfXhhfRyir45VrmfME5LGAH/sH6W6Z4TDIS/lSuyMogX/lR+7mkxbq/2XEv00DRAW
VpNbfyjIV3IQrspvUDUyMzHdTp6JQpV5n/bYUxXimYmmiA94FmlefeBhzizY0n6jSVaGSe1KuEue
Dk+fUBQJmaz9sxNFU1OV6Dh11zCJN1NE9w7+NCrVw2YkikutZefMt6CDTW1KvXzcAsgr5JP0rDjh
dsfOKMpgt+sjTYsQsoD2ZA+b6MD9ZfBla0L0zm7T77jTaprYvFAMVnCdFpWDL2VRTwmy+wRpCh8S
bn5nb8sP87ISv/yyMilxnPMPW+UNgHHM9080BEyGWdlwK7zbPb9WD5HxltjnJiOzEbvf61MOUiDA
PO6D8VbleOPidNRr43n1kHyd5PRm/kJBOtufb4xQ2sSxYAMNuJgxHrCmA831Yej5a+c+PBr3rXhC
tBCbsKt8+s/fwgQ5ZkKL7i8c2+ARRkm/DnFwJPhMUdE0kFunVxvzdGtKHzMPIAabHPfJ0o8ZrNEH
ymDgnlH1JESHnwDA4Lq/w0wM3haYFcNAjht3p2O076tvR/a38b5b/+3ubS4rIHfBKqx+ED1JUuRj
3P7F/u/VGdVbyfd7Ioz1xsLpZIgFVWFynEVXkJuW1lwbOew4ROgbKC1k6D/HyrtQFW+4B9KqVCio
eOSXdlze58tK2LwrE1OZduzn9JRZx4lUPoWaiVv93AHVgADeZ/xD50DFhsC1Uos6mYcel89kTejE
WJruLhXqFcmtVEjJq6joL77aYGPmCasJYM9DAHJJI1JAki6XtDDJEzvVBIYWUeq0OXN+5zjrkYC5
FjCcNsZt/dmHLAsfvS7Dajgub06seGHBPV583q6ZNPsMJxV3UeXRzgXTUQL4SvcOYniMKVzpwSya
fj/yaWramyRXrb/PXt2xov/1+zWMM0AiW+o0UvM20omjBgTtDM1scwWv0SsJzfga0WaiGuI2CQ1v
7O+5GdcTyx75Hp9QZHCmr00kqo7AhD5Vtn1M9oHkm6D809MO1r1Br/4/AbVR88985NqfdXs5vmnc
/43+R55eiZRWMLoO9JL7L4eLam6iZX1t2vRtdG/VYYjuUq2EersxSWa2dfQHK2b3YbfNtBv69cvC
8z2xmR1glEZyeuovxz0em6qs8AmNk1OpocX5cwlObc/EBLGETm9RVgkMzZyEIil4GEGEXMoHNkoZ
9fvSQloIOYvlRpbhYGTWPsPbOzX8KWYkwsMogpxFwZNlBczNFNI57bSgzPy+x6jUcuRfg0iy/6Ta
M1AMtWhe4AYkDJeE+CWctjhVXJ65dWjfDX9p5VLH65toyllkrMN0zGugbKKqIMYTx8UGTkHkqYGB
U70sa0dEKql+yzIGWWZj8OLxIYkEvWSzX6loKkDCj9rPocuBvlS42au1nlmbpPncOtzWvFC0Pvuo
cFYv3uqKg+rkiecmmvZbm4zKNzkJAxYMrWeUsXlgwJpyteggkX7G6nCl4jjdS+2TwdcscODImggj
a7paMGjzBCLPbtunFtbkI79TeEldZnxxRwMjBsBs2s2BOUzNLNiuc8M6y4jPtr1a/b5aeTIRYpII
sYjoXjeDAr9SNoxrjPSxGqQ89X0zml+m5GbmmlOk3wH5/K2/VWsI51RyVBxyVSBFhClJd263t+a5
F89hHqzBRdrldrvZIVD3T+kp4xvWN2KIybzpQpI4XqSPV4hxzq7TrTRtzEINNYn3eGln0aC4PsUF
D9bezPy4rXVFGATZp0Lpv8ozlnJnFlV3x4VYaEWvn50Khmt+/qXtWLRQC/vBPurbDiP8Rb5wS6/Y
kL247PGv9FKHacEkM3qVg3/7AUCctGaW/9mmkW8aKxL2qlgqOboFomRGPDiEE1+7plLZ763POVh7
GuKxV1B0lTHLewLV1KqVw8sYy2DM+HxZ8m57NH1P1Yp+FpA49lfrmp89/XF0tjQ7/QfjSgX3vcow
KKXSUUCifgH7wU/fACS8gWPleD0pmx0t2XVLBuqHAhcYdKP8iavmeCaXGt3+o1RONAsuDUmIEdZO
zVWftSk+iPbG3QgoI7GMu2tO81a2zzt+DLp22dBvyfS+PXc5EBFMkDqaGzetkH2tmF8E312ZwBub
31Ap+IIyK3OBJuBuu9RZMVl8D7wOH5YKD/ON3AfxVWMxd1PvZlTQ1Nf3yM/IHwhw6WiosX86jpP2
+Zj4sQBztlbnPd5WKdTFO/f9IhyJdDWeafKMd6lIeZUcAUxh9q7KB9ztCHbCQZ4WUiiPI9HavGjQ
3TG0iPcS/RXv2UhfBWiAJrH+JGDDvWJ2gsXQLM1Cw/53S4PjdVFdmckOkG8a+0bBJVTF4dh6271I
xyQlYec5Pzsk2QKn0LFVZBGfix+HZX2TJqMX/hHRDNiPOYJZ7k0+eVkf5q91BPn+zc6F85ZY0YBM
qGwWGAIgB7TUT0hPvBltUWDaSyHMkkpoqStL9lm8QOR/2yLlYS6IKgeQaGAS0kqMlSAIEXkR3Kgs
6pxlfMqqYJWQxY9frl0vZVcE0rdJnTH9vogQ0jfAPY3IYnh6PvfQ6AMX9ljHKtBVIfsSutnmDE8O
G86lkwBcVNkIR2AkXIZL6p9f7cht+s87pkh5s3oaNKnDGFAumfXonfSIo7vAlptu/OSjsQg3BqHY
7+rosHvs2tfkPYrnR/gI0SDW9PAnBk2VvSKo3pblk1+yCM4u+YWCuubYZZIFm6itBRF80YaKsoyC
wBUvFnAGJNiVviNJ4HCIgKSsTquO++juD/Ormnm25gRJTP7fE+Ce+Onc2ZEw+ILjRqASbvhj6bNO
VWb3IFEYJfDoMBVZ5SfanXna4mDO8Rirec7XkSEpFMieAc6/WqlQFzpgRvJB5B4QL/vP47xBWo5K
rPJ9j55xIKkbfj8o7hzSV5Utw6f3JS6zFt/v2XPToigq3G8sR1qVF9pRFYYN2DonD1+2/jvGEnjH
MoX6dbkRmSd7SZ0sZQJhObbkntOBSUOKMUsPZhu30gV29mEes7yBjVfFBNOmEVDYD7tPJ/LDzW9X
Dk7w5jep5qCtgkR2fJGaVf8aKvoRMtduD5JbYgHmXKmmtaKV72FyspR/AAPTa0YV9/ymYWCSStIY
XYRkywPIRSYlb4aR8IGydlyCWydH1TpFGsszrM82YKN6FNdZ/obs9E7TFYIAEGQvhwsf4IAJcefk
8InCLILh50gJHKRaxAu6xmKU5bSqy7ZgaNtI2EWHSwLGwoaCf5ITxSMNfpz2C7THwgr6a9VwCX4C
lJLPu9GADNxP17JUfLwB6QqKIYJW+ga0bRJzfqoaJmDzr8i3Y8ekshVfloVkFIcWBCFfik8SiU0l
Xn6Smf+liITXxdtStRttEtncbTKZBEZ9EPCZngKezT0C2LJQGARLHw0pPxUp82MR1Cpmn/Qs6BUT
5ABCvsHUSHUo7ldjyah7JoQAAbyqtOY39CeJyhWKXZy6DtBAW2XPuDxwj2Mx9S2MD8N6np+cm28K
V3qx5y/Id7JhaOBpxKnlMsvX1dgi9q+dMDqhdcYAFdC5SFj50EH9ustYv5HY8+h9UPcafr1N/AwT
8VAfU1ymqYoc2vfAUL6NCyien2KuP3cfGpihk52pbddAGCS1sjHUZVvG9RNW8xgOgjc0SHyxE1UW
tONMVt1zEwyUcUDcT1i2II0GEcygsB7FSanSk8xBgoB37rxevPWaWl1zxbp7QfgavNlmFNXEJDtX
qYWHkRwYjwjVYKCnzqDT+2eZUiYfF+jzGZ0/Jmd2o4EcPjjNvZpBLs4UNCs6hnjD/qy0qZSewygv
P5wPsmeU6SudinVgE8IPHxjoln/57v+0F6XoJdlqFjblQBMVhYyiRQJd8hR4pKB7ST42BZFhE3iC
IYhFHm/wWHktVuxje93iNuGyxGqy1Jq9YRvpoHQ+soe32ZP3ZFE7UTWF2EsBLZ88OfhBV6Siqp/2
MjLSDWApfq515wYBCEa5Mx9L0/6yEMzvFTlKYUsLXMZDWabU6YR1WosmhHISHBB32c0d3L94vXtE
fq5MZc+ajWUUGnAPZHB0sfvoDdehkicOi4DOb7F506QUR71+lxkGh0g/0mmVTf7SbVSVOfH40PRA
b4GuOOF9QfSiUc2vM11jLynnCKYml6G+ldIttfj3G6UBJIv/9dYAY5tYAIIKdd8jKacdPFMOc2mX
GAPA3ebClOfh3jesCxaaP2oBHfYCSfMHn6s7rYlK5l2s9clhFKwMdzZg5Q8J3DaTxprauVMfE7fr
cjNSWDZZJConoxDh+WFjfQO2qy1wZUDMVFcXNKT8oFrJD9MIeAiK4p8fwvvfEBJdcmwgfHjucIuc
P1IXW7M9VlZ2KckpFtELmrRoSeCPiVKvtXmUf5U2kPxupPBYd225TiCsuwacO/0oJqLjLeu+Ztgq
I2axNQNbtYwqMbA8DLxjYLOma6eXo19faVSoN6ccnoPk4FJVTJFu6mHwQGGWSg3ewsvhKdTlqOcz
toQxbHVF+ZOLVaHR2g420uEzQsDZhJbl2IPFtsib44UmrzalkqiZBWA68geeQIV8lwG9xQolX/1o
iyHOMUzR6oipmLhVxHtGGuG2gcwJpHA48ohf91VtTR2haA8HelUyFqcFR2xe7MKmiCxbaxNyakxd
3BjhCWdIuUA9fX8ARV3Mhukb6/BVS6QWQuQ9S3AHiEVpz7d9kDVXNxCR8rY/AWXCPH+EaHc9QOcQ
2sa5gadqpBbZ3WF9tkOdoeflYZstz53Ihm/M8SG/vGtDPH0kFR9V3GxE+hXscKYCWzP+rNDJT/e3
S50Jb3yweSM5mf/mCLmc5PAVrd8jNJpZ1tNN8WHfiTlcpUSLrxz+xKtWTbW8RZloVTdpG2eddOUB
5ASe0RLHNFyN6R8PYenvw62MtZfwJutCc4axXwn2PWDJu5Ku5Q+2sIKb+iMOMNeqCV8ZGZm57Hnn
ezJ2sw2Zvwip/7M0OqtQGFxsO8uTYHub9CNQ++eVELCEjrslCGYGuyqt7FRpFiJcxvNmdZanxk+6
2GYBdZVUP3SRoN6PmhAUh+8f2GopOVh2uYfcuXCPv1zZkOay3dwhkK/yqD4hyTHaibTfkO0YyXk/
rV08p0ZpLq0igvCf4IRGwYq2sMFssHviWpiRatM+E2A5Td55kfYv3CW0YhgSEcmHOLW4QAGZ0+si
fBMJhGl7ryBMvM/JwmPEReujAT205IpwbpQ/uA51Kve1FN5P19unmbXxTClHKlXtwiYmgjsJb4X8
hHXy8YQV2fx1txe7sK72wNI2q6eXD67WsVbzmx3i4G/9T+aoKcuOps1za+9zx0e19Dq8eEKBu9pm
ZgZO/Y44jaG1g2OfxDzKuJJ9gr0wHRD66XWF+vzjgMU7Ihai+69m9ZYfGjyHDKkn6Fp629CXrOBk
q2wxwUyGJeP3KjxOLaiqipO7fy2cxayODUFcfAHOJirddUN1hrqPs2Vn8zW6xDN1zRlAs3Leryh7
mwsWMBrTIQfeklvOIJa0PhYhIsvREWnb4cRV2SShvQr3STgfEJSdNSCQh/EcuEYiKvBzGQ2c+VJ4
VVGQtrUmNavUhanW1gNkvYUNq0dmtsCsi2ataCxNo0FizQgqaZLEAZv0NOLSHPX2UlaQDPW+ySVo
AE0Vl9w67YhMtHk/ac2iTJJP1a3O3FaNiFmWfzvFdsI5NZVgtd/BGzGP9SobP8n1qKJCPDVkE5s9
QrnE9x9g3FQwFAhbp4DNqCowpsFQ3KRN1ajlrio8t/oMtwtqdXxJ4QBDaxaXbz4FMFgaKB26R2ls
P3nmliZD2LOVPahfpOO1gw70GjB1ACYH3hxMedYhhfaK/PDgq1BTLg2XpEpMbvn2suSHNWoaGC7h
NRo2rko8+TF/XX6DxMShPcTwPKwK237vuD/ucDztBS00Y2Na3+peFiKmHeQVLxTYk8EG1ouV9CFP
YDR2mE9c4HRVoueLRy4HD8xXFPZ/8aP0js5ypUFFnF4DzMyTxTfmgXFTnN2eCMNc7R0H1Twk3n/Z
LIl2G6K5jQuEc3Jd+LJh05bJnAQLw0Vit3EC2oHwmerGhn5hGCntPr1juRmncCvuXGaPE2jjjV+4
flFZu2fgXNfMPYQR50rJpa7h29tC6RnxH8FxMuznBrCqi2w1TTzG2INjeApO4zPAe3qO7039jnG3
5E0VReC9u0hAWN7l/KXrtSodTINW1OwrlZn3Hl5kBJGg0IMczM5bF3CV3QIvo9140vGKESaSAx2d
yHfbDYSJnOBmy64WC1tCp8mKZN9EY2lSXE/qgyNh2R0y/6uXNkHbJHdh8cxQ+Ip7uBJYPwp6TwSp
BLBpeZJPCl2L0qRUi0+kXoqG2KsG+QeIpsZ+dmaAevkaQerPRcVZXNQsbhxY4JXyKxBRDzPNxiSM
GTq5WbrBIGv0spLN/R5+J6MBP5+qPgqZGAoFe1jXYL3QNS7GM6Q1dz3z066du0pd2QqqYdZAZtUl
KeUXDTJ4tiGccVe5TdfFCFW1T3Fca4GHzrveCOtoqKV/lhCQdk9O9cw86g77k49ieQzs/B9fCrdD
yvjB66Eq1rBKByoERzQ2vDAQOOIvcW7JNC82nTZczYrZBYezQbFBXXrSw1c3qJETSCF/JpeYwRrb
KYbRBRHhnLWu/XN7MUvgu6jqFwM5esnI+08LN3o0nvmlcQOtRIYHL3r1vKZFMoIz7qT+txQIFglv
uYjATMICwNV8AtY1MAOD863Nbdd/wvLmC58sYf/eoWfmKpjwoIZ8h5IS4fyv5/+pY9YSkAHJQn+F
ScveYgYayfGn+3uoRlz39gQWjiRQ7v2/NoZEop6HeRtKpP+Lvcge/7drPx3/Xo9Qqg6/+SmixAeZ
AnMQEY/IM0qjxVS4qPm6racQbUjqRfEu/k4Sui4uq5DSj+GczVZBx8Z5UZe+lMRReIlHwqPzn6bJ
wP26GRB3R1JUPMsGTNh5FaYaifQ9m16G4Un/fwEt+ihM2K3MPK3wPPCfONxPv08oCx+5v7aTXW5y
mAONpRbAaoZkZfuvGpyu7Kp74J9qQJFlyYS5V9u8fSs5vTcc3NHN3TzqbJYNsksaZaS5xtWVU4MT
z4uJr/lUY8EjOydc7qOrGr2GPNQEWpV8cOUCAb5x90A7Gz/bs4a337ONFVmDGoSsFeGZIFjz0T5l
jgKVioMD7hj/YRFaf6Yfp7qdO1l3jSjzbZHl8umHmmEgCfCYkdO2eHQ1my1MnpGh1Avy+Je9+sN7
vOQ7tN86JYSep/AHo/CQx1OD8yVJsl8Wctx9i9l8ks+lnIk8hIw3Nx2VEd7s3iWO3SQeWGSPr2eY
Ohq9mVnjMNZC/bp2v5Su//TPSBfH8QWtYFfIzkt/2fr7pI+8J/J51InvN/yxiAFZzbiRsmAEtXc9
cHwhB4S6NGL60MMz+Hmp+alGDMW1ztPKdUuNQDDGuuwAhHxV/SJ9OqFljKN7Lks0ADDrDYwhzn3S
Htwx9m4yb2LtvtVBYIQ5EO2SzPndpb/tcUuIiLzUM/YK995hDhpys5BYcQW18LuWB83zQVRlmaVc
kv5DLsaXee2ZlPUMDVjuptJSbIzgWlO0T9cQoXTkq/bvaKrfA/Ieehigelasv7m0LETNtb2Ok8T6
puQPfFi+QEP3RmixgzEa7+c99IY7bRkNIfFC5EAK26o8zAZSPlWtNUsXOMmUOEJiTxT3lqe50YgN
rRdcnBFIYy0lOknvQbSlGL9KQ0uFGUj5kM+MnRIlZrYowUlWw64COU5unC3QaXu4PtyXSO5t2Mk4
hgk1oXDDk52FamtCOHgpcK0WSxOi01+dydf56rFT26zmNAebt3kC1JPgBC2i3Hhm4lXxQyoUkaoO
+AG7eosg7TwqhtNIGhWqy2LAd+430Sd6JVmvj6DQvep70bVHIGvfOhmB+DALHvUsJgXv2rAi/ICK
jD4TB3teWvoTiVqLLxC+vakc3JoEUN66/1iGi423Iji4bTKg43rofHw9anayvf0GEMfzV56Fg4NH
bTeIe6WZEeGXG5KDsSgEsORDTGc5vQG1ECsXqsIYyC5CYcLE3EB/wepOuXCcg9rlVeWWwLRIa45C
sW0PXKGyhTFrk4//zpVlUJpdpC7f5SO1bIDWhrnUN/PvqNpEWuGKBwfr9qV2Nzq68dGRoBDOwbsM
8tvjPEGThrjSskvym2ug8fXk6rysU2swBcXdG7D9QtTx1kuU2294986jxrLKxMGNCs+rKNTTqKj2
cNyGs1DB9nFFo7MweHH/+comA/ZKyoj35RuCWAdQTJ6RURjnfGLy6r69mbuEUJfUj5ofizseBbUt
YMOx4+HRTqDucdeo23Ft/jMTdve/TAjZVd+r03++HGA1YqFT32hjzDfeiduwH8AajoMhDmOeMjnZ
SWDML5zf63HdkmDOYvAtyuHXIt+CRLN3ODQXZZQRhFTy6uL9Io681Y0ZJM1SgGdYC28oITmKmVXf
QhJvVlT+AhlVG2l16KdWsKAVKhMsLAtQ78GEGCO5bupx/XGusSjbQGTBVi+wusTyZslIGBlvEQPM
6VNclVbrXCaOz3ELOS4SlZJb5NsTYGq11G++ow41TuA/DKPPaOnUDX6sF5el2bpVrvit0A8CySXv
TXN5SSiDnTjLvJ2a+RjGVF1wy7ygLJFdAe6MhrBIdzk2JlVQ7INF+B4S30jkFR+yH8UDH/4N/TLt
crqigREuBOA+LoUYNXP7iAx552W+i0vSaooHsUFh1A2cPLFq9EanmEPwK82xQaM4T/R55ESPQQZf
GyMlooEFGPF6/Yfu9JmSjJMTeGgforJRm83RQ73SNah7N/CIj4BH5El20r7JS04gC8CSA1KXx0qg
8gUvy/0UAZL+/nDFI2DvobJyRmpmklF7yf5CTNY9epzBUFjoD0jlYN0JLjBTLOneqlsBeepjI/eL
l9ixKaNsjeNIrpHm9px02S6a4L2sDQQdgC4VjS70uYC4Qgjxg6v3EuTfDjZ6mGZ9YkTxBMW9OvZr
ergUZz3xnBlVUx+SiJrBmzS1J148pzLws5fqaL/HiIdtQDs99ZyoQSYHC9V+63wYBNy5urPn3ziR
5em7zkU83z1VmRyTo7qyVAcss6m9P88AUWTNYmSvQT9MZnMA4Vke62Zn31X/4nilD/7+643xgx0e
abQbxaqSrUssHLMYj9pIhxGeF3USoEzjVwXK7n24+X1Uz6WoVpLsMI7Kc0tRHPnT7iulurX+SS9y
L13nOcyRRh/J3vGnKFlqgsF4LRk0EyTpjGLI6NPxYKIKmLfTrdsMH9reIxzsmzIA40zVRsley/0k
SoXEVfG9l8/KSfxN/YjDZpaxqisdzQIKoig+hEKzjr2TUpnmuNE/L2BiS+vIe5lS+TZN12hlv6A3
w9F/IIuAaCWqa7sXO7zhHS+IOhDe9JcKuIcjMn0yyeptsG3AyHyBFbLUGxUTXciTzrMJRh8TUVC/
qP4sDtagq2gpOqdofuR0JVEXDRlDJDgfqCEdBKBPENokS8+ZfQZvVsAEE4L9h/mbvRWNMfuH1aX5
DjT3gJ3jKSEjH5WKgvMN0hQWTozWA65ci5RyssWpiW5Law4Os7T42GGJi9P5SOC4/VEpAbTHUHCb
OUI7pQipy8HwuH/ifM5eO/hq0Edt1HyiTBGytqhplVhuKCwwIQoAX0w+t9RFZ73ULkK09DDRxJ9a
0WtgEoX+1w88W69wL4zV1zHDTTPuzxuieXWLkPQyUw0tlssNIY73pLs3wWopWZayR9ZKiodb0xVf
djFghbwCUrkmA394uKVA0k1TvQwnQbJLZeanfkvjmCJfruAiLKMYENT/Yvs+Q97mqqUrsdDtQhUK
a7MktwasIJOOjvsbYKjAXPD9jk5nnT+ez9U9o3iIF/7YwyN4ylNdMgD0sizvzYx1ny9+Z/7Y1Uy2
nTFNIGEp45Mo8DtcKEPlK6SIPScXFwHf2YtXS80phbMSgMVVSZ9jAwPSjYfvcZbiJy8A4yz7TRMN
Y2l8pURdRk1CrBFoJN52CmrsZ3MmyFPzuAzGpizGqJmZlo6I0qT7sGZXMuvGHx6wt/UAZphAnx/3
6m4KuozCB0YFP/c5v00/p0Bdg93kuupVUsUmF0wRNV9Dwu8i6NxuRLBS03ZbTr9w5MVeffLMCrX7
SqzOVwF4I/o0sJhRSZoVTIpAzZNo/oS6ZP2j6ZpMtdOlFLj5k+EU+YvaeV72D6DIzhOFgKiS02DL
FwkcRF7pP1YQ9Ci6uYjop0ayRIMW1wjHxtQZLLCCTG4XXo+qgu2kunjCe3ozgBl1csSla3rjnP0+
FuBx239drYkkEJrK83BnijloQ0Vx2ZllCvgDhtLy7GrBnCa8sAWDgE7lwgfINyrmTo615GszMBg8
iTgWfvxW4jSSqzgF9d2U75AMdMEWguHRgObJ9WKkh1aRV1mOtSAMKCBIcdSR8Kd5YG57PkNUa78Q
MTG4f7JlgCVGognPzY1TAlJkStNkiNHmVu8vWdnfiZhYxPcYawSkWQjsxXcpl70opsjC7YnvjcxL
tG7ts0uhBaclcKW/H5/PIu9rsfHSYwWzny0E8N3qRZ6zr73c+wz+tDI8E8td+sRHPUaqsjtNPcx7
m8wEKMwmxzDeq2CjeG3EIayzalVL0S/JfEVc10YR2TXyEb/U6ht/VqcM7LGw0uCn2/CI5Sd4uYR5
SeHnwptVbmrIVUFPxdzhQsdsdP1N5rvqRmwWp+DEzWKR0oLURE+3VJY7VDneaYHM3h+EWk1YDmZp
993kuqci9CgW8Iwso3Sxy6UfSTFqYP5pC2sc0z6myqX+N4cUvHBgXduqpgVm0XTmTi1QQyw+Eznl
Vj0ePVj+GRt4dlWkQSvdPur7LUAnFjQ0cDuVNW0ho6uu09SK0S6Ayd5ofBvuyvB7Uu2Bktp5cM2s
qJ1eVkvl4FKyhnvUrSnad59sS6FgsM1C9NudVNewIUOst1EfBUB3Yv1xFAcefomJcPNLFX7DEM0I
3lJrcHqyqlfCqIQ4R+vhWNYlU08owF74B8ND9VLsrGnW+A8Pg3FbOadDfBEvfFyr2Cz6VHnbUCs5
0IEmniAxgDnco3FlIbWx3FTSJj0FqQHiGJnzdFMmpXIvbZK9z/Rel2NBL2uIq8IbwE0Xl1KA1/jI
a/QDTLud7rpan4zGsty2DCeGu/0701NfQEzkpPco9/KfubRWnInujjEyvvnNtL3xAWQEkXqQPRgp
ya2Z2GvT6Isq1eALJL86CLFyqInq5BWKbYECEsMUHWnXiqJJFLCQCKWkhbIvts9rKh6EkIMyfiu5
UoTi3S9BlN0MfGUjEl5TfNtqVtKHJ3oN5bXL6834zj1ChEhncQm40g4WyTntq8WSCPvXBUI0mE2X
cCOjR5SZCvm5aaQ0ud/B7M1DLvmGkht5JwBRivdVBFHmjuUz3RKR3LpO6i2MDWSQJos7DRefO28z
1RqCB0KP/JNgsze2DPFKCa+IZBYxByN5Njq1swW4DS1itm3VBt6/vv8c6VI52uUtIfUeO3bzOawk
z3WEMx/ER9Ep0auyH1roukWmSz8nJhLv/UN1681VDmuiRW/dsdsE9rCCBJKjAZVosWtA31DT7/Oo
H2IvISOMYquUPsEMRS+0ACS0Xc0bI2a4HaQ9RPxvDxO2Qje1IB4UIyZKNrnl2oLcRroJ5eTc6jLF
mmn2Op7lArPABLnAyddaGxcmZPBRjxebhS2ViC8ODMUtXW6lChNApd/0oyNbKf2cqM6kGBINALrd
C1ocdgX9E8R9XYV/dHZkTiyekN0rwni8eRyEshdelEGJM6HKxw610Fhu7IVCJ9pS7KkvSOvNWRP5
aGRR0pJG987DzGukYH/Z17cBvQoQwSeu5nXDNGXiQzICc/eET76Pn+yzG9OvN+a4AeAb7frbnPBD
NnAZh8ibdpxtX96u0KMhIlCzm0iRBEuPQHJxE+YKUSMZSi3599lY4jIDW59EucjLd1KmYWeLygLt
EZ0H7gD06GoRbYi713pHL1XU1d5AGD+AE+5BxWU/3BbW1MvxICyHND2j5p8OHZtQPuCAzuer0IHp
uJCb41c5zVrQPnkUByrByXopVMrKnqvVMGsMtMMJLA7IoJraOl9/wVIma5dFHv3KE0R5a7eWkx8C
upMADg8SGTXVggfYHv3Fmj3YuCjgRYnuJGdN3rnR/ToTLwtEVL6C8Shp8fTvYWD+islvMKaFmoiA
BKN7uyy2l2CI4a6BelP2Vq+xedophxJB4OFqSDTCrhj1cIR/bEMxA7sDJbKg+zKdiBov2H9QmywS
J0vKeR7y9dH35yhquclcuM9i2WT497kFZhuMXCfc2jEecsGUhB2BwB5RxgeCJcgZtJMoJWnwDYnA
LL3xx04Y2e8d05Unn3sunZXwJ+rKORZESNXff9gU/c+YzrWad03qgYT4asO84A52YJyMHPEgDU/T
pSdDqgWmM6QxMKBSQlPx27qR8Pn3xpRQedP3tFihuhPP8atm4fSFJRsYn0WNRebRSx+5GdL/ASis
VRcpeI51ORn31ACpz3uzavptIcpqyrh6wlV56ts3w/fpnXnOBvqk/Z5BhJlIKbRRVZqcXGzptIRF
9TB217I11jr3BKuK/gP0YrbfeHejQAPDGCNQ+a830CJ82Ot2XJgexgyX9PxqoNLW4qisgTzhcpak
nhC2He9olV6u8obtpmFcI2HOgaFsKS9w34yvqVXTrllU8su0+bnYi9kworKpuVHn56D8GB9ikeYS
DazyLbxWR6gAo6x+mBmiRvpY441WtdUrdAPX+b79Wep8T5CcGezHg3LrphQ4YVLfdLGCRaRx6K5g
tAvEFf5WC6wXQ/fYKNyUoKXlfr9ksuP12sWZxkv4I45JcYZTtCuU4Af1lhlu9DRhSRYUlenzhOCk
JI/uC5Eks7SjmmwWY90YkFxjH58jVgrH4EyHHDtGMZIeJz78khQpJ9oby5QZWMAWuU15Hjxo1lnf
ETiry0/2u0D2ukjs/Mrlq7HItHZLiWoAgCpBMp4p5NCcrczXiOAJuc6DWxQy/BYSOFfAqBgf/UCs
mBTtvhIS8Gdw9cKyrVkFNCddrqvcjSjcIc493KmQz1Sv5Q03xBhtDmIiTVoGB/QQmBwlfj3uCm4D
vgzBe1WYsS47GoWhXTMKPRUjb01RymkxBS02BIQfX0/qefXa5vncFAXPWcGPieXzcvTKnoCy/PNe
wnnOGPuKnsvZyhZ3td5pxYUqIfaILTSYs5WwthAphA5mkW71zA2Dp4iD1lh0QgSX9eGboTmizdX4
ECBe7RBJnsrP99mZSviMU6hwwyLoy++Nyv0ACktLnm7ukBAsECrk9tQ/Ida7JQsSmN9ZVhsEXrXf
t05QB6t9VmWeYTjk3LTAn3QspZLbSOCbXGs2zSws9t0uJTTxFyzx/XLA8RtB40GivKH84lvPhE6v
Fq9vJkHvyrVOrLzJoxfrXQPZ2DzfTzut2YJdfCIFigCfgtiVeUGHLVeV7u20EWgpMdkfTwkZGJPT
APP62WufC8US5lOER08YP6VbdTTuyGXfSAEB90MRNj9YBZTaUrqg/Giq+fDgBXqAZVLo2UF22/iK
t1GFnWUrhFnWDaIm9C8WQpXuCs/8c5EkdK0d9B4tLOV73qs4RmEMe8IeyRQoElPsRfm6Psrzg08d
XnC1fF/v59TwzJcDj2q1EV4d0xzHo+TwB7cJteDxGJB3TWdPdm7eZtYVOLeg0ukby5NNdoXD9ZQX
3jzo0JQoD9WLHADh7CrZ2Rnw/LplAsqc0PEcpPDWmVYwdNUBIW72CO+AyiUstFdm4Es/tkNUYVK7
NLuf//kLsQJ6rezhGuzMXpHqJkxIuKH39N0mjhjJRoDs5uaE963lhP1svwCAEH9kfwXFoXiomqdD
LensqQn5Hf21OkSH5CKLJKS9W2X1d91JEq/UhcVi9JrJiU7BkV0zOBNZhjvSYqcqs811RmNAb6Eg
1cCj0eEiOpdcafvkNb1Qm+rRz5yg3/RAW2YuCAhBGPs7SBnPk34ZkE8dnc4nOK2n48b/oBQCHL6k
mG5BivGAV8YrEWVkH+RStpstQpGkIq7B/r16TWi2vZKasCO0WPEG0nXNdPcBVJgcESccAo6pxEeh
v4P97vnIAHlAPbeqcTxsvy0sFXjvZjF8hzAX0TAk7S+xycn3QVhxzylLHd+0ZEriNANXdIaSUVAU
OyZrAHkbdB1/PoDXsVZaFydM3/t6SrVXIkK+MimD4njHLO/6YGbhcM5S9cPBP/R5NLcaOVsUpYyV
5oDhqPHpT1URjuSOBBtEKS20JgJCCfeSEcwbkgFmQBKkSVWEtswBut9vslAeLhuDFdYFFIKYjLhD
yH79z0lvSdRPSIFpxd38H0wcRVn9O1CyGTSka/67Q0mq3hBmW8MyPUCXESCuXnD1ljNtAxAtX3Mo
3hmTFIquSaS5D6uYAY0GnIHPMGSIReARlO91Fao/m+1d+O3mDOekSDuhKQH7x6OHJMl99j4haNQ2
G1sE+ITK0S/4FUqSoqYB3Mkbi5W99NSvh6H/CM4Uu4ihKBXRkMdEZ68MtQNjftzlNN9OfUHxUZu7
FA3QAeydbdNIsSYWVAirvWX2EMPfYITYxaebUUp2xmXekrOcbeKDdrMjF/dsXc9+3y6bSUvE2hin
BZDe4vHTuubE0VFdWxZhhMwx/P3QkXn4e7oRdP3tvg5IRtECecrBcj+MOkGEsPTCeBlTWEeoxsIw
bm7VYFKQVSUJMXmoSmKfcg9uJ2A9ml2ZPhAtWCspkH/JpAa6vVC0njbXdW3sMb/oqQ8Yr/xnGDIg
a6okkWPDpgOaIqtW+HV2WPjkobxiKZyY86ZEbnVTB/Rg49qJVB3ckJxXr2i+5lWLuDxaz4XxquxL
h7xqrTqQ/YtnxU/a+uNlOtMhT7q4QFqG/EfI/ss1n7K7x9G4Ee5wO9R/L8wRFaTiqrK/lrBeclLL
Zp+7oTP5P+G9Q9Sy3YVZ4a9LUpMRhWk0LQUspTGiU0UsUBAETSP4CDACDjJkqwvVo+49An50V/jj
OYqng7KYeQPjtwyk/vptuP9Ywyybmg+4KAEeOGjd6y9CVgH68UTnktP5hcVyX9swAbn+p+J0rsuF
QUFiJRoZdvhLZL4UTdvyK567BuDQnVp6Qez+tD7cdMZxUuEcAf+la2xFTtQBY1tuZunRUcynbht6
sVSeBO+8kIRU02hMoquWGTTrIVaAJtYFRmyyFOveDtFNevCNmv6Kgu1fHvSWVVLct3Skuxwbm61K
P/XZRs7HRVwdp0ke/JE45rGG2WiAnj/VRWMH/WH+p+QzX5d4rXaEZF6bLXbVOnG88lzUhXpSuvOc
bXFI4O0JM+RP6ROF2HnrB1PWltRSnh3QXGxEfQCFkUEaIR4LI85IfQSZbrnM2qbjddVVhwyXYDi5
ZVdSxvl4Uji5cvsd8W5m0d8spywj9NqMRx13xXD3YTffkSKL5pxYR+LZ3u8ZzPBf6e5qibbgJL5m
AweXfFH1JIsWWLiO/O4vxN/SopzSJikGd0HRUpExQH+F7qVMjMFO4NmDpRl0T7SO2pXPgFWcmWCu
/N6K34r65y4szgSPGR0LsBJgVY0MOR9/iV97QmXcFS3WYOVpTz3wJBcBk4e2nNsPbmhXLdNhV90I
A8iJsdRm//BECS2jJgfovKLG2HceWCzNnCyB1X1RqTB5+QyXoNyHVBwPlEpYDfBSPknGRxau8g9U
PA+nGHrVSPrGipsvmipifb0jh4Bm4xXMuW6IKmI24O54LVEGor19TGFMUWGZjFijC13/ubdOROIP
HKsVFu3V/6yyb2pbRVp2nDBlCWx3Z9FLvjZ7SJHOgPQv3mOwRpF0O+9Rhy0pAZqSUwROJ7faMuJU
3p3AlGHMV+1yeCUum8fytGvZIhA7dfEy+3U9fK+5y7tc9RKHXZfdi+i/LOTWBCAG/iGe+vtHF6tf
L97r72OttinhB4IOFg7DhHXucMcMDY71/wKbRTQHFk1Tnxa3z4oK4EBPxaWJ3zsq+5r54SaNudd+
+c8bD2OjngP0suymiSMIadxRSjWeclN/7ob6yvkkKZP7W1VQsEUfX11qwejB1F0/HqqaSA5EDXZu
hQqOq9ua9hOKgCDKL+YQ94nBIzM8kQdpnoZxDamkk+/b9/AmujpO1ZCVsycQS7cnRcLv+woWpgTA
l9q/F6R6G5faOCoPcW49p28r/RTAl9FUIDlb8NPHu5S4HPrjTwBTOD+SbKtpH3m7WmOCFeN8LiRD
QWs4Dwgq91ygqJ70hkMSc+jQdXMRUYzrTWq11ICX0ifzq0CQQW8nLYo8zTPm5sGQpAXL2Ce71kwY
iHSuxX78rf15N5Zn+V6XOctXFf00wA6nOdD2ycEyGQou551MmrKBFXZAMQAgbyz3kd7Xn22a7OxQ
X+9lY32gQDuufASSsH12fmdJaCeXzQ+EBx96KgIadUREY+E/3lpfeCkRoJHY+Iy2ePtmlyefZ4bB
RqtsYwWybPoyBhAxh5v7d8e4wc8JK4ZTaCcoa7b81CloQHNrOFYapnPJC/XHFFfvKNzDUwKIqcka
Xmc1lJKZLX11lGkCX9HpJKgiYnyDQ3oWvvXYK1aAqy39LY/2Ki2HPLGXT0tjjHhY8acYtfY7Pida
0K3qadrxl+kOXiaQGaMd5FjLXSj0+Uvr4Ijs8QWaBOnWSvh0VhLQKvYFlje+VT4oImZeGYsWG3df
XO35C69oxWBpcX0ENvlfTuA1XJ3k4rrbG0RI7Usa+56IRgIOpDj8mS+3GwHUd9es+yBtkZeSSide
xRKnilrY0wsspQQpB7V4Qe+g+vwQK6Q75eHxEad2zFY8BvcGxhCs6mkjblP7fLOq/r2xK3p6+ePy
bHGPMAXRXUtCp17tZDek4N8sKn86ZwZJPFYM8P+WsiDY0k1s64SkTVDkcXcmp0CszA5j/mqD12YH
GSqmp7Md4YCTQhHkRkdVw+HgV6pu67CvSx12fA8CiN03kxPJRQHqs4hZtsTheidZ1Bz6jL8qNMbK
QZAos4JivjrtsrDV2PBBl2HnJoV4+FZqPsRe3KFwaRtOiAtg0LsQRT9LcSbo6ISgfG26g91A1LCK
AuSq4Kcc5x4ohduyaeW0Xm94K/qVgTAPrMJZBHFGNOsvZYt3yCR5fYAuHwDTCvSr4Ucz9Hgt3Kbm
/OjHaCQ0LxobYNSN4St73ek09hqvCArASDg7CyxpTSv0MhPyLmOklu7wdhrSaACzL9/ZvDHazyWl
VTTAsZm9NaVQJJ3gfIzACTZx0Wau+FKDFMkfSN8kSM2KdxvbQ557jrAh4NjuF4uQz/cwAF6PwvDj
jN45kvhCPf4B5r+omsOthrnuXxyc6labhk2aDyW24U5WHmnpbhiRdG8CV2UTBcwsuBvTOA7Jkn1B
Jc23YHYwvPQwRciEyNhcqyp+c2ty6SqozVKC1NcQ17Wd/lNi/AjTOyFYuUcCohJNaspYNwpzoMo4
iUiJHVdsL2VTy6yr0ln31zkGz+/YYqTmSdszaGc+NWciFFDsrCJ/0aJEHJHmvbL6nPYgWjo7arLA
PcCMElugKnWyHb5mWqR+ggXnaW4mZGCe8WjkpxUMEMdYrMXypNa7sz5nQeu3csQfQCY9HFKF6LIB
D0nBZFsWlkqsPLf/JwATBi+14l8IEwDYWy0hCDiCua6bxQ0nf0Vwa5CqSXF/fb4Uym607aVuUvwP
h4eKBhHLfZTGhb6iiRE6uApvi0ZMSddAb4yDoi1C+yh/TCEa3D3Ii8UsYI0OBaz0spR4SpsTDrF+
boQl/M15CI4V9QNfdmimLO0i+JUmWWGlFz49szjWLNFPJ8y65TrdLz6M2I8y4Wac4ICI6ug8hlB7
k4Ry5q8Z7/Usmw0JkU1a3vTI6Ohnlr4XnMPV+9QUjAWOYm5jLwDWw/EVLU2RvpUf4CKnjl0RrXVw
DDvXcZx3nqx1caliimKjqQqVGmKPsEpaEH9tJs2w9ldtpW876cSdYZAf1Tk/6sacLAmQJASY11w3
MaA9MjMbn7Jn8Uv0my4CCJC9QT1dZNVMLVCdSNyxadYlM/MDGdCPF6CyV/9tXFkjbZVjZlZgcvNV
HVqvATPSZx3BeZjbVDzyiztpFzsFqoU3d1Tz14biU/B6r3cRkfZHM9uz3VZO3sjxJwDnqrb8ApLF
HTGOt6a8UpH5NIf+3vRGTAHYG6ASCXzVTOZFeZHwFf7C3lw1GxBlyTQCWA29/GL4+94WYvmoAmTl
iy4UYIj5i2BJXlcUEE/169Z/fUO3HfQt988vQ9WJevInFYbHipHz4yNyyyBL8s2igNNoEPD4/zRQ
JiuWvnzwDSTzOreuHlfZaMpB3Jm8rJdvT4oU/DlYk3u9FOAJPJILPjmmshg5xlL+jctthbF+5Bmt
EWzRiw7X9NJ/E/Ay5e4eISWzOZjGA+eIMgK1fv7M++9lVYK1j4EWKlzrWNAKKjvtGQ9Xdp2o68le
LtELIsE2pAGUrITXKuskOKizeNXsBDW2PygR/23X+bO0PFRM4SlGHfyklm4CijCOdkZKEfRxs8HG
2tJNJ2xK6gziaOPOnZgL5H6f7nPUATxy8eDkULUsoyeMeokbLIw5blBCSrHuk0N6lfHYHjhgWbbP
4EAivcx63q3NRokawb7Hy6CClMcNkpvdMK5o0JpxDIxYPco7AjVqQ5Tf6MqFg+MtZGEaO8Zcg/8g
FV2NUKnP/CZaddumJVop2440RbYOQf+tvtT6lEXJjjkUAG2iLOF0tYNL0eEekcRs1CZrZ6p6W1tq
HNdfjZ3viDt3SfFS/WuscUjL5YqzP3BqQ4JaAn7mnw+CIs6bM6uy0vQOpLb044GjPeeUYDj1AsTt
E8pnS7sDxHLmZJTdhCA3MbIN/dfqIxqk0TB0Cq8XNAWVH1yiXUFzUlT9P+KsBcqTawLhrHN7N6Bl
SCHjEGRuHfe9e/x50cw79oOQ9d/o1vRyZ6DpgEood1sHYI/w6ReK8UZUpjMM+rUR0BEMDh4EXzil
XYSkFqXVQTuPaQgGGvKvS++JLdxByV6YSechh6ltZjdSx76rvrn1GK+8LDAxTCsZKYyWYVdE3Dls
r/qjwehYR1SjrX/NktI8x3GEqlesHbehuUQ3Wv5sjIJo16QR/p1NgGW/Mc/2SkiiIix/nckunQor
AGtmmXXjUVydqhPemw77EMeq22dMzxvYpEPnm3ajkW972Yl8o2XGq6uD4NFqPnvci3pCUFOvfQlP
TA95TvQmrZ+IeqqLff92N3wku9MgfHqQx1aQ+5A4HWNqIdG6Br/uBYqiM254pjD3v9Dj6z0bSnTG
3EUsr4rMtC1JQRP9Bbn2QmSKRMPnQuiDcfs0mc3uvdCXljxSsUQ6/tl14zUPFQxFoqNTNAVwBACu
TDeEGKgV0upnJbj9ad90eYLSlPMyGdX1i1+Qw7eDWwBIr3Bs09H7GPCApfMo/ng5pzBWEe7JxNsF
Q2HgQkp7kA4It4vNLeMG0rHBySVcyb2w2epIc1kDay7gVwGMx3sT4d/o14kwn+0vw7EO6aeH1P+h
X3J9uPp1KXv5YwmelNyeSj2cZlVVBUOmj46osioQ1zXPsMILkPfswX3zpkF8aAev64ZkfcSuWnU2
yYTEGDa/pF1lzrCzdISmu1nsLTXV37D/xElZOpgkzt7gIOGMzvvlPhOTJ7Lg5UBWNPW1n7vSgZGt
g/CuAviWczGbv/ygGbP/Jzz36OHOwX9rnKCatBtxyeMdMlSaIrYayUoHvVmIayQxekgFPiuVhaif
7QDYWYDSiMyPosznaj6sZ3xe/PE0qnK2LipHQ7lzwVo+Zygj5KtBaAmXvkJ3CsMSF/XdrGW06jSJ
zlMz6JXCC97kF8nKcBdie3LN8a+kBZA6VyQVl9nQCqWzTMmrc5zq27t8nh6Z6IefF1pPv5pIQpaU
jjdfFExHr073H4/U+bJwy6u1SiuWHv0EZbH7KV0hycd19zq4Cy05OvMQ0ABizPqAFpVojbUQeQmr
SiW6PmwKdHDYzM8lIuc+9rtLci7XUmCNHL0l5zS/ys1hnR6aNwrQlMD5D/vgE1+3gfgr6VezbtQm
azBUCLBw6sdmlOEVMvRxfEa/HJHqD7fSBYd6oxIRPdf/mR3i4ZMN2buzpz2rnczZWhksKUopSi3d
iks1L8bYGdcJdmkcBZDJEqgGiaHvl5a2NvaEyxfFZkzwhNbzsootrfs1EcvqlXR5l5JVOERJHrYf
gP/xGrPdEkCKRNXWxN7+EBCaHbDjM+Ye/mLr+8Rn0/Zv1wiLrynMfzdUdP4QoPaQeh+4c20mS3zt
qhvtAZVsVGeIH4ysbBPpYbTbZ8uH84ckFHyFGq78a2DWrvQuLi7IAKHmVWpC1VrO6mvTQedad1qZ
7dQ0vTeFtnbZS7EhOeiCnUsQZH5rk0ZQ4M5UDvm4yXuyYhbitvrzT+HKJDAI2dI+zBvtdvxNzxeB
fUq8a9tmesu5kEWmTuGrHLm1tJCu7pn6Z3Af/QZTJpKCBTulVkZJC7ogiIxlIAKfoe8KZFfc7lpN
3kRuLK2nPufv0pFs4/4hVvTvX84HAEpfEEQZnQTqeFPaaanOBM/DWvwlUUOLdmuWSR6DcBjPKgfK
Gy26vwAJsxyBGd7vLfBBsOW1+J7YLJI4ELquV3SjRbWni2ku1CPoRmdd7r3kdnA+7aW5Umm/naWU
7b1RdYMDwThiUcFPAgLQFkgDNWdpOPhQnU4UsYVP50wRN9YYD1/ydggy86SO2Rsoh6jQAo/EijkE
Cjw4/gG3d/Z1jM9ueFB2Do9MWSnCBtfBUFWFerOrrlwlVPROj4lk36c/tI888xg3v6B1hF6DHfEq
pnWA9xEVb1m5o8otHydhOjx2LXTbW/yKyihYDH7qt6EUrWFUANzsF8JNihdKQTiMyZS5yxKtxQIf
xlnSlxtFDj8UF+O2s6/fqUHeAeNaDslhukRXoQ7VOTpjY7fpwmYOEOzO6cAwwIhYmkYh1w1cHLT0
9Kqu5l4U/7Jh0fTaCS1MHvKuONbYdHoWgNdD+k3jSnVvmEYNbWHecCyXLdcKPnsddIRQIqaDTpdi
Z2LKCQVtaTj2S17k1JDfSle26zKvjK+uEWmJtXpCbB/cNnS4nTYLEEcQ6j+Sld1oltaLIFOQijwB
Ut6EeodPZwK0UA+j2a67OIzjXZyo4Z/qdbLH8HZWbp4AUrf214KTi60k4k5rvLbozjVK3NGn6dqW
M60OrZ21dZwt1xvK6BHkaON4zWkwiRT/TBhZdA3RoCyKJkVzXGyfQJ8h+hYxK1U9VRUHhoRHQAWm
X+9UAPW8jXpNLHdi8oAPXw4scgaon8Gd4SMQmtla0sxaDloE6um5BwMA6DKIJr9FNAxzpEmvea7Z
Ul+reRsL01Cs1BaghM2D1uAvP8wwlvasHsyq0ZNXhRid+FQxJYZ1t9Ov7QwK3GJBu460UQ6atxiQ
Mme3eIUsVwJaH6Dtqagofwrgtf766eFyMN+VN8zLEtBGqYUTX0O5nSDuwu5aXFpnWp/n8gtExhpF
wYOOATsLFz8XqinDpO9TjKFwCuLq4+UDBDEM4KT460NHmQ/LCRQY+o+9FvouZGctWJmMaItbrzB0
UX9keyUXak6QrbP+DoD81eVIfQzgI6EM6TOb7/YJwAE3Kk+9p4XKie3mgnOKFZvVaVbLiLfvc1NZ
SL5vaRPSHsC4mYoRLek9s/JUuwxxNQpuzaeNufCnBPoKNAE2UBsyQ/xETvs9wRw6qmrI5eQcW4VE
v+W+vBF0C/r3qvG/9xFF3A6Lps2xJADJ13w+2EWleq6gU3/aTlF2Y/z8gjRi0CTDnq8+4YoauEYy
BbxQ521n5Z9gOBiMAyIIXnhmTM4mjR1v1iWdYdYSk574I8f/s4J0HQVLrcrIMEhJ6gRJJFRJmM6Q
CyzSvXly5TSAW6Bh03Fg5ioSbTrhz8zVps0H3bQ5R8j1gMMrxqxFZX1nWzZEBglteV4iV5uRarzx
91ne4FYqtiNvWQ4ZTJ2sEAbHOsV40SVVRGnQR+waYT19vCE70LNq8B81D59oY9NkiWF6u4SS7sGX
hQ378BLC6QLU5tmL80P1WUz4A+7zRlZ3GURyQ35pWUosVLWdm6sQS+wlyYH8ehmemTNzIJcr5z9p
VCWKpWXtYq8kn0V+DxFG5luv5JS10PvXfnK5kWd1sGftWnU8qTpYplLNxzNzUl0j0i6lQQMEwRzd
sHhC/qC/Zu2SR+TUs5SAtAbhhtOjxFc5qYx3x5MhafU2Yd2PaqeYXMrllfYX0S5Zi3u1vqEVBEoe
KKHIJDzu/luJ9GfvLqkjCNoNpr4mhOFVej2zvAqgliogY30PloCNndB+EGYaS2xMh+15OwnMnWUh
eKJe/rwHl5L2GJifet6QKwf7rZpwJWKfdFIh5iD5MoKvSNZ40MVmCPYK8P9UKjaRByQSu8gCjT/N
m5dmWxMJXdfyn8svqi+wmVYsoPTnNDb61CM9ewOGUxLN+tMffnPCcGW8U4V8mPdWY91+DxVwpQt6
gf16iaYji1OvYB6QUDNpruDBCMZjVjgojuIotc3eCRxQWI68pJtIhFmRjraf4Z5KCVBVDX/W/bVx
A8vQU1a/SS9O+/9G1MPmdNGXCxr1XWxy7knuHIhiquBD5DGgOXwFbwCnsWD/Rgqp7QIIZtH7Zq0S
xH21TA4Z1k+J+wq8Yv3DBtG7jxjNoAIx3CWf1W4aGn/888f5PxSAWsPwaYLG/WiVLrfk9lq/mrlk
Ym69k2a5O4rFqifzZa38vW8sxDv9cBd0M/xGIH46iZl9G4KD6FUQFLTHZDDeedNoVI7A0HzcM2QF
1943CUmdFeRieGcC0pK3anVv2V2KCs2mVAVaaSoYFB9DxCa53re9qPbxchJrmaHunO/FrAhugzhI
Dk2x+mSBreQLM8JLjc2PdZZiOoGNJmUHrHAHa1mm7t9F+n69+oCunXuiAUa+UmJop//59NDkOwql
XZC20z8Hv4ht0gW/6MtzWOlCV25xRP1DWbqO3Zc0JzQI/b63CKBPfA6RQclqBn1Hq1FtfDm6K3PQ
l2Quj9CvpT9Fy2Cz+oIJ/qMU8quRjxP65Y+jcVj3t9yBbaETx740f+sYb7WxCQNmHT1s/HaSpu2T
Vfc2Y6n+R4sPUThxueKxXhtTREYXSXXdzSeEKCYVafKpL97SDsH1DYU/7QAFGsZi11RsfzZNQDn7
l5rWPuZJHiXylyNkGYMzycgfMkQoCK0kBh7eGsxL0Y2VC1fxsyhpMGzBaNfhjDE1JHTOtVG0Ryl1
psxErRvY1izNXo1jbKD6Ynivr3gfEwTMsvevNFHmWRQde3YqoptW7Iek+Mh8VYS+dX7DMEYbzefT
4UqzZKoeQU/NWNAikfBADy7NZRbfXC+OnVwOZ90TxHp+/LTmeT/LBic4GUuW8zdlkw7U7xrIIc/Z
3fU5l7D9an2xXo9elJ2YSgC115pX6QiMeOHjC8iHXwjMlOYhmrZvLbUA9ftaqYuqbbyZZCx9nEib
bfhu+yvDn8vqB6qhFx8kc8JpNYbOw/pVf0u1BrbsyMD/4nC6fYZBKfyN5DinfHapZKh4CWrz8W31
yUBSmH4ZP98yYVF7KZkBzCsjqBpax7U3XaNQZrirgWJHSzARVLrDyOJv+wH+bwwIp8k3xWeXJSpX
naylrkd1sY4NFdlq6paUqHmSpL1sm8rV0wblWsdY6lYA6TDfZjSQmsoae1OHbcg+0B3GWlTUBd+g
DCmhFsm5NXLRlIVhPtFrpAvbMxu/yyctFNeWUgcfe5tjHkHWgfv7biqNsKF4e3bKmeK7WlJch5em
IElZNil2OCqH9Mw5o8hfsFgU8kohBEMpinF3HcvQr2iRNQ4Bxqg9jPWsqb0TBSotPxapMdENIpKm
N4ecETIw2tShxvnI7FsPCzfcy9QXyUN0EdwSc5J0BKgp+BbV06ebr2CbyM4Myv3bUZCujwvMKj3l
r0KHTiq0vzIL40UmKjtlQrzzYO+egYnFtL9xAUup71wu9HOMzkNytUwXe44VmMARsoxspgyjuglP
J6x0Lcs7jD4SQnR64IIya/nEgaPjL+8OnxeViSRbE1GeW7YBJeKoqmLmOY1U+tnoX8Z5Fjyu1d75
3jfZ3/WqORfFVUCiMlKeaRzL9pv5/l7eCqXTKOQRqi+nxhSKO7d5hvhNEgzfRycXo2dZ+C/V6fjm
qPDnjfaMezAfmWvhjLE/ualD+6jtj36PaRB95dEaRhhkFjY8SC/EfxP9VhEy0kGdClhkVn5o7SVG
mT+aRuYv/4EfThaAyoFbAN1aEKNuXW7ijPuRDv6eMgse9CdR3qPn1heQwXhwTXeMZ6m3gW5roQVy
bNiFMMeFuyOgpnPV9mVhd05vT8q/84SkQXn8LvqxbqABN19hX+K6sTSVCpfABOID7MdHjoFaMXdA
rRQmloLSg02s+E+BlGnjBk9LmKVAvKaFxccnyrUOHGJ4zhP4yINSwsCHKrFoOS/1bvEEEZXy15DP
87+5BoWsBAXvHryLV1beXSwvbwyfJ65sVy1kXBO9kuSk6wxeovKpF9JB3Bkl66halZFtpvc4HHOD
GkIrmf8KUhXvxCNDC5MNVodckVRn+WOCVrd5MvWQ/IF0u1zkiLeyX0torwQLZ4tCRGx/apg2lAgD
dnHppoAhreSca8LxMskpoi9/GX0iZl+POC+BG/3XL/q2GHqgDv8yNCUOfF0/Zun/5W3kLxKHmNh6
HlUAPQunPUVu+ZZtkCcPQMZTVsUGNPA6SsK9A7rTpTvtKhyBvPhyaRqJ+mBeBNXkbVoqeUVLvYT+
QIVUrTgMs6PiHZA1MG7V+uuJ1GzQvLpiuuAMbGNVk8bsX3kQ4rKKySJPSPSPY8SRPEZJ6Kp6xUwW
EwW9mObKDWjXw2CZHsIu6Ug9r8CDEC4Kg/SRkDEylXR1DhZcCUdU1kcULwxDBjTc3pl4n+CexFRs
9/BZ6cze8bxJuVVuCd+nGGSGwtt8wZKorU5bQqvDrYg95gYMIay+v2ApDlIdz+5XAd0CLcFSHiQZ
GknrZW7iQg8zPTc1ddaK4LQVD/hdkSaj2GncKpzILOS6BZdPDZPKbjJ4QgnXKXi+REFCCsCRyveG
K/f2iIJT7J6pmSXM1H65GYGJhZFgp0tvkA+EzZfu96wwBWafMCmWNTBesOXlcvOmSucL+DmaSJXx
Z3QxOy1A+Q1Rm9lZHQlqi8psyTIqNjUMirnOqD2VrRqsr5q9C6kQD1db0772UZ7McDb/navFvqCP
8TNAEwP111fs7nOoXPLpNv4ORg0VMwD+21p8WDxkWC6B9ZKMbsLNybFB+VKIvWYtnTUf79SbxgfH
yIo+eiZiauJMiHpFssKuF8HXbbULlvatHE3TSRQH6pB5MsXymDXzYpuFc21U64tHNywvxku3Xn1h
envjpGcJ/uxiSzJpzkRu6bQuEeLe1S04VjRPNlAKBXReXp53d/n1YPH29tECKRits3D+Dz7mwFH+
aADMQ7+gf42kqod5OplxhlxGGOwlrSuADbH+ovYvDerPI5BbjOLrrFdaH2hcoCMtw5/+omWGqiLQ
FHMYusxAouDhCpz1xR9P1X79kNBRNldR0SY6u1mQ0IgnbZ1M1mRmq+N9dgGPpD744+PfvjuDuMaP
Nwp6m1FjVDAa3RuIv4txY2yICPzZDr4t4UeY0TiDxiNnUMkV2N3kVCblyKwkdWJ9k53s/ennErFG
BMxK0+1K0B4R/MbTmKPYcixLubmloIbjTyGwf0t2Em7nI/UCZT6kapVgUEw+jISeucXOqvnCOcG2
5/F/kJv6eTPQslM9KWZmJrBcBFs0561kd26IiMbLba4MjkAA+DqKaoAi0uDu9BhuPdnLMsMgt18t
CfPm/VWLfYG5WrDWSRsMtuowipRP7XBgPidKTj7Hodu8saNm41VgsFXl0suYzJU/6iXjohuByrcw
8UEMDNeR2BhhvMUxS+/MA91h3Hoe9Y+PsLdpHZSreXMAdaRnz5OZCej2QJMcuFClvL95tAPkkpKq
obuztmqvdNm94YLeESkMMf2aH2/eKMTcRO8fvWgvSnb4wx4szm7HVGh1ePk4wxL9lr1zbrr8B0TO
FmkYK6ANG/f2rTZbX91CDSrtnKVGRnQlG+/a+v+s8+YdeMpH0gvnrd9xml3+RkeFU9y54zHWd9lF
kS1UVkD35XwjnbbqnklH/tF+dqqg7NLhPKTzAAFo9/uBlbbKL/F0KTqJMnTjrI0uYQdwdeB735Oi
VrutTf3wdewQ703Ul4FQMRYF9LuinK9QH/EJlG8UMrns/H3LY7UXOdIe0Ei619O2c35XIgUKxDTO
rJ0vGLLS/13N/T/XEfB2cCDWywZPfSXxZo50HXK88a/IFSxJCQV6bL08IDK0qXdY6dSo9ySFFrvh
qaVCtXCHnqjOa7hKP6KCRpaY1UFcrQ+GrMGpSWea83NidWZMYgqVGjtBBGz37T7BXAd4YtaJwnMO
M+mySn8I1yxxBTQSH5HAp5NBEu3ZpQYg7V7ASVS2X4gU83TxGnoH8vlHG+5xEknDCC/blSV9GJJb
wU00cQlw+IvcSmK07dzVh4ZA1Lpk0PPgE+mrdJTbtANpDlp3U4CX9N/Ld9awec1bkZ2ENQTUjw0I
u6gEHne1waMF2dUkfRX86uENI/PDDytUSZKjVwqtWLAPEYexCb0B1bNcbtNS5aOkUWXSkZY7X4eK
FVuCnL11S/j6Rv9h0WTrHMSE2sawKvGagfo+mK3viR4WJwjBBepVQZXLXM5oFNIl6hTV7FVq6Zfu
G9mXyJghm/EgtkOqx9Du0X6E4IDE2PoqELLODxjCaWVk8H90amTull/k4cyYncEeAGI0pmq608N7
hNfvlt7UFyFQc9Nv8nknqOKmOXWSBQuR+OP4DuuKBsn5OID5lUusyyXlRc3pSVvQPKLOCO9U5tV4
sncQKMVLMCf595pyw8zO/na5yKvlhJqwbtIkBvZiEzQoZParCbTbM1L5JdrKKi91tD9ZqChkhAWQ
6UasCiKKXS3B5jjwKyh1paY//Ze+wMOuPsfaE6MymF1V8VKECkIoo2Hy1gaNZ3rcSWrYSFgCNJTQ
NmAjGgvpO0lpNndECXcrUwFS5i17DRNnfA3QQQDkhCWUkUioTqBNljc//Un55UjaTJ6bkVg7LkqE
5uIbR2kQKqH0QFeNYxrYC70W6BirV2/Ce8zfWsjEPHuAxg+X06iW6KvhRJ4m6mQflCu5F9Qs0Mx/
Y2Ue8wNc5reya+K8bUd0HwiKrs0UhPJPgyeYDcgRhpVLWdEdKYuB55YiBpbjhS8hHTns8xIUcFtW
oVGGTarATN/8LCzt6nBoPR4BPH+IMugb3MgLPrxbPvMUDQRFY3pc6VOgri7+KRHLMUOP9YZM2LY3
D7rD2kRar7IV4TmT+4vDNoo/jNV2STES3OzI2fQN2qAbwcXbZ9RQQJrkbdr2VhAQVZbZLS9tujLm
BTcUzzzBh7AMTOFLF0GvbdHim9lOnsrLbdOcuEjdYOHWqtb5kAZtA+Fzuhcv9JNWiSQK5tQlyyic
wytJauY8ueFPwfkImIju2y7Xbxwi8XOrrRma6rRBeBVPE3B/UU5XSSwNCVOspFH1mqLIgXkY8Zs6
EY2xQEl4AzjdN7/ArFVZUDNmI5b0jpbxvcKvuiQ0pW+G8lR5ZLGQwuVS6dFim2BiKTxTmSofc+07
mN5PR3IEZeY0gUe1EX/PU+C+KkfRBkewGWVEqmFbGfuEHxkQah3zur95f5e8TNWlxW7mxnsEZcPg
cT6hPy1Dt/dPCT5XvvX3EXQm60bvvigvTe28QirvOvcg4bYmTXmblf1cwzMF/sn0xZ51Nug7TFxl
MIKPnaGPcFDTYZ3tbFXwpPAJS7hOdACWx4YXtb9xO1jHurRDBgEP92OUmRUYGcw3Uc3D/Rpm4/5T
qiIQPVuKAfSyrm7ygaab9F2Nj5iq8LT8/rYAk5ffoB8RvhhYhHVsrf862mZkeZW2iN6cD1Fb/EPh
4Kh8QqEao+2d2lQcvGKHFCkEvlJHhV0oyEVSUuJc/OYxtMm/j+Mbg7UVJxVGl4a1tv0+i/2nWYAh
+zt/lLoCIiDBVN+n/OzibmRI202fGWpGpj/TnOLMYH2D5D+98rTPuqru9ESwE+cDagycJTYwPoJ2
81uiqNSgUnIruv/YNZbTaZJ2CbnTp5Az1uDQ4ZYq8L98f2Me5SEZTBDylagL5w+PFXL0beRRaucI
LZViAo0Oe/A3fDvQzXH0Mkc7ufO38x5vezKaOo/TNAke7Q6L6rJHfxXjRPCAg8dKfKRcR/bLGjYT
ttG7AO2+4kaIoRaqHKFv59A+XgMnO8LhJUlMiGIQQ3Q7TD9QqboAsXBb+ZaOvBYpLqVd6WZrXUhv
aaEwGOZOViBv9qijFvm5GhoMZpnijvyZN4i+S9+eLGHS3FriY1ar/7Svm7BSKZkxnsdyQv2GRBnZ
+SWCY7FRheqWkZGfQbT5esyFnCzC1I5lNTsny4aAkl8xuZ8GokIqYVihM/K81W1sLssnmahp4WQZ
0gu7ScZtSK/1b2W3iyynH4ix6ad/aTKxNZ9117ZfErgeRcgwFSfGEmqHNtxGtIaV6zII1WcA12AD
eMY+6qoVUWHa8bHgpmPN3BZQ55973HD6JS7wlGF7Ezc0h54yzYFN/mw8EDzuztHG7l2to82KWG+f
rRHhCRDqhXHborjXHrp8hm0AFz0OhFyxPpI0nH4umoFqpBgoXnP8ak8SoJxPjWj4dCuX0Bxu703M
YD7VES+ZYUXL8lZvcZhBFsLF3UkDVq+TbvLUk59c3teCWahCq7jA97fO+BQ/i8KkMTpP+s1RkEOV
tlpUR6fD0JbNtbhDK9EM1AfR7mQvLpJOeRVN7OynZ48L8foHXQHRxyltwm8tRdrV/T8RuNVmwH+x
EonAwvBTlrYPy/HiX8ff+ENQIRO78eyjBsoMh8iSUSMx21DfOfoWDeY4aolmGGRzcgZi+Dgz0+di
A9Hr6IAbeJLXMYIFP+4IetIQ38eDgp6BybOHazrg8pb5BnJxkBK7Sl/YVrqWW8KeP9zdYp4+tow5
GHG6OAGVIHTy0aPpZxwKVcetQed9ptzx4kAdy8nHBublmxGsjl276P4oX29j/Gyxy60Dqz8MKraY
nThyx1DF6hfGbDpBqN/vriyos89Yeph0VRU1fkKxp1bADcL6loyTTLjr9iY1u7tHXbWmcyIzewNn
EE7fvwIiQ3S7oyTtVARBkba0RWgpIKMsBtOdO40bPuNAU7ZODQ53KnsJiNIObevNHyjXsolWRGH+
xW5aNy8RTWPiHOe42MtPn0wcHB8d9nFhYuaRsyZ734sBBvxttOe85kU0RpLTLxHSEeBZd1zztS1j
98PkTu+y/DHgMMNV9fJ/KJmbgqZnWwK06rUkeM+kac5PnYpNlWcbvgmUIDxu3qMz+XHuAx/LHI7P
nz88wKPsfUp0nB+MHirc14r/5JMzaLJHw7uvrC1zrHZvtIvoiaHaW0IlzqUVVdkc1h9sGDbVBHz3
ZygeGDomo6UB9bKSdUjhg3JzW5Tms2ee8GYZoIAeMcNg/dhxbboFGmh/ieFgLDzqxxii59gMpLoE
FiTC6zlUkcjI48uec9E92O55mt0UTegFDHoRwzz9gu1GR8t6IlZ5uaFnQXORWHi3vaLpMEdSEAuA
bB0l2faLNplZHWszoXUvcSNXc3OHp1flq7Kd/LndkLXL4rA/io4SDbb4k3cq2JnhCBN2ejxC5CdW
3Q5PtWUprFZxmlqhlt1W73xqVEFT7w4OUPNmh5caIResPX12ZABeiWS4IQrq1CoBPBjsb1VLu86+
PV+InPrZbUEp+VyZyrzEKzICk2VsayTsMqbB1ICgMEz/0/fROS6J7Iml6Vh1DfIMhiYeEzX77F+8
5yKkWcK92r4JR8Vob/MnVaNBH/RSkrgGj27zckQKqYYDYwZXeqFthdBzt5HFa4Gqum6c07QAasAh
PkvH3pZ/I/KaAPZi5HMWhGPZTuh+iW/UhP5B4thRjuO96+ycD9+Kor6dcFlo6d8lMWVN0kFKWwF3
pzQ8Ptf6lKOL4Ezg7ggjOf2JLHwiqK3oCAn0uqfXad16H8XQLIMB2FXZPFbCFrxmexpmvFezKTYK
9uTi4ByTHPoTAIgzjSqLGDRtcAgFabHTE4HqpSGKQ+aEmlYdkIGqvcA/AQCQ0prLRwo3w5Zjv/0s
5rERmm0KrijYzd9S+YeQi6QxYcWJTZRUKwPspd5lGdeo2CUpEYWUU8s2Gj/ONFmfwaA8ODUYc8b2
YPznzHuthVbG9wtsFJabhjLxbckqMyEJmvHBlSjcP9iwyn02q7yXplaV0OdRDg4pubkHU6ZZ3eb8
7Y5W6E9AbJmQNofYkKC4iiJYwT5MmGz4DjBrbswLjYqtSHgt/gDqNmJ2F4FiQmPx78FJe2txFEsQ
fcY39rGACNdNygBdxhq3aZE7E4cGo5YyTsnfgrgMLJtnErLlAF2CQ89Pv71qCbenN5l7X4m5Gq2j
yrFb60zhblhM9UW8jLqS/pgOzO45qdYTWqu5o/0SIY/fjo8+5N/8VbntkI4Uw+hDKKH53ZKsnz5b
zz9vQATA3ucPkdkeXMy+bF/xf4gnWCy9Z3vu9DXVYzC0MR2WURubBi/Hu/5qd+ed6I5VcirmxjtM
fQ9Het/OdVz3HNNOSiMNSdMcDNuYym8ymPdKnQVW+HvFit6k6jv9Hak8Mg6pz72KPW9Ys+W+RBiX
Wr2vYBmFnHDAAhnmL2hhX8D6GSzTTXAvwo2HGsRvdB0m5XJcXDx+GD7RFy3GXHlB81rwDwVs2OdX
CDl1vzQn9HUbBZcmSOQ6Boo6buMuaNZmcihBjPJ5HA5mHJFKj9IUZdUcfcJBOH7YQrKecnyQTkpe
WLAg0Tz5qnFgOfJDgH3Ai3eN0xHfH1K+YhtqqADPV+TDotkzwd+2SRJppAKsKZyUbGlxCdR736r2
BwAJtd8RklPLWxQH8/tRHFBesN3yOXovVhxBuQ+pKLYPUTJjvlgwR97z6s5LATxD3MIqdHgO3xc9
yxsPsWRUUXJecwygNyoOTITSU3tLbBrbZ5Q2gVf0X0+UEcvhjlP9ns4XyUGAIu5fKeF/Hb+P3SGG
WUpu+WO9YgsPzmHllwV0jmMRHRkGyryZW7eFTEvJSg1f6vyzDy8aAtM6rJdfnTD9ywO/6YVlWfqa
D2hSZ/dPjrg15euUbhQ1QjZti1jip1ElhaLUMpDqVZOUieUGl8osEofoQI/54fYldnFvq93e/dp5
wuVmoHZjYNYVRq5PQESQZwYnA3TOlr/LU4OF6U/H3CYLoWcNsYnZAvBWicnwP2/1nbvT0bmQ+wEO
rkDEY9KS4bXcaGOQmbhSbB2+F6hCIegnT2GPjWJgGcQadBp+h0nX4ltqQUjnSMwBhMLMhlyk/CAq
ny2DnmiTtOUJ9ycQGQlPgUHqYuwWDHTEh2T4vvk1UMISgoS/6ooSZIU/O1dwrnjSx9fEGtX//nCJ
h17U8JxdpOH/Qih4E8uc1bk/JFFME9kaClvfIhK/R1ia3+IU0N6i4xoDJQcrwdbaDFK+QDM7cBHO
lVjEQtJ2Jo1Abou5KgNHKCzpGjqZN6h3GZ2mCr+D65VkqWaJlaxOZHB/0WncvRLEJzgFZcjOtNYm
DgQIhx3YNeFrqnTr0QtLdHSY6UdPfrxHHljzGtfuN0tnWuJtHR5jYY/yg2FpC1Fotv5v/ez4Dic7
YHZaeFZ7FFWDgU9NjiD21iXI+OTXuJuAQ2+Nby565mYpm7xGK1WRFsxD58AUyXoDDYKSPd6s+IIF
5NZzBIOa4OVa8uvE04jEzwl/RZjR9vgmpAICAHKbLF0dxYjYose9LR2jug1AUX1H7xVdBtIRDCK+
KyrlppG4r+IGLeHNEsJDiB9Qxw6MJl72tEzHZHKI6HebXq1+6t6OO1afCHzhkwaWtjsL0ad3wxFF
SgTR/oM3zGZKXHGYSsS0Z2Wh2WVDOQathPrwVf2aDfRSSS2UfMEXEPGVpPdFcENk0Xl9TJHstcdb
hVv3cjJCZfN8+LlpFKbCI55Rfe7UjDXFtYxnR26DWoqGFUDZNhKAboC3i0G4KkX4fYUk87zV9C4v
s5ADI9QRpQhEdn8qpIb4bihSw65ZOSdn4KiS2EDKBnjcf9XvxA1I3NdcMb7huA0K0ej9Eyd//ok7
UAfuo7tOWqGFA6cFG3R5Pu8BxZga7OTC68gFYIK2sYNNLQChaK31gt3EKX+TsOHBw/y4N2lqH3RG
ZGEEkkSnJ6epsWK7pGMKiP6MWS4VBGe+jsWxV2oxQOnn+wB7BMVKpwh9dhlHO7NxMYeZ/LYBQpxT
K2VVR06ZLR/m431n3bDdcduo54RCdrpwt9VdtD4AX/OOK7q7nMQ6rpMIz35Ge8WA6JNnaN8ae2dm
rZQJvQmOnELPtik8glQWx043S48KQ07a7E5ZMTZn2PvqPoXpatCkciVkOijztuuPeGTbUR8Gw3cB
TLSqbeYjzS0JLpx45gdd0uDHPX9tCtyJLRTrl3xXHjlGPVapDqgqI7eSjcu6uyQEpZFbc5Mjwt3B
knYriHfITANhY5j9ehI4s/OwcHm3GRV/V2Q8ww36dC3Yt8A7mOIRmMdN5rBYWuoybjOAPnVyGbAi
BcokjWHY2ralOsB289QrqO9nyLO/Pr20kBateAGMm0Tvk61x2ZC4qOolIYABHfMXn1cOJ1nXP/TQ
Fly7f7AIM6pPUZmfR3Wesyc29f6cvHbpGBawzWo3F3xQpSJn0ornriRK75iWfgHG/H1H0ikcVg8W
gtrGwfMGaURujUFG0wXIRuOLqAjJ8g9mwrgObWvXzwnitZ6CfqmudwSv2zgtPPxXXqiC47+PUT87
cbmkPs5qDEoeTD3OiCJZVODEaCiLnJMRpDvTbQ+Lt9Lg+NRKJpZTzbdOULqIrbHxfPR048gkoYxh
bmkCsgWoz+uxsnAjYCBbp/+ZoVFWLowNuUEQe4DoDZ+RNAFDk+lkzFhKJWgjSBHZr8asV2S8s4SA
dzPjG6rKk9I2s8RrdTl6pi/4LdKWA25lY0x5gJIptEeVqtRqPRnyMfk7D9pbm/Us9B/0hX9HeMD9
J6RYO3PdB+ORLydUFt1FzXva331ZNcTeRBLli5WsPO6YtIlLcx8KFwjEt8MSdQ8821sBnJGC721T
Tw9qqjtztOwatNPVSA/z9UBw3OXf4pSDjR/a6y9q3ztlIwXU+CUwStVGNjVFynLHW3QVaYu7dPJ0
wQvFqZwaUgzUFNd/MnntZYgEd8V/XfLaCkvQ3GQ+iHG4tLjnnueFamiOdPdA1LQ/0TEybO0tHl3a
oeZTucGQD2BeKOqFhTl3V/dnqMXp69hmbs1i38k2ipEnlJYJdIzYHLSk+LkpYVG3pZfbE2FujQwO
MPzHbCoysBblspYvzxCm1oF6T6NymsM0G9TmAMr0GNVTZ+h1hXbI6O/9IQ6oYKDvpyoU3dDbHL98
d8S97U1v2Iw1AKDEZUZI6ufDBuItvw2VnyQXzT9PrS124GUsXECgexiUAZNMbUYx2LALE5DnlC9H
QQFZuz3+fdRkSkXLn0iSIdp3Q+7L4RlWiFhWNrMYyGqwN8pMYW4OrlwTbIT+Gob5kqecDpmqlh/m
yf5DVBDO5DmPF8xnTwVBxYuxcniSzr10F1Pk+aln+jk+8AZbqD/du7zjHqu34sq7jtn7a3smCmAN
tWIR24PcpwuOvc9Ffnl3kz/Bw6PHj/1wVwKprlkCGNvaKH6IKnqoY288VUwmICyoF1yksQ1TLNy8
dxdd2OdVnjo0iF1AwJDr1PJMP23a15rZ2VVvFZfKQP57GGLKQeQMvx0hFjqu87wUb4HQCKpKv/Wf
w4VHoa3CfQh0rO2xVV241ENrjFvlNAHSl0WOWeBJsHydz93zCF/VzDdFiL1nJmQpgKHQXZjLZbjF
cILt8tzJJGOF+fEOvdz0NLnINh7jaGW0YxcymYgzISa/5tor5ngdxduL0fio0yoUc6g9Gsg5nMgc
1YZrAq/R4SX+1Lq5ejxpGy+dU5yTegwlvI2/0sgkE0WToIKQ2lpmvWU8cMWB1lqrkDQ4G4eSZfuL
lAdzK+Ubz93Er33EUaOtC/h7lfb1/WJDJ2+Hbi9Rr+Coy0AZdoUIAyudMrJtlUs4UWERZthLma+R
dmTy1CSljUpXToo+pu4ALB0gj1eVGmfoF9zY1pOKSWwMhCIoF5WHH2J+9N8ZLqTvFKg28Sj/h4RG
21c+g0sskixbCqBPijve9/ZLuJ/65ouzwR6H1BvXFrce0AQuvYPL2Xtr2eOahvb8JnMdcY35eyfX
LxYBQHilhenY66BHny80RWGdQlosEDHUIbfJfXJ+ipU5DcYZ0iY16j907SvNCyxtlCekqScXaVGA
57msJ69yrVMVn3/xdmB4tPEOPSyOqn0meTEMf0qM5q4fA9H5QlUWFIBh3FhReAoIHi4CJNzi6tSW
RXzcJQs0J2xZ1hbLRiaJqAHeiv1o1gAYqJTBsV/DcvrLwbbSCmpuIdZRh87ER29+id0KaH0HVgbA
TUfqPhgyozARC+/xjxMDzm4Q0z9K4cqkdGCzeLXxye6GA+S5w/rEyBuZLb2H4z+HoaZyzeUpRHUu
eznlXjGDvtLYd6JofRoaAuf7N+mj/skNdb0lFDuBrF+uGlG8aA228LWuO8e41tqujB/FeZGWMNgF
LHV/4TzpgfGNmMCC4RKZ1ydRZVKFuqOf7ZbKWyeZsQ5XtgmwNHbwOlGOYlAp7QQHSiip3EaFk5Qt
4Y3tKK47cU2nxTdbv0aQdmYkPaTD/YXgi3BiSkYIcTz2xfFP2qS5MaB+AfuIt27MZO0PphCAhHhC
pGw+5cV+rqIRjSTySZrt/OceDrI/SjA10zEIxMtdJCCYoXBl1WOyeF/xhJoKvzciFDjDXG6hjrwD
scXVpORSlHpVjuXO4BebyD/XP+UuZ1YfuDNUl1bzR732vWIfDV2hl0raLVok+H8i4n68GbrtnKj1
U+MOLKfG4N//vD7YrPv0iQNuGSQKpQ/5oFCwYN3Z1yjpQo17pWVuW95Kf/2gRYNTr0sNn/amw4mu
qrh38QPVyRkQtE/DwhrQcDe5dtSrnM+HaHHFSVILxIZTjH552TfUJsoKmdr/RERgXV8uGGng/VU6
pgt4yXRtu16gQWOfJ51IZWG7711RPGjfP8z5tuXX8dKT2pbTY0VuisbQdeOFhZJSQqv9ld0Emphx
h7afZtWg++4Rl3ZZv1s6P/MRn9zVnpPbi1pjx0o4QGD9HZroAMQi8KmFywSPfow2L4Llumlp+b7t
XaqzyTyLHWN2XDg8aAg8r6jP0KB/1gBa0pkiN69UmOYQiuqGrbb69mpat+ZcAlqoOCFITjkfOpnA
shC6SY4MFplaO3caNMU8kpziYZ3VlKKV8F4grGbiXd4ZwYmU+HnfTelq1sA68MBX0XwaziimQ2I7
cdawb2VK5SbfIADVER+SoDkQMcxMjNX1TcGkVJpmXgabUSzDRfta5hRDMPotj/rqez1+49LQURjX
0ym8dwy7yvVrcnxWh3Bc54/7ngBft5yH1v+NTmjWmNVNy/QlqyUhJSlTppZpoYjjZ+eE1ro6F8js
YI42x7LIAxaQ0g1I1gd5RbK2m1sLRgYP98UbKn9DgtVMiW3Q7+Xr1C+yEUfEstMK7AEBJOI3SyyD
sdvFZm9QOpEu6BahqV6gIw85kV/EjxWuFiAaE74Al9e1o0pvFWjfDomwxO9cciohSS1VZBmkNzq+
6J/AqADN9CeYMItc7xoy1bFsNPK6qKqy2WgPvAnBLsSQquE9+enucDM+rEzgH8Wc/520TQ8cYJxl
uw8fjGvBAXiQNZXsjOcxU2HzUF+NsvsU1PCicSd+fFbffJIC1Fcfiqpvk63ca4WjbOLvem1Twpcw
JbT0ocmaOyRRJTcPgF59NZvERXATStdD8ZmwYlS3FMnirqdreOIhgFQ7I0fzAc5i1tzwO7BUMDyo
XTALsBkYM1nkqrGn2kdZ4brsHd/zaP0AbFhoXh7Ul7y+evz8MNhycrD//KVatseLKvp5cN87yeFP
JAzJ3Viy8/5FhiwYwlInrn92UjfnvX/nLMooYzK3s3BlKVXuDglZjkNKlgsBBirf6MA1r1hW4d0v
gHh625qwzH/3ou3w0VmWrozxCvGSwCdjA4BnyK5Rlib9AfNyc2y2Xc1xsGHnMXGfTc+uhFbBDT3q
hgLGluc5rDd5r7HD/IC98YTJ1wECgMk4AchH4jGNiYnkx7TZu4xa++nPwxBieGegH5ad9HCOMldE
+jLaC7IOyzhKDFfe72o7xSauoutjQjFEGa2T02CElw5lvQz7FAhtT+753+JY0aIyg7pbV5Sy0dyw
Y04CTTPW6wUe+XLYmkYP9m5qrR9WF2M1rHHHBek7C3rJqY9OptF8Zgv60rzgdBsPulS8izfQWoru
Uk8h5Oo6CZjFKdbnAYik4IqCrxAei2BfuYmzjFWG8kufOpi+VKAtKLw54QrvC8jSHqQzhNhZGpcN
HSvzvLtRsmeFOyxFFaVz/CxZE4V+ke1S59152PyNQcutdzLtpuK/m4KnMEbQsMfBklCoDxCk3MfR
xGvEa/1++EQ60dk2whE4KzVSEafo/g9C1Pkz8bZA1ez720eG+aiG2+wVtls1mN85B9GWglQbmLMr
dHiAYh+aCir1U0KEVSVnddYsSsVNBMrPZi0g38J++ELg1tsiLAexVxkLGnofN3YcI2zQkj8iRWRZ
UDyOMCUa1VUOQWNZ50mObkr3CUS51J02Jp5VDQW+cfpUc9CxtDHUMeu3Jtu7w8k/iQnHdW5HvGgE
hkRmgyDrbz0FGMUjnVECA9EuVer9SSiERamVqlezEpuJs9vOYNUCVk6x8rDFbTgA2KhSBbg0r/Zr
TPCRz0n2Lzur7YxSqmSHsibVMHPwlHxjbpaNB0VNkfdY972fXtVs3Kox38WrSE6sTdl1m5WNzec2
JsVmWsgG3kJcKPNnMNr5Z3hDCJt5WG1vTFS4B/SqPin1PVJY5rO/NpWGoOFifzX8ccNuxMvDQ0hi
RlIc38JX96Ajc5E/PvIOD4DBdUYze8MTrR7y2zvmqtdsZ93rGqTMhwIzoTjT+o1vuauYJQEkzbXT
wvYJ1QgVHCW9uWoOdqdO0zlG19+h4P6DBaG82HRY8VdX3U2iNzQNhK6fMSmB7Lp54MGFW5yf+xuv
yk5/bHIdG5TXcEJ06MZYzlIT0vFp5PzmkDSiD0SM7mwB5aYVdgl6GhIWwBFW9C7GHcITWvzMg65R
vIFIVVEParNO3Y5izHuix4kRkwwju+2+Mg6s/T7qRxHhTE7v/6koEXNHPpXh6yplp4sMTRb99QD7
KgxtEGzch8lDey/ITYmKBvgD64tRQS459ueLIpPLF/AIH4cEIJsR6lEuZcTohktcbSP8WrygR0G8
VUAlEFFDO9fBuslwgWBibeLQTyCxoiK3x9Zo2t6LW7oZGcYT6dtViCB7H3154Ie/1pk6Dk8ofu0W
9K81lL8f7etfRRjjl8W5dQ+EPvvD7qbEjjk7Z4+pbnKBBH8Gqp5Opr2EfrrvTnB1D4PjXujGnN3f
rVJMOEhmKJO14tg83/HjzmxjGMRIqGhDfpuPUbsxI1s24PGv008+UcWutQCXlSSF2fMtD7jOwg0o
RcaVRbDs9IM53Iutl/ikAHwlT8k7+RvIsBophO3Ck5ahrwLPrPCm4f1AYijAKBlajmJJFbhG31h7
gaLqFnEDS8Iu0oXPMzLWBK0jxQQSllBwezv8gMoXVhu+3VO8bebKEcgKGEv4o2afTA9Cy7vT0faD
d4h3CRFf8VB7E0eyGKcYgBqiyQQnNov6hIHdDl+/2xS0j97V73U2g3pqKTs/AOfS0QQJ84DworJ5
Hr1W/ZZ5DYATOkc5NGDoTawEG+e9Au9ulI38FnopaPF/2+ll2FPAstPz4+7k6AiFZmOooIOxfu0y
80NRvZ+qbsDxIposRktd8wehbdEMNtgnAiuSHjstrJWJ/lzbNW5Ajx4fmCFhp043TzEu8zgQuZ0z
FyHUyL9g69j2bHT/UL03bXsoNfidzf7ti63O6OjC8gWMHOzoid7h3PG7YsVr/AYRv3fYC77SL50i
61mFnw0ZE3hORfAi0qhzJ7ALPDS8awZsU/yTVp9MOLzEVEZhuVnugjWVneqv+igryVyScvFKrq7B
WG7ZON2cE8wmbY7YOCjOJaIrEilyzFsw4JbJjBnftakQFOVpEkO6SJHgNPj2wbgYn9ydfz6g5Vwt
4aDYN+ia6ALxDg1Buujj14f3+WeRtokSV5qZ9LgBjhJZb0mdGXw2dx9f92sEIvoXtuWhVQVfVijw
9Go5VxagA71uHAmFkQLMEy60F1kJmOeppjsj2DNTn/6l5QwG8aAtAKDCBfoakEDdZ3/pjYW8PGMj
EGgxSa/9AQ74s+UU90765FDMVchcK8BHs3nLxUBI5sZUXSNLYePN9V5w3H8h4NMXwxauuyzA+qMG
ZdY2fybC/KMXoymqnhi7EpVlZY/T7Xe5Ofu9+xyfquMQGFIIGocn5wWN36xvEwlJGAnvnqbR1E5w
lFVPSQKuiWsAoACmPUI5XwV1H8SaYITsXARa9+v6OX9ZSdg9Ys1eeNUQZgC++n5bjGUdcAc1bnf+
WOjJVrtAqGUFGp/IxO/1XbTrCZLw4RVqCdJInuP1/cjE7fBNg4ATZHra0f9coi5TuJV7Skk6/2iV
ghGJPxPB2a09d0uA/WTrTA3HOdyboenF0hoEt1ckxIFV+X+LILFwZI/Dd1q7CL67ab7VHXoZPlce
+CmWnzf0O3sieUtob4azOpNK0+y0thBjhli5DMEwtI1cXxXjSmViBcNUbjenrC+i5++HV4vvb1Jc
OGGHWJIOM4iHV0xHRb4ye+ScCV7vP3nS1r6yXndIXIQvNU3n1JQpKH1m23bGksGujrnTQngmkUbd
kBDFd7CoWpGiwpoCchcN6a7nl2swstIHJKWP2sPZe/jlR/96bbxe1c+yW0HkFpp/5r7BLIoEb8L8
GbH7Rwh3oVol29vwszsjgX8fzrjv81lGmYZ6XpeGBiNl+m4w4+86j5Ry9cL1aFyLb5+4YR+qJ5QN
83llNOARhqw8EMfVqTUUW7tACbJOVnludb5i+KYPiat3SqyTD0MrD1zNOR0qYlQqxhJ0T8YeU77c
7ZN3ip/yYtFai+qrEHzEOHQZfJw8whwe5CaPME1C3Y/rOze2lH+Iim6/GKIn9mce/XWmNMObie5s
Cbc8crCW1gwghLteOtA2drcPxXnZAW3II5ZhLDD4siSaXCMKF3zk9GHMSZaKbUo0RklZFV6MS0Af
1BCUyPBUHckY1BAM5wbs7JbhjVuirNxpF+DHUkYldAbE5WVRCXL/tSBdpPLebRfk/lA4LHypXtLf
C2iIxdaN22QhxwHz81TdnmOKcRKiYlDY76b5IryAqrH/rjEWX+PJvayDMeuYgWkWW6JwjvgpT5d5
+I1aAFClYs7r9OK1mlnU6PN5QjkMa9g3G2dsLFiTtzVfXNPCSka8toLxyqXmNgXV0AtWhwmQTYzu
o5Zkoe9d/1lvM6YvuCJoJvfl8GSea++n62rGxvhIP/SKrFOeRUlyAw7iaSNdj3hClt7IkKDmZKaP
ffRyEqM0GqZGol0/wyf6gDnVaSwNKt73Q7//UplT7Vp3YqI/i694ZLT2haZOU0D4+Xa+zNGGlNy+
gwiFx4bENGPCnfbOA8suMzY5q65HstxtNamEj7tKV9fhfbn/kBi1+14NGxAGjbaW767A4xfoM4PG
rmXlYAEXbCZF/UzYO9qCfNF5H/NPlVZnXQ4rixWkyhKTl0l2YPWAdZfSlvEAidgMpj5jYfk7Z2wK
hI2/JwYaMNIGccJxNCP1QY1FVGhHjMVd5oSZWl30WgVlEpidPS1sbtVYuZH+MIuQC2Kllk21KSW9
1OTnmy4MjGkZKTdqvHfurNVUV8VH+ILQE88jt/i17oi0YMdybsYtXGLmAIx8RyHCKtqghVlSYR2U
tG7Xb1gKQlnR0967yUq6OQEZjw68wDvd5bWCO7LrTrWEQk4nEBBKHyPeCRp5KTP8vFwE6w8tdBhw
b87MlpblnPc3/cb5uoDeNAJJKM1ecKKjpEDOyr8jkS136Hpv4LHbDCKuBqEbKWxGIpMtNimaFfWd
JB7OaVdHuuV5q+O5LTl74r2aDP3a/Xhi0ntrX05aw3qkBnaoY9daEReGrRqEfBW5saUXsK2YUxVx
0WKkCOGR7dLv7rgpPUwrcNfHOxzAFNHh5vMQoHzTFlasAD1rDiVbgrCkev9w4cmHhJsN58Iu/tAu
JMMM27mhLyBqqapabRVqTv/+r33UrYh4yF7Lwvyme541ifQgkRgrZRGkEAEcS68oEfatQv4VrLOM
rij+C+0if8Ps1O68qsK1t3RTdRceyUegmUDk64eTSXU0QJ7caYKgJAbpZDOZZjZu7bhekMYSr2b+
yZ4E9NKUJ8gmTxKMUX1wYJNMg+9ClhhEbJHYr0lCQ8LFgofu3pzcyo5A08pQhLFlks/lhcVIZzLz
n5Ci6kDzs2tclmbsDDavkshdWb+2AusvDO24uwQw4begj3Mn3umVmJOWDift9V2uMj6aoHbtVlVF
ujqID9x75OgZHyxvMWfvyMfKpKVfu8BQGO4JRI83hoVAn4db8DjaIbZ6+tliN8iGdML7VdBEV0UK
Fy/WLhixnZH4EFt92lljjY5V/LB67CZiAksMD/DitCcu1oAZgSChNImZ/wPB7tG8CVukK9vAnsxp
7VmJQ2WfdZAd7J06inZIl4AqXyobVA/0sRRoLBl9xQO2nElgUFlcAdtlaGpb4FFDvRxsFE51gvqa
DghsNLRpbCcNWZEVL9fEfVOzk8Mhl/RkJFWNZcnDUjT4m9dxdyGXOdboKT8fs6VLs/sgFl9Epe+/
vtsOycDriOe7Gw1QS8j1idrPrIV/3F6HTtrS5l0hy5+TCLGN8vpUDGYzn/BRsvMaP/ie8ReKfE6g
Tu9SXcBFz+9+UOo9hJY3TqsWkeaCM5q5WB/NBWLUUXz/Wbpg997TJfOA2ujsBP9Cz6hOq6mSDEUD
ls5KVa8cVycD79YgU6JcXuB4aiDIyw53wJFW5ZJhnyNVf38LTeLeI1bNS66ChQQQjFKuwNqgE+3O
Qy9phphq7IV7QT7ib+zlrhvdpzq2okIf+Qo7+20KTAN/4iRRUyik+IXiUvnczqq8IPk4BOKdvrjX
EEIZP638I5N8e54/Vr2AOWjvVyZkYZg1v/pcIh5IzIX0FR3jbA9x2Aro/Sa0aapSDTVliUvsx2aa
9AtQDukyd4MRwWauxTQsZglWNovvqbCiD2SMnk+AA2XI+syyYhsbnIwmAXPNjMhGHbUtM0tbZKXQ
CUITyxKaaBDFwJdtgUhlF9IZ5hHp4eR6cGLB66V0Xhrsxqo8XbEZKvZBKTYYGYjejO8VvmIH1Itg
nWADhBKyNNgolK5AH2NBaL1aRK7cXx20S5DsYkctWeINz6suGmeY6pvUOSu5aS/5hly+UAeG1+JD
5ZhDbu7BOrhAXN2tEpXWAfu68rV0YoNglHuNjT/B/nMU64Q30rcqcURdkPZ24OQ9b+XB7oray5A+
jo6Hmm0Vpes6DANWWKQ7DzZy6KZjmRDMYVjz0P7Iu7n2AAveVQO2BpSeBqEhqoQfv8w9NLRO0itK
j1PkTnGItMm6VqXgnjXxQPKe3mN64Th7bURMDM5VrWgQsV+FEX2o4w68WRUj5bPDfhol9Fw7BYqc
2Mg3kNZVCXfZMMjL21icIe7KzpuPrOlBOxOIs4U0PLLzCOL0ackBT1VIEI/cx9pd8hrUAj4ZvV4U
Kdwn44IQUk0qqr0OtYVfpL7+K8bU7lHBbG6BynMYlhO4lRtIoNEFVVvNDig2ooArJV5hZhVRdWLY
mLix64aCnhMKc5HdxTPX5u+uWXiiIgo0HACO1wLGFr00LytwUATWdqDhPCnP6ymSZ9L9u4MCcqVI
Gvg5mpjY7ONK5wLu7CLASa/fn6awhIhlWISpdSM20RWrmNEznJ7nh/3xAq4h/RQvAuLUPcmt68Ye
zrW0mVRX4+LMFW2bGEUhQHVpwovWdjYpdUG4JAaZcvNy1w9/+cbRJR30ClT9TSoC8yqwTX38Joeu
qL+koDPE/Kkx8cK+nW2YAthOFo5Dcnav4ULuFsk9UtB/mqtOcOcv67oigavdAc0K6V+b/RO/RFaN
xWVkDqEoqHKZ6ofPNlPV0LbdA/qWbG7sZW32G7798NO1kpjrFW9e03GP8Z2T+HabBkVqh8satu8/
OZeflIyiN/fYJwyBZSy8PhQGC+jiURVNbWFZPU83C0oDtNJdgujfJXW9nxWTsFpFarVeKY7GMWHb
aIGuEIrxa0gSjuPx+xMM40IBG0DWK2pAwyCpgh2bNUcz9i+drtflnQ1KbeBPHKAmMdhRLohLSyo1
rzfOAm0BF67oL8e6Mx8Otfufj7NOeegWYsxKzjVyP0zvuJSsbuaqfQJ42p4f33cm12M9/x93QqNi
wHbNmEbn7fxD40k5gOoCp/s4Pjq/4k/Rg5FEaaKlY5GcIwE6DrwF7F8ZcYWNRbepGNyPtzEXRn1D
oRt5ZpFtYMv7O+Q0Gj+sCdszYBA5RhSPJzzqynTAWFetn6MYGqOiHtiRxBQlV+6YLWzuZxNNzjie
a+WVs6yoyCjNQ0geE0mXd4S4Y7zNIIZuEXZaBYEVpAJHXI895aJ15+3/C+anx839HodAmhY/8KNL
qZEVmsjXsdh4+U0DI252TbUeYU9B4C9r8LODYj9ddebPlF/YqyerLY3AsdnMMbNGqWxwlUODXDUM
IpweyqXkitSXtN8cDQ8vbzKk7q2gRfRYzRPYvkx3uScVjRWdJ//4OuHkQ7djhUrPZMIa3Gtw6eP6
BzNtLiezHqFK+w708zjaqumTJnnL+3J/gEWaBL6ZL92jvFpvRILnsNILsj+AU3Z8d/uz9T/hWELF
dpcqTpGaQYoTZKBmtLXvpXXxDLRMs0R4Zn7ktTMLbmWw7kIBe20o1fPxGuoIOFQZ76F0zF22ZHWE
T20AVWMoutBu2svia+hU18FSjr31X195mxtoYI1VNUGBiwL09zpcubY5CxeMes4GfLy9u9iKKex9
qu8JWboYJvqsnr5vnpQbEFnov4MLySeXN1pMgBuVkFffjFjLnLp7RljVx7HU/pzIcxxdcyb3Q4Dy
nFdo/16SNmpMAEEVHmXU3iGNiBHGEsYx74EiXC3CKUY7bEPhDdx1L2Pxk+rBAXSNGl45tI2PFrCk
jKPuENHh70ILiKHvt57UxUbFNpT8nUhJYG8H2th17fBJ3rwhSyALVf77/xBmpVdytgGrDXVE6lmE
Z/1AMdDFcUCQt/rIoGG4BndbfQNSHIh33lMKGnjZrqiSKgZKb9RWQ7rbnSHYpadN3VL5cSwBq6hz
aW3NHfOFgd/SZgVlBHphDehhNzX/UgABLXwQ94ZTaGgXT2DOakiRtrNh9aIaevLZauxL088fWNIK
+x0oZQQcE+a5WYKTXUw/b/FC2nWK2HjDLSkKnUmbf9fh8P0ZGhQywcNZa+OF9oDfH2oRcb11C2aX
FSmAkBwubyYC8H7OBHq0ow0R0mZ224MeOwW7NCHVIKS89+8miYXpf3sAkCeUzboChws7rVsJ4u3w
o0wqxx3m1AIN577LOp7jm1I+yELdf9+V3pHqDpZHg7pOzbNeDZLLpUVCpIlSNNh8SoFlEidL9PWX
AR+mGiWRQEwR/4jw9jX0UukQBB7KGrA/6ai9AtrrLtDhIICPgipd4xbzdYNnL1GptpHgStLnTqTN
gy6y33E7ETnzlg9bgwetLahEcRttRjaR+oDvFDuUe1SFhUqu3r1CJ8iq5dQGjXv/ES5831O5t+6p
ByWEuMctWOG5Ygz+JPOVrojmWtnhN/MjY5muPSXFJHn7qShRTxZBSe+ykUeo661dyGfqpIFNMA6S
ssS9E19DbdA7Fl8rnyLZJsEgvkTzRDo6eVc2T5/9qMK55bIzFxibpeg5I6Sk2x5ng7JefXLXKx+h
EEnn3ln+1v4QObrFIokDjE5OMb/4dPapw1e3mkx6tDdex9siQw4iqBZuTIGepHFmc1IjaUwW1nh5
v1rC5ZzAcUsKwH8GtiNbmOAHZp6tNc3Y2aGtWGCD5bHMNmVjk5BegxcMKRh2rBY8eeXVnIlg/bo1
3HVFOlG0YxAw1Jw8xGae+CvP8U10NFOvcmYKPnn4u0xlswR5Kja5cHICvM/Zh3nBqX8lWc8Iwb9n
2vc+hpI96KaAQVrKtdqcSwOdb4zYivATyTBHRZfHRHS4rm/AhfIgq7SO9C+7zcmd5SZ3gMVxjGAe
C6qNj/6koMACiWuy+KXkx7POy+eflrhc8v1Fm7piKxi4BBjx0jcmMluL5boTIbHCRhneyX2ugMt6
VkzI+vE6CYpVPx69GGvmyxuHuM13oiONmKz+P+w+Jl0z1mSPdlHHAFodDG5dyfR2fXaPnX/HfyLI
s7hNls0vJVI/2fXaLQsHg+qpIWYbia+VOLkdr5l8x+BLDzTFYDIkn5qAprEEOaU4OEue6MEZCWPB
wJTYe0TthSiGNM9r63t1VYDXOxiM/X+lY43YKSwNZWDRKU7Vvem3vHa1SlxmWplanuWpHM2ArYhX
ok3FZ96q4eJQlLgjLsd8qNRtgUnPJyD0CPiIl9zWIfNxmXdeMf7PD8VD98hdWIYMpMFOJ/2HtVve
2CwwKWCZqf/BqWFuGobQ6uU5KsjCXzcl1Wf0PLHcA4OypIWBvu0z2/XP+Ehcb2U+5sX2k94QG/s/
UZmvWouszAcyZSknmyaVxydZZYOKsGID3R4l0kVZ9522nioN0jdVxQ8vHX+vNB/qVavsUkYWM8S2
26JJLmMwFmjsJSzVK2uvOTo0oOCWjI/DxDxvLzEbr6Irw2IjIxGSBTiyLINwLjv1rrGQQ6Vl+cmC
c6SN0RB7sx2w7VboLJCmezRrIw10v02y0JNZ20V3oBzUOlVBBhZpyCRmmi8WEo3yH3f8vMPDa2Tv
vBXR+sVEKAYAvwoU3lGkrfrqajxUz15fPc1Eg36ufq0zhR8KMmnxucD16W6aUM74udHAFCfDhVzS
8/VNBGEv94mIWW0Kg6isj2UKgwpiu6bZuEAlZKuytWsMGkJvR456y+j/FhKEcy8Ypbn4WQKG8Lo0
2dK2lzxvrUXJSaNforYUPhejCQd63PzMGpRBBKAyCxF0jgIkJNS1vReYyqGtsoWjkF4x1TmJsqIS
fOyh737L/kYHNIpT7E+ZxKMAysjrQnfN8IqyqO2VJA4cjMPOlfGdJzhohm1hMwTBaw2paTR6M6JB
fN/t1TfZPkfqD5kOhBy//xsT+ClWCym1UVbsoOEFmlo3ErRyt/U/li9g/oJBXuDw9T52e3oqV+SD
8uzPMHV7wR9elgtqnb93j4tz2PP0l70hJhaIlBwY/fWtCZp84LoQRLIOspzdGey2p43h1yLVEHXJ
yfxTCOc+5OIHTEoF6+o7vNXMUUfmC+j6Rux8yK3uO/5FfCxSqSnItHdq4+kWMGBo8Ye/yBPqCeKV
YJdPjrRded8yDUzEysLTKa6XJ4T9g9GlKSlRL8NwTFzZuyRliWszNwg22nEZD/a9eoIB/9a9jVZP
dTYs3riLrpXciO1DPMadQHAIXppWOW4wsRUN3N3qgXdvjuCk9L5IO9fZNoIPahrpJba7N8Iyh+ut
RDMyn1XTBKJ9rfm5q1WnYYU0EFd9VnOVUaQNTT/FbQ1e83XGFPiRYrhrWINqh4qe8qnWWQSHlL76
gTsdIWXbjih3JQeyIwy45rBYvO0aM8L5aWV8bWn/+w6csQTdzZ11X/slyBxkcX6Z9LW+D516JKha
8c4UmpDLea+pw7hpiWXTkdvnHAPqvp/ZSZBK5SJBluPmcxfJALNH2li08OFJQPM3gEw0xROxjJY0
+DrMoXpVvwOrbb3iPWXH/Ae2PvTCV4brHLzB6wYeifhi3d+GAqR/w2HaboO1Njw0bYoPge5H4U7F
GgnwoF4g/KmWt28ml3Blpmx6EpO8pufbU7/KYHSR8xLapGMT0Mb1CGPopey/lqCgBKKIDplyFYPp
hcC+DXL/ZA9Cxt7vr1hwCGvJF1sLQMxtocNg5miWn+iQlA7k4gfl4HPvXxw5K3n1IiS6jpnGv0bt
w5TRtJ/WnT1vRAEGnhmxTv3CxHmf68Sx8AL+Km7696SMECq0k/Usk8ngh26PxrtEC5pvkBnWO1fE
ZFdEkpDKp/sXU/B754Eeon0VMnfADLfdTayTMpn2aVfEeu1g8m+nJVOtmAGyZWe4EMD+SbcD7Fbk
RqNot4qObK1cvjCTqgUp7v8svquLmCxmK78f72nm+QhxLmWLwqBPtjkvf5Z4Oa0YvxCYA0zxb1j1
uvXishlE5zcBQVOBrUGPqV4bGLQurWOkQlbJLCcgkQzryaZvSgxg3+jWWhE9ORwo1s8c6ei79m70
gOf0v7n2JtXe8oaRJQlAZon6JxI9kcsCjgQ0LMZlvsKddpLaqbsKa+He4bM1IOe2/Vye4D+sxUbg
Gjl31LTQRne+wCdBeDvVHhHBvVaQE3JM5Kv6bTGZTa63q2TlU4iicBtq1ptCv8KFNttNpGSXx3np
lnoTiV8ZuJBJkPH2bbHlH1XufBvK6I9ieGdVcZov//MhMKXfWiuX2zqTWr4dUGB7ttIP02gvN2xy
3A4CVc3BU30eSDkmKa/E5AkhiLvqiFgrrlccEaqXdbsRugEP3p3CEk7LQFPXC+Es6Pf44Ay2Hu0A
CSUzr/wlVB+1OKoBYaFdWfzfr3wS9COUX04i0tyqoN9Bm/BITKhi9IQvMr+CgBvRw/Z6XOiieDlV
iS2UDtxySxVI4sH9w6zLKi8TtDi4AXLMzer0HbcEvyfWxwMmajgM7huZ/Td7adzOJFT3iMS8JOSf
ojxrCPecANKtwSIp4YWSqng2iAsDn2Ow9IdjAWEUtgLUM60dgWX0a2h5pU1mHLvebo1uT2fUbYIk
okL2fjL63w72XlilcwrshbHGMh7qKwC9/mp1mxEqrYz4WM2VkK6Wsj6conGf3s2ORZFcm4TPdklD
teSu6FBgwQ8RnBd0JYvVkmHjQUv9iJkEq61oTfXrg+Vbuies0y6HExhbj5MnSFFq5lGwswjLQmmR
IAX75dQApeVJAqB44tPYkoJIJjwNKnn1f/tLjdYVjWBY5MTZQMYNg2nk8k0FxG7hyyUWporbuoTV
InDa/WJCEMdOqefPRCOAcDnQZ2iGngeLVPAj689yc4jziwus2jRu8qAnb9fe3eXQy+mxOnz64phe
E2dah/H1XdTLHicpDKPwwhkDsR9Z9rn+Xitgtyq7KeGAD0WuscxzzWSxoZOwhRRmCCKFLxRJhytJ
Y2lRRTXegAwGT99QoQrl6YpKNmNIV7j0lB7ss47dW45JUVDVWXXRYa9hQoYJDIkD++3p/950bAY1
fV69u/wu2v1fjucdIK5UZ7RO+SzE3L4IxBgD+KK02Wfb25Nrgm3MlWdZXmxyHy2fXqIh6dwhPtvu
zKHyJ+TDcQgPUo1zbnIp3CaPurLA+VA1y3ZGI2sEld/0lu9BKEKm+GPYNkX82TgUP9JrITuEHQnp
r+awOhinoWW3tcKmVkD6mxg8uhJHZUw+LEBYounvVWY8ugPAnWrcW/OAUsRqRTEpjvcdRH2DT2In
PgNX0xiQtgCTTcmVqPwyQVfAS4wV5cF6wDhP1RBvjQjfKN+N0PU3hUm+3mvuJvt3lCBPqz+OmkoA
T8/fOMG9M4gD73qcxVRY/z6rufla6+QXGGnT9Jyih9QkJMoNQus49ClkVCTnYRmN7Gxf9lF7l+Df
XwN3sjo6Lf3Amju86WZVe90ed3/A//cYM2+YRont36kTA6GwBEx8VE3fFhdTVndCyymYUYs8hObq
unRUw9jJq1Td65H94LeVMs1YEmE0smRI3AefL6y8i1hy3awFPAGsGa/rsY+fK+zEoCjDZ7uHu6tW
bypb115sWqEec08ropjzhonB6KLGJtjprRvPxnat9pvnQa7KuMRJmn6rBAzQeF35Ptn8w2zPFvH9
Nbuxa9dgq4xWkKGki2VCakpGaFe9DvGnN/EPzC++nm6RnuEep2Omv1ZUEFWEjUY1bVV6EDsElHmP
O/Xj1ipEgk5IVygSO7HZaU7lWFxLeqXWfZNY36QdZvjQ8t43BLZZxC/AQjVZRw6pxakzbF9T0nVu
xZGugeyvTOIsoZlhuqUWXdljFzu70E5opFStQSeGipNXDsQYMs6qmwBwiBPIG9z2QM9QJf2w5G8i
0Sv8G4yABbAXme7YSXkViydck9dD0EpKSSy98O748FIAO96J/v6J1RdcGcomZgA+xvtEIMvNkSjc
h5t/LckJeDZuCs2bbQv00AiM95On0z0qf9EALbqc3l3EI14QEq9CyV4nzhdL+3vbI6/8g53lrVTw
M4dZsS8sqQlCzfNVKW5ftDBC8LJBqolFwwW1jrisZSnEV4keqxLu0TsQUG0XkpFmC8zBk+L2rSDc
kC+7byDn60lKiANkAuP6r61sXQet9DxACFSsVZSCMkcn90h/j/JrjSYYrAf/FQUm7vmAQWk6+T3d
tM17w6bjCakXFaNFlI3/O9RJIwWFN04Vvt2wKzcuCVGaR+ZarkydYlDFiZduXpIdtjy85Bs57df2
DWi0i8YBplgpgIC1e75Fp3fYmnpldxg7dYKYaWsYfyBF4/3p2SqhZaztDrLnL75izcAXSPORelAe
Z0UjcvFxRHNvvdOvonZs1LW6CO7HCFAq357FrE5l/N7ShB3zDYjthvQk/R8PWppAkArx2AyHy2lF
aCrnVvPesRRcaZtBsc+0DUdqlJMho5dfoKWr35dRX10Sh+dBchJDS55yQKM+0l6MM1uSkr1uOPmw
ozxcLUeZZ26UtmdoWK5hVFPYbwXuXvYFJM7SuIQ3iEa/tjm0lPnuCjl+bNQtkP7Zj0l5l5I9yE57
9Uqo9AiVS+veiurLiYKOaPKpiJLz+1Sty073d8fgwQNXPMsnWI+CgSQw8De0c3CXOqq2djFIJmrx
XFmqw3XxnxmKI0x2hF3jYufaqV4aAL+Aj0XPSQVREYjBo+PNs2uAWTbQu94/qPaKqdppOFr5oWjM
ofDOqU8lN4ewmvjwDRj6z3rHxIDdafybbLHsyV3+yv6pD6F0rZNzd/WSgwW8SSDtoasN0/xWNIkp
yOV79jGYHvFqmld1F3k7JFM3tyUGGWQsDsHJ2XThfAXCYl2JWGC7Blxtiwt6vDpZ2qf0o9F14N8L
NRolkpENn9xnNQ2sjyXk0NwH23NqOZrO4+Drc/pc5wgpGRqDjcHVRapBZ30kGS9LgSu+7EZaZjX+
IsbIVKyICiXOFJ9zZ0sxp9z6dF2KuH8pFag0QEFLBkRyg4J7UvrttzUeZTmA994coJaglMDtXgGF
rQ3lL7R7ugF/GdnIbiGexU5kI4AQ+q+hl/KgIX0Lm1es800jb6cz4C2lKAYGoAlAYd+UiFqKWT/F
BBp4prTVJ0u5PC71rbvbzkRP8x/Q0YLrOpAdqDn39VhOvs05NbD4KyfmkdDivtPnV8e3jSYsb/Cn
CfUjauYuAU1KK2PwVW13rCM6Fk54pYnQ51syG3t6Tt1h0DhZp84IVg+TpJwBneDukrYi4LNuqAXP
YOzL86O769XBYm4cfMpnWLruyBvH/gR6ETm1JYHZ9c/uHx4NTXEP0/WLV2mXGTjkrRo4upDxbW8H
EfZ9cbE+/DXDKUWLemzmI8g0xtbKow/l5Yj3NZTLk0gJo+LEiB2QAkL3NQSa5oJs5emgX5AIPrSK
6gm0ifUIRl1c1IuK+X/JBSnK3q82VSPXg+a7+pNo8cbaiKL6qGOGkcaQW9esbucrwxAS3vKiHCBy
mUBWi3UV8jc1XatxgXxxtBt9fukOGZCeaj5HMXd4Ev4gU8d4fik811LpLFX1IgEGOg2ncBHu0rXG
h6vu35ceb7qFiJWdBaA619QArg/bRLEYXEx80dfbqcw62ADX0AyHzxuLMsWWrveeqH5dHz1c0rPx
e/omjjAx5am0nyXv24APG0e3gJP63D6sQ11LR0O8o1MsqPtLbTvJKlyQDzNX6gICR7pLSDYJXHgQ
1Xe/+R1rslMFvHaaTX5rd+nnS4EJf4DVzF+omwIkO/55tp0cC3DkADk/zBSSjzAG49KFfN6dUBIs
z3S0JSmooFaf3GcOgog42MiDDtfLESCLPi4gxLFYS6019aFU8yT9iLL9i6wuLkNBxo4pKzflpSMq
Cg8co8oYwyyZMdNTUm7bnoTAsHxzRp6PUWiX4wJVySoMB2Tt17uTNzQ0/XIe/IWlOQ/3IjZvOPTN
gB7xffWV6jxNJeQ89cdAa49ZebR92J7WSkfiwHNu9lJyj4NY2/OCnmUvFzc3MhTrQvZ/UgFcMro8
BtT2SNEc2FbQbS38nHS6PJtQB4zVwe85ix11fBfH3XDg3tGUwnyJcmqJdhYRpDO0q2JTjliW0nS3
h6WzqbwkLxQ9e7ZZX7GXvzFBEyVDtZZ3nyqExFOOgHZU3TRXbzuj3ZPf4g1Xm++6+wrxHCmpQuRW
UGlpqSMpTGueICwEOb0KaFXJTcF4gn+VAOqCsPmxQ2N0krT8urYk93WQ2489khI8jRWinH0/WbGD
kpSmF11a+8sWzdaeaEHDatoKY49CRLZZxtrdltEi1Q9/qzkPKsSTZdKUX6MXsfzx/jo3vt2O3x1Y
NcGrrS18O7GDKLzIwBkkzTef+AZhelvtXTLg5ajhCMlWxLRIByqcPMIg7MF+w3E8xGYlLA+KgxE1
IgTmklXyOwDaGz3Oiw+i4bXBl8e9LX8uk67tVTys3+Wt9pzeOx5kUjaycEvxi6OQLGlWgIuz2Zv7
w0If3863U31X/ebmeLfoPvEj2vhKmUH9TSeJ3CVcIDVNeIg3murp4aOsswlCbjqtDoCpMjoDVeO6
loWyi4BmMyysee3doNDCRI3SEaSc8ol4CPRfCWzhvqhFe8VBYSsOC1zlKBDy6b/HqBrk1DCJAVwG
kf7OHSlTDbcLZv1HIPQCsd+N7PvlOuM0g4SaL7sj6glKEgzhmNB/kXKVatRs1h43Zb5F4Gx9Thy1
hYS/0cpjdkMVsggs4wZw/JQGSHVaWwL5J1eNidhvUGGyZyx4uVFAVZHSjU9QB+NDobBLriiFXANh
A2Wvc9qIJwGMb7KV0U4PqeB9eOThImPoNp/4sMzPS4DoSZActad1mDggXLy1Rx+2dhhHeBy56SRd
vK86E1v59D+oBvscpGhydzKZK8noPy30dlqpFyzrYbHhlg7NlfpNII5JP+EYEssRT2JBSCIIf7Xk
YtpgGFy6bDkUNP62NHtRMt76cDMC8qNNEDFbON3jkxitnLmns3ZJvipOYjXBi00oxk0lTMBt3ne9
JN06PRvywWULxdD/GhOjBcQGLP+KjjAT0Zsw0gpjqE3lHoXmC0S+BBoN23exa1kfWzd38Fkf0Dc7
PbxEtt1kdN8an7OtRvE0yTTr2Hq0BAzu6Zch6EIclulWdbEMdzRCermmSE06LNzsv4x/Pgeag/Zu
FjhLqtVluqwXkq0qJgwQQW98BFL25LaOA7G6/uSMFcPfH3/EYJQf+4KaLcv3H1SEl9u2zOSX98yK
j9T+RNbSMwtbHmYyteFnBQkXvamuaDpRLZi/gYQBhM8YqUm8EGS8Otr84j3wMoGquOCkSeuA+ojD
D3Cb2uiF5BuKfgPiTGXrYd4wSrWAU9Fd1Wj22RI7g+l0ozzyReYWgKlDIEWQqDqr5e1NMenWqXt+
h3j9EwDKVKYuRshgRIXDUhHa6OeYT1YAkIP/yD3oARKP5W8ReoeD1Wi0Tk/5UxB2QEdvXUYowH6t
BwxRzZsSsNLRiycdA73gAAUfSZj19hiRNlsXA66RXzXXWoLzop6fsRlOsaQ6r89gyLEMiNFKmuUI
QqKQzjaGJnBWL7yYWTUzQq7wEZU/hAYUs3UWblhiatxtAeoG37GUSqEzibk502I6G4sEiTTKg9O3
c+nfmqj8YJQ0kQzBUPhfq7SFlrnHrBRX7PiOJD088hhOjNFlNozN/QOVDPvJ7vk6jfLLuMAU0zSb
M3nntPVpMkKUbldZ5+f1pwi5eEQqgfHyU8Qpq8QOjCiUSdEo2/zZo3TZXQsqdgZa3b5rC9lM71yP
1CPtz77FhURQFwMhdyd0r1JnOZWL7TFuCDAdZjHL78NSjUGG31XPzuvGTtNQiXA2vwzoikSYcEkP
X5kt1h+XtHnwYiIGn3Kff/BPQJuQ+pdwr5oxHvX/BHShL0fu+k8rL9m6norEfT6+LkP/2qPrcvZ9
ZeqYVkU86E2/Y60Dn3rTHx+7qx55+kfoqTH4LyqceDu/YPK+SCcdyTTPwtDof+V9FftIA6vx/TVH
Mr7bQsQGNPVbPyqOOl2/CIoUMPBJUu2UVkMg2LqIQtqpl7opp8oyewFYhfVzh2nKRfWX4tJ3XRI4
1XZeNeRHLVfvV7baqGZHVZyOAQR/KRVhZg6UN+dXaXDQQoLxn/poxXJ6BCEkb2ichv7j+UH9fxyq
We87p1CJ89ASYB72MjPjuPLp4CSC9x2iKAub44BrAaBsnNbWO/TR+oU4IEHPufxJNgSgWEk9BvMu
pHRtG/xC8IjetYOnFTkS+poZx2rtCO1d6pio/jecQkq+fp9KnyCyipHXNl4Pg0y+2lYr1e4Q+4PJ
tKYORr2HF3bJdw9qTs6Dh5q0oe12sdMVCd1pR0dmmQ7QtgZsH6PITiTB5n1SFBKKuZLvYzUA02nV
gVCSigdVb60HQ3OdNZcpbM/bWdtrIDL1LApvkT4Ivl0DVpOtVPokg7RyCCsHLylffyRuYiCKMVZF
lZpV+Sary37dCS2yNq4rQtwFowzdmJzzRk3O/pffi+FhLRp5nqonFnMa1tAsJW6buepzIt0ZKo/F
WZU0HabmUbcntzBW/xxHnhdWfBD+0Xni7e+30NLBf73QHxPmS00DyJ38joEqfI9gRLHItnoPKlLO
qP79hHwgJBvFawGTlUXoyOkj5c9JjVVJpIbyNhgaqxkmjjUiOvRf90QwrnTShAWc77Dq9Dy6rndU
XAxYbByrQ7bQDI71FhlRgVM8eL7Rz8P0m66iVIHWPBTn5yuNhdK68WPyheb8xKk8lErws2RZrk4a
J30upE3wTSp3Iw0+lwyyu3j2PkyaUEhlDQ7OVFkY8faX1FVi+zzqL0R7/Z3xRsnFjItcFL1CYlLL
UcGsOx/T4bFKjDOEZJ1l77z3WfVpN7x+GhYogfL9WlSg8I9YetB2vemib486/XpQ3y+Q9Ce/arAw
2FKdGcgovyh45wPREHZz2rrsILidY602p1C3e/lqrzlSe7YuyaESvCJX1DGaa3CO9fzIBpWHVXFQ
8Y1jv5qQDOHpOXwK+2sfc67vF7Gc2JpTI646QP93vhCJ2V7Hb6z4774Y+3jAMsFs+Vdf8tRzIIbu
4kJztuwOC/RPKjmoDr0O3S1qOCr6HItFF8TAlCCacU1TANwjZQDH5lmG2aFf4T3JUDqywwBh67M8
mzZIbjkoDAonImNiRwlxAgziVTQgunGo+eo4yIwxM9BFAi3jpvHo2EsGUwmLqW0prgpwHClG043Q
RNg5TNhFT80guHGjK7H1yQluZsui5GuuWUl2Ld3ixxP4Be1+wU/c4XrRcrj5TEHZ3IjEmrZ0kl9q
l9iQku/+rE93P4TGajmQ1zN85MpICRZXtwxUoYTPpx/Gldv8/y7dCivaQjDVPEHpPMQblFndBZk/
Erjko4RTSezUMiaiXpP/XjPEX9nNM8TTgRzX/mSz75BEZ0RDYJPtvmBtwUd42hE5e6K8Osrt53lA
OgmZkVHyzMJ3P4ive8w2Sl2BW8PqF9L38am/w/5+41ririuZTw6V8vwbRgVAlkr4G+nj1CkyfGvV
50tmzbhpoNwUIw/IHojHYPDF43C6iR7pgRxSovGXCr79GeehKGLD5mNQelOghqdklM4TwiR+TOja
881YXHKJx7GebiLdHb0/trPaFYPdtkX9a8rXjSAcxO/65UBmV4pK4Fsb+/OQYj9xofScfg0vqiEi
gf1zhLm/KOtWOyrfsALQaW80TTpwWTp3A0tWAS6ywCgO93/fo/ZkOc+lCc5by7Dg/t4v+gdFwqnE
rBya/Ki3eOO5eGmuVDtaSb8jufxzuQSO1solk4/B9yBi0OAjOGMLF9N5r2grN+OvodYyFZolHkdw
SOChoMRPO80PWb/OqCUrTQtxC3HgLk94+J4Aftc0jZJcDlwLeO/s+pfg5jiKDa+ejE/29wEgAmYX
pCBGbVnvN1oQRCbKVxlEDrSk1fX2RNbj6iPLtwCqzgx5ZPG4pDKirYV2NBvZZxPasdyZFLHHqe2H
xkmudAa+VeXpZZflKcLD4TQYh7Pm/Wq0EgmD3HOks4fCs7LD/ItPNOCKzU7QATION7V8laCo9ixP
dS3PeGX0R25Tne6qiqGY1Qa+gTfVXnH8oPaJShTpvsc/F58sFu+o0WvRqUo33OJvU4NXotMeqLG+
j7C1kLeEfvCoz5FvwaB1n3fVBpeFsXPdRct5YeR6m2rMRnQSV47r72wKRfh4fN6FCo47QQvxZN45
adU9fLyaXPAbltLO8AVrBLS+mc0hfBhSiN4pg20A3O6snMjMBrWm2uJigOS4ePdSXutyKRYqkyeJ
XSm8Cm9MnuFo/YMPmlQ6PtkPkRZPShfdbxr5HwhyO6gzltyIjarS1LE8p948C7absCnQxge4Cv15
81IAK9/oka7Srpl1HHJrGTdzw16F9dGzS8PjVXwcy+qk9ppLSPHiQ+pzjRvT5UW/Yg4wx4a+HD+6
V2ZvnDBMg3TyTKZdyfxKsVv31cE0RgGaJw/FTokNAu6aXXd1B+Hg9fW44c1HUxtFdsnug+uxU5KQ
44QBbbXyRhkYNKV4fRnsY0oRdimuLruv18Hv9/kCCv4u/BPbwu9Zh7aECXT7YFdX1W/QUU94dtAx
R+7ZyFX5ReZM61IdA5wQqwS9pB9WQrXv2DWPaBTbBAjLc/imGgWzOUkdVG/ijfiQCUJEuC3m3lb0
0lHIpItreyK5ifJbIETTThe6hcS1Mn4U+HWc8wLL+4d65/x7pF4J0/YmXy44XRAbGtjsMVo+/sIz
HmYmDhGnz64G1CxB9LhNcu2kkVuFT9OK75iEsOAH3Xk+L67Z3sjmZBFOXjFdT1iUmbh+Dz+dS3lq
ysz7kRGqZkXtClK2Yq+8ZtGDnCD22zoUfJ+/th5aMEwBSocbaz7lecENao6ynSH79L5KA4bSyWiB
HMo7C90YhSyWGUT5lOb01TaJ/NH2SayZEXbRaksg8DNhPzTRjrviPIMGTEYKlJnKaFvx1902DRgb
DEj9A+YZ81ksSSEtjdN+kJ8Vzk9xt8M9uTG2bAP+pXIe04sIrvpWWVU9a6PGBvSB4atnLNDkmYGB
dxR03huOUPu8slwsQ8iEYgZjmlowMHVaJtSMYQ0xFr1HvckBHaLLyl2uhD0x0ps1HDt2gdhHg/Sl
fQu/8N56448TiNMWkmM97yMcfAFcBqooTU2hVSq6NrP/fRkN3mEd13omj2MisQibDZY06wl77i/q
3hTSfGRY0VOs5shgFFruqlmSlBvGkYrClfyP6yWtc9XswOKPabHI5TSNiZSKMu025UeiYkrleycO
mimLqfHCymXJXBETHNx3KLyuC4WXQAhdy8dy/EgBkndZNg2tTGcvD0q7zsK7vfn1N5vW23QXuoIy
PL2pZ7Nmg1RuwKS6kWNcO5OFVy6sAkZJLLO2Oqa9M8LYiULRCQrA1FkYrBdoTMHtTFekil1PWcGI
sypEGQahscF4ATYx4pbMHMcf0qwz+8cj1ZeeWnCHcJwdI9Nd+UAPLHW1roeWpElGPIob6dqflCkD
k0l846PJ/zCdcMd3s/kLVonQTuaP4sot7C8rTXEaEMUMgODx880uQo3o8V6XaRKDp8us7RoGVsId
1lEAtTrvA+QAvChaks39IAaHn4GTgVHQCUYZcdPttkrigG/Npp7rjXFFYPe/T7SRXiO2ZZcxRD82
6z8K5Q56mBN+8jbr8xVuA7nfydFQKnKbFKgKBWFLbm2J7c9q8qnYNqYLdaX39LbL6SKTegsh6d/c
tkmHT3D5q6YpQEkAS+B/rF5u2dd0eJL7w5Elp5uzE3xWbBUJUhrTpPS5ZTb9YtqaMHK+2nH1chCm
DDOPDVh4QtUbcjkSLYCvsCqp5OEAneGOtnXrJkQ6hLnjQNpj2R+LtaPkcqJYenSdrhiqXOjsryuB
mWUOnKpdU96KSyK9EnLTt5sVWPvwu7HslCPqn8kOu0FdR0S9ljhpm7xgCk4s73hrDGh44zylY1nq
ilKN1VKuwZ4mI+zMiKRawcXl2oC7gAwd0OFcOVEnE4UcVxNuJuHtRye+U3MczFkrLJ47AgarbE7V
luShnypV0MzFBlOFlLQYZg+RlVi/j+Rr5Y2Ct8tUIaG2myZC4Rz8hCYwCred5j6tqZGRr8cUzpxs
zr0WILAe8rbWBw07xWd6pDzaJdnkBDDcfOHO+tI7xEfkQHJFPKovBSwJQ12GWk1C13YY3ZOZ8rLK
tNU7KQbngc7piTI3c1ujmNwWJqu+43s6E+Us0cf0F2YWC4V6cNgdzW5e0f7BNEK2gk12S5lidHVH
PRsT4B6pufmuu7xtAMnLxUDRypduSUM+SmbfmeuyIBDhLV6ygcIuNCdg1P3ikBuVzCb4nW3a2fvG
lhvdugvoYpYxcK9xxtxCEbOuwFEi+Wez5BZuv9nnLuhxw1PSkzOX3ck8X09LEFZbc55jr/O6fz4P
QY/rf5M1dlztIWYIwZqlybBT1+0UeDLLUW5+f/Tt5dAbg6FGVhPqOPXsBNX0nYtwHXsK/dMM9/Gd
bnA4RwZccp5ICa8DgHndobonRZfLl0bdcZN0g2wGOn5jZ6L2vjpKJV2Bwa/oRBeGWs/8SFDmsc0K
99gbEBI85FUdfcSQB66EiJduXAYdecVC4oPZlgYzgCH9Uzr8fesG3EaDq5S04xLnqmdtDQcqmoD1
enrKay0gZh6cPGKRSnLa01PuZNzMUeBAG0Nbce9RNiIRE6iI8aULzF1HqTEFFdUP1ZeXk3GVUivW
yEGC1nsuMZ3+FUGMTHx6c0dmjZIvmOfrtsJkI25pEmng41uii4LYmK/IEGOrol11nN0xNIXdJC93
Jxar/bvIhIX1Cinsrci0UuuVwcSGMpwUQcOkRqH4Xz3Oc5aHYd5xYjxCUqDjYPMNStIwLGNMknjF
4HFioqgMF9+LMQ7L2abhKdqIKTzHFvzlsqiLny924ZH1o7iPknaoDuKrqh1OB2jQiQcEH0sHZHvi
CknwAPMPSBIdoSkJgofR0uNYq6LqjntvCg+PBltJ/UigVuObku7PiD4ThJre0Z8IA0TugxT9L+3t
g2tXoofo/qkmmcnKqLLaspvJNOn1DAK0NARp9cnOqlrmqg8U3sIN0UWRViWcAw/HpA2CLMCE+tsF
xmfsyIRZozjhi5B5mmZCRgerZcFVFj1AcMEKR5BUig2IH3kmiQSsyVE037K8PmauKdHW5DoYeBfd
ABwsBzhcJbm+7DCUV41TCwlNOcJ+tLbMOXLhxpQh3QQZwpPxqac19H3GUrjc9dAZXRa+qrullrpz
OyjNadKyWIhDaY1ZLN9I/tEmGVh1H3+fjPgDTm1k9n1BHbQ1wZZeDhkLiRC94fJPc7g7qJgk/meN
8H/EZ4/RlcGjKrrtJ9qUEMyCzT9t/7PmLRkBq5FYmIlu0zMNZVw8jdR7fF64YUlGer+hQIHCQMTa
+fto8PLcT0laYfXHcnfD8p2aUN6/ZB9P87MS193yVEqlW+7AXsZ739p7XWfE0nV4wDRHX5W0gWXD
EeV1UfLIwz9gvDvSMBSyHv/NZFn8RUkJ72Zj1dtpnZpwMBBXv9h2RbmjlIYe/WQLLHAHCnXd1KKl
Y7ETxKHtSD3MnTz4x8EPH16VjUTgpo/+8Z0kTJdg3YEk6rRyDabTa5xjnmSnvetln9uxUztQo9jH
Z5joIUCrTj5HZFkHB+ktdEQzVUZnhYzYlmmk3lkrbMOWzDo3h8ZJBQ9T0pu0aGYK3KWHAtjNK3DZ
IF2dk6yBXOvB2wYCq5XDnprU/lq0p5bSaQ2dHGAdZthzvnGNr7uFvNG8dtlQrz3n4oQQItBtceNo
I/Q4ChJn1HstThV03ObLlz3KC/2esNQPyH/9y+TqW8CFU0cXWZoTAmdeSXdEVwf985itn56TgTv5
TevSrapPejEuZBQhpY5OUt2yxOZI/5Vmlm3yrN6Ns40L/nn83im5RF4ahAQukXn5fIqG0iXn9Tb7
UmRKA1ylBNbLGB/Blru6wt+lE79hwEYqUULxCVfjX1vbcd4N4VUoJzR0KWZ8QPmv2fKk7yabwZJp
xZXGo0r9KPnKhgx3rzvrqo+VaQnPuuHJZQHl69VCA+KvLj2OJW5igS35Ecxmc0jLPkLiD2R6nx79
gm1DuWkEb2Fw40PG1z1Pjs/mRNgXaZDBKNFerestFFdKXDryKuYMc5peWQaW9zD3v5lTuUTuA43G
TSG8frmSuzzwgOXvcD7wzDt02qnZvsivFgcuCUje4KMgEe4+Lc9iCHpq7pNI5udl+3wJRAdLyTJ6
X3QixulwoESXwczwyLeh5yYzdL28D4wmkSyQJD4dPUkwHSe6VSGk1HRZVuw9nhqYedSbSO40dElx
MBW9uPVylFzwAPHzbT9SNbdnnopX3+ZIE4KlRKBj3vGhjzskFm3XtYV6WGHDsqRP3fcD8D+3PdPZ
YRpbm/iY3c5p4sEyUKzKb1jq9J/Qtri0HZsjBSNdQcZ8DUq2aydKaol5epCBiw/aoCofP4PgAjJe
eS1cyv3u6mfDZ+Y43ILtLGO3JB5IiuNywfr4fiMLtd2lUnMwh0E0QoScOEcVWuEOfrLVf81Emfr8
X1Y7stLei5FDCIB22C+M1zyUjJH+e9Gj0R40CsQJOfHzNoreP8oKZweo7x4xiICy9FGDBWeaG2ry
OJOYYeiDz9Hr/iSrRMGGgR1fnANbVvXG4z9sgtFvOTziQ+dPA++6ao4+niw+8gjgBQ6egLLTLK9U
FCPzWbVr18rFKL9jtLt53IddHpeNNhnrR0qAS4ELRZtQWY2sh/HiCp8LuW77S1qVrCp2h6PckGy9
CHih1tWzxJ3tdXFi4ELZVNsva+grdNHEevhagjHJeCuvHHyjV5lfmr/eTpZlRFTYNsbKsFQexIMC
LDBbKqdjs5mHJ6nHEnwtZZo3HvFY9UPaAtvcJzAcbfbeuho6RRhrHtQb8XvlcGDv3OQX0N/3TuIr
Vv9XW7VnIZwRmuSfDygfH4zCTw/zox43qr9YTgQGw0htSG08pUwbYbmDDfG7xSAXrmjxtivUzv7P
Qi6YgxCnVGdMm3XAB2eVS9racLJiX0DTmBeV/Rg5Is8K5g3ZUCNZiNgcIBhQ38JKH4kjf9V/8ugw
z/qPAoBwvP+KS8vzQFUVOh6ADG260ijLKFmcXjdolKWTAF1LNKBNW0IlRG7qCLIyF7elS5f+vceW
e3pneTzNHFeQ3GXhqimfPiMNDHVcFQ8V1psMtkPcXbIIVtTjqujek3k7lR+k65AV43ha88e0oYTc
8PB7ah6W3BiZTTkBZgSfljAH6IBd9GVLDE9OAVgFUM3LiuBJFaUN6PnRlbhYuFMEuG5lzUK98KsW
jBXscp3VtUS4fUuVA4WHQYUVRRCaS0HzVw3SAFoVfzPS14P4zxbtGl3039E+AxgnZgZ3vgm/uNrR
Niwsm1HKpW80KSNo1+witPUcRWALPpJOCZ3lK99Ldn4eugUG4MBD1fSVTBvDIfserTKjchzNJuUP
ICHfs+6W3QSGUTwwsAGXErcSg98iDDq7jZN3KJszJVpz3Hkc+W3lBCBJGsagV5jA+xuN3G82ukLj
E4NajV1pBOeqXwCY7YAQ8WlpiwCJuQtM1sKiS5T/sIpjsuTTRMGq90V70SqXSMl/KJbUExrLAV3o
OAtWwjUQogyId9m1Aa0Sk3lULpoUMHlt96xqzKEErUruwWyNt46IOUc/a+3dJbOS7lEQOvlFYXYG
S9UZOwWkztdlo6ZK7SviPMAwMI5W3mTySqAwDGRCuq05l5MrkEl9WvN1vnv2Z40cBHq4TwCoJOFy
0us5wEIL2FTi5YGVz7yM/gMGfTDd5CC5+ymXgvgtgM/4LS0RrBxFD4SDIwz2XI+TxenrDjXxljpJ
L2feqHD04C3OSuYqF8TqwpQ+TEZSCUx+gcoTpdsiOU2X28KPo6NA0wHOjCZk4qBdcv088A9Pwiti
Q+K+yOvTZ5MKiYLAos7XmJf7t+O1ChYoZrBDJ0uUPEoYEEKqgU5fCzPvxr1SQoeMjPk9s9Ca/bma
4AbOW7E/9njAoySlAsrdgj3Gc+4jccMMlvUiyWaRcPenTIU8P2GhJdK07wY89Cp7Hxft5nr3sh3b
ZxEGcOLZTX69NQFs29/bE6D8QKLQqJckwP4rDVDElAROnjUP3WyUcpmuD795oiYmPJpYEqtLHrlT
o3b2m43kxzm1UF9SRShbsS+3jKi1IdhBnOUROn615npy/oN6kJJ1/HvowdCA6epzYb8wwghMr8Mf
IeV/50lQ+vEjnS2i38FBKdgb7mHLYrfKWYw0epFEU+i+STSClVZVff1Vzq6fKC32WGjBEA1Br1Lp
L4ZCzqv9SaDBJXXm3sITacA7oK8AQ5wLiahUAVSHU1YlqSdUJb8JmnSoyaaLfRdzsbJXqD9HeVMC
RhAJgArxyR3miuxMDPBK2SLXS1U0KvWDLEfUN9lJyMef3vBuJ5A55a1Uk/LdfZ+1Gd6oSO3kRGzV
8EzLPkfgG59bwmhKHNnsXSyNtt9smS69s16W3BndoVk60h9etb/Gdzvuk/Rhm0mfDvsFWqEigtu8
suPSdXmtVkn6Jg9TBVABBkbWvwQj2xdf2M+VEEl5d9NVSMR99BTRzb//AeeUL+ywPQL8S93sFsPf
TItF1fKemO6WgHwO3WtMHhBcGjtNFpQBknDgCooGoV8MdRCMAitBKfw6R549SgLN8p7j8ufe3JRr
aUjvSvdHGckAo4SELkcplCsMDX8oIZ7LakEoWjuJd3kI/wylLOXG6K+C2I+Wsh0IojbwoCA4IkSt
fNUxl9p8AQF1gus0QaPwH5oJGToXtXChN8lKKkWW4u5U7r5aKXkvqUytmyNtuSM5n/WXSR4lAPmk
1iGY8dmWgqDEjFltYK2T5JSbEwQrXappGcc3YwwOgwoivKVzTuzKNidjVoWSrdCR+GidK9mO1tCe
+Hch+V9x4jJrbNCEayuMS61DuqBN+2euNIsL05ZjOjGiHvlacy/C9KOFAup5xUFnZlKUU67OuCMW
aqq4aMN9hZg5eq/mm8pc3ci0TPCvU9G20QHLOcucy2TcJWlrcKVoiUpPqubu/pEjdk6tE0sxtO4w
KoXfiAZzhh1iApMdX55Z9ZlOucvE+OtkGj5kRo6UWGUKcSY7cJM6g5OM721e5+tVRfddx6cMyiaC
Q7IqPz7x7QLK+UXWNirKryy2Auv7LrtWkA7Q/UJUq81T8PkjnIr6ArWOKTpUeE/e7iMx7k9JYf4+
boQj6HZwOyn2j0IXyszvpqbIgITLozCjceBQSuHOMFbs7fo9gdFN5cYKdSVZxT8c/e8uQkB9iqGV
jnxXnQHuEYAgKq/DNThu3cmWkwyAZHXJL/kF0tnNrJwDsBNpBENxGqA6COEc9Ov4HSF4Nq9S30x+
Yg/h69qEOXdNhaDriAiqYxXjDKH1xCBX5oqpSzn/H7Xy1cWXXEyhKmwei4B5hdw1GnJNMrE79cU9
N5aQSQj6dfy2m/Mn4VthwsYUlLZabZTFBiIwUYYxU45hkqWv99poMCHZxISPvOeGKzwR9hm9uh6H
MtfX2sjF6CAo5JDHZKBE7tu21BpGTWcRGAdqn2fo5+Oxx9ayB6VaCzHoGy/2tNHUuyYn835sLEC3
kobQ+PHB5cO4L9LiqXlmrhWBvnTGmxmpx0uhif31UbH5U8LJ5u0XZTwJZUPG7aboruSasJrJJzyP
m7pvaYZsCr/S9Kv7eohsuyWG3DJB9VH3SNx7f3SdWSxDQNfBa+3Ls7HNkejdrCxUc5TfHtefjpUp
9fyw2i3eceU1qPfTzcI21a/j1fiHR/hhNG8NngKwgg/UJI3G1vVDySgDEn+LRcwsA0OSb25m3q+F
oN/5opEYUEHsXNNtHnml7Y7P7Plq2DVmKn2MyHiqG/A+pa3Fc0lGtmEw8mEJ6stIGcgCwhGsa7Pv
THMxZ3MBdbCrQJGP9gy1051IUUK6CfIuNwMq0pMCbwkL3ATlBM+oG1QDPCmvDwuple6WIS9wtf1O
I6275A9fHIwuivt0SfQrm7iZ/8iVC1tLEePvtD+fiunx8a7/TUC//BBvZYgyy7Bew2vGvZQU6EhB
PbLg7dfrCxzl+vCEDC7L9ZqX4chHELHZ1orhOIloQeYTvbSdRe3NZ1jlrjt81yqetCBJMmjlzmMp
XHgzYxxOCOUiOOzSsv314LMeH7wuiR0RDWlrjaoWD3FIfnFF/AuFx92+FtCfCJrBNoND36mz4Pop
BeDTcYRE3MAAkNjrs5ep1v3RddXJFMISiJgGZwXcRmfn/UM35eSPhJzkR+qQMUW9+KHPx3eAY4kB
NfWCr+J05jpqEldwRQgckD7SK3F27YamsDVHhzSWBdQp/FWsZNZHbMOZxXQqYpyt7nUn8uRA0qKb
t6tUsIq3wwPIIvRD3YAnQ6ipuFVvkPsMZvBDObSVAwWDphoHCOcVziARiPIOVc5kalNhKLl4Wvaf
bsm0gRjdWkPJrVzANecgIMOakdgf0UdvPCGGdB9J+o8LGqzJELx1abvt1Pn3m8i0Cv87jkDmbboy
qwcwmMcGQaFkkvGT7JDV0boFaVnWVBNJEETKZF/9MhPyF31qrHRlmpJgphqUhMpd4u+akBefQ61Q
GL+/wYNVYwsrs9t8BMqyDA9xpgLlYBshAk6z6x7n8+IC3kNKok4vAgdo8oCbWzyVtSP0rlvSIT80
dLkjzOmWAPCjAc+p7SKznuikXVGxBMviwk/lxHy/yy2N1aM4aBBM0X6koawKHggfy1XA0tz2yVCw
93W52EOzLgCLFNKi7Ui6t0/vHMvGTrQ/ouDI2bRDPH7nEplBQ7jU3evoA1K831oP6gWJ0lohKN9L
qYaXTIUUpoTuf0cOcCcmIoJEVPcGq1zDFDWbhHAtUVKM/8RfUUKtArO9Qko/wgkElqqxvw+HmEUK
n7Oixef/YrbY+hpddO2+15Wx3a2hc4fcKljoxJSr32rIiL3bBrC/w81RXUAAhoC4VG30g/xD3H66
s7DEPHQDixpwbqAYe5tqA1AZPH8Ravs9V0MRUR/29fqQsXxto8TAdqG/S+T2JI09v3TrwZba2lwH
sMnD6VZVhZZEsxIKJcKRxsdWgGMDrl+4dr4uU8+bPv+Xy12VDVCsgv1tKuRccKKwCLIMpLdaTuUU
Yp3bdP5AUo6JPCLEbh3WolF8OKpWAsdR7O3La20TVZhH0/AYsgWOor/yVT78qACfri8aMI4UsIkQ
8F0iBVn5XhiTwIEnCCjjsdLAj/FfdzQhkhArtXkuO8T/vxPGFYtB7uXUADrQ5PvkXmpJbzUoMu2O
uzByPj/cU7lSgU2sRMxrVQwIa3jc1YqSHURQ50eoplkCfzCc+nzLFN4gFAdKV9EmVy9qef6AIyNk
NnP1XLBo2b3U4DzE/gvwi6uoIecGlgR1PrvKT0hv8QdHwuZhPCDj/ivQSNZTld2B2qZ48k/oQVNV
TH2I+6IIS9nd7othTlDvCnE6iMIO67DfCMEPp7d4Kq1u9fZLNz8TL0vaSUjhmym7wkIORXlCea86
eY9S6AYUqgp/oS/UzxyHrFDqnEF9KDW4jKMYCrn8tnJ5yp9lVIBRWJTKDw1csMqLmYePxXT/cJRM
JFV221VEXjL+Q0W4/fTsoaf846xg3abVSUF38/jBaQpTVTOlZCmLQvXL8bBlL/JnzzWQqO6jXqtq
K1kYWVl7cuo3u740jeLmiK9dscHVk62AR4YEGDvwVCwlZalrxAYAOl3w+HM4oRv8CfYrNAWmIzcb
5xKnhDoS7oyxFF8s+bdY1jAWOiGVMFCd0VsPSMYVUrcZj//xVzxSzdVjVxasxo6XCi0dcP8scXAc
NH6gpO7dETPt/fUlutlvJSntypAlZqi/VKgO8MWpTvETFHrRxBg7hZKO8O63qTvYCSifQbKdns4e
6ELc10kZbS5l2l4VcKMMKsuoPvFjBQ2rV9OGNlm95oW6DGuU+Q0F5ihC/wwQ0foTnfiByTPLWAEz
YxAUD4dF5YcE2bw1qHzQi3oQu6Dj+92fA33bwpNOYfM0DV735orfWhFLG09lYFBJAXJz3myWhiUr
2Bc6/E4SIOtqCpLheuIWMnP/vGFRakrw0TiAg4Mb14lEV+wIKyRMfi/nBM7Xnckh7C04TjBtZeAv
Bsow7mo7fv82hJwdGbeN25+03VhaOts7qITfa8t1gYQmsSvBje13v8+K82EZC+JEuA+q5GBVQm0O
hJchLn2A2RwGZfqmCETbQuN6GyTVvOciZQGYzo5mrnj3Le7QocOWceXTOPWnrtYwc6dz+liSzafX
5q0JwmTxe0QXwra5PUA2mg6ArYMYye5C5ElwJiKRERxT1KQjZBrkOI6TNYlU4bZGfZf1lhSRxY1O
XHS+q6ei7FywDrMo5CIoZfoaTuWfUBzAY5lxmFpV3/fv0RFFaYtfUrPQonQ23fDVRnkb9uZP0pMp
LztJv8QRERKU+872GPML50EP3PwdkfnMiOOtVFldAuExB/N5v9QaKNk3np4yeAjKVkpQIFQshAu2
yCnIRMXzIc5XPsPm/gw3dHazJS5EnROnNqRKg/W9xoxq6SVGSKUXpMWBwqYCWJpano6URPzilS52
tX83tJCZ3VNlPtgicwE0cPuLOfuO02fphbn0tBGZQu+cEcJm0OjHYJkOdCmDqrKomtxne42ttRVf
s4Ogih58X3KPN8zAjn0L+r4knwRonoMXY+HWfBtJtsdAhFLFVeXO04+nhx9tr0qTCkSAcVUFf0PA
x+DelbrEyUCcToo2cTp2eC6SNgb8NmaQbvSWzPTE6L2hOnYfDzYRx3W9xyDy6jM5IKZOJRguQLiE
B200vnBq76D2hQYRP+yT/s9x8B4/c/0tBOVBRNZFpfxza3LbNUllhvkf+c+RcZixaicYXbRGzTb6
hIynyXaS2ASPisIF9huVXNTp2RtkfCWRcy5GM9aGngTjqkEVU8vB2SqfuqTsUw4ZndXDTmMGSq+g
f/6tEdbHFpKFfvU+Umz3N7/FD1FdJmXdsCx8C65xFSA+AEmoprmOoC4wMSC76HEjp1mVDZyaGNop
U4lPFS/WdMR9ksjDgk1vov+oEj2WoT8gumCnx2NBwc9QcuIvokT6kJjfFawsxXajM8sZ8TEh27vB
d5Cb5fM6MlC7plbjpotKmeVBosAeNEVMn7vwiC6AJD5P4rEnVVIRY9bIjGsyPrgSD8FJvbSPwGHg
oFdgL0IPhnPSDr3J9mD3lmYlm/FbT2/ghisUtHKGV15Y0GMvqUFB+WUBUMWQ3X+6/q3UXismc2tp
18v+ZGTSd8nDaI/itF4Jk9MRB0oIxF6MyML6Qzxa/7cDlLKACyOQDe/KoLVgpScCoHneBXyBkRzm
zKdjp7U5Y1BSFFwLqU4kgRwdQZxiVB6TKEq58Mer1X/HA57ZpGkDXE1LJQ5+HPOdS/bK3JwEg16Q
5JKRF1Ekf6SmLdfhAuW28zEYzpo80HRMNve/gO/6CeYAYbaOf4W1OaVf/BCMO5kYfgaX/PPo6Kf/
CBZyzgAfPAgGxyyYgNcko0ZUlj7e41BKZlY3yMaXpYkPDf6XidqZI5SuP/WTfy5rDZbzjNjMRILR
lYqB6ig0KZlL/A+hPSinRGmkDUukmTAlW/fVvaVDvGe90BLai+01GZsiskscKKVwQfq+4d18X95e
q+JJ9dWTDVrlmK3Bq/v20BTZONAqCP20v5d5F4Md4Glr5o0Kt+CL7t9qVQZrMNyRWFC4IiNT+ZpU
2dj5cw0mPAhHrr+YymyYmbjGKnqPGcA7g/A7FAdU587RyyYG++LEqW/UB8aXtmcpD4WRj2cyU/0R
EDUiy3vIG+gw1RC3PBPPcLktBJsZn4uwlEebMN8i2sPIouG88YLJextbTtyGWI1IC4YjggKkk5fT
x/cMmiWDC76cdZI89HLkQ66rcBXmSL7LRCE7BTz8ISb3BZSM9GRfEy3axP/MMBO9c/DLULlDEcs5
UmWhqareVy/OPHDKIb+cCYWRht2nXU/STX9JaKSvPZKj7rOrhv5YcqXP9cTgErzSHE3Fr2my8kkd
jDRB1cnIAmvCNW5aJmkBt0e0hsVZdpwnzdbJdHC0v0l4Z2lfa8N9CmvX5CacQ2PAsdx3uWzczvX6
AC2DoMJZOM8EYJtih3sPN41hJhW1fa4HIGgAHMT40B9moIdGNLlcUcvb6HuSVivhye+J+56FqUsw
N2Nc03bYpqAInMd1R3jUoM/Fw3LSaUcYBFswnDUP2QBpz021RrKRvhAMi/KBK1zwlwj568NM+XVt
sUklg8S7eCVIW/SXEgTLlcKeGjWBjoNtz8bfqD2nLKwCtP+2tnLZGdoMheBTdPwkAnxbAoK7sOzQ
zz9MuzwO0SZDvTCJfJrnAKCC7GvuSMBYogE6cUxf6GBefw6abN4cEUgE/zKTIDe1PaYSv06TxqbO
gzwySiWsSbyF9+NS5QumKHLYH55Jm17TbHu4/vYIiQ0ui9xxMmEsBcGJOdIogMK+SZytRQK6G0Oy
1laZktO/6Sojr0yAlpzE6CjRTOPLEXw9lVoM9ZNhdbZXTPgNdRR84l3DDCeZps7tqwJ4PRztuO/3
Xr5Jaqx3a1pSEdE0TCnyvyvUNU0lerha0lV/sLhEbFk604pY0dAn4tKLrIz6ItCrcBy28agocOY6
aKMCNwbQQXRP4TvpuOk5kaLp2fBOwdspNfLJK2Xbkng4avflYG7v6DZxguqwaFUDwkufwLrNBRDF
fSdc8uZ9p/4m/wc0AmF85NMoT/3h6Y0I0USi5Xzh30GsPGF7lJZirWQo0O7AqNjoEZ1r70r8t/Yl
dMH5B0VzJQoN8wCgNuSMpUWrler3rOLlqY7RJmdyffXrtQsSBGJpj2ucMoBQrpvTvIZLPL++RtrJ
7MHQay+wpzouLHhQDjIvw04YEkeuBO44hBMe0vp3c5K98LNPFWoI5IPfuVE2RpubuSQ+Lmxkvvyq
wXcINXq6nlItmF8H2fiUR6BNee1ZxiSFbbQyvmmFyCSDgS02ILrqn0Jm+LsdA6q4SNyxYhK4n6Bg
W9HZpChbosyHo5Ux9JKAfyGkweUl6zAtjz+y9wF9tAxpJGvW7Uj1XlwitFpUSN/dFWUWeoOtqdSe
lL0MAHFshr+fehS5gyt2i628gy0tUSOSdFcbMc4VNn73ox6laYIJWNKEEu0IjUUNMo/3UDL+WHd8
9A7qoozCBALhhDgJpzLKZjRSu4VJfzuVQVgU8HGJ55jEV4gSzLtKsOgGnOyIgUM7PJ1E9uPbSSP4
iqsaAuo//5/46KdsZ66zkk35Bq2+c+r7radXEigNeiMJxyDd2iAwNIv+rtnePJvu89xllCPfULyt
vpRFOHoFejuk3PN1npjQfG7uD2SsNOp11YEoFGEwCcBYwpnzBQ+7/PgImc50sE2Nj9wr58JmjGl8
G4b2aCtxht6FT33D2InAs/CAPTMxOWFZWiVaT9pZuHLWr99H9ecFikTAQ+/p4iBQihzlbO9iQgWx
d3T42auJHu2bXa0mw3+7TCcJLfhTt6DO51YNHEubaVfOVqeE3LUg/OwraxKiALzzS63Cplm4GYAb
Pc6soBXysBxYoCJ5ApIivQ1aR9sH9ebrwzQhlWN1l7RuKKHhZYU7KC4tqIId2aJyirxriD5nuQQ8
1OVvljKNg0VKDO7Alwhjpz9HLkVM+9xhIB2ZNwOIVl8LxC166vB5yUjlqP1Gm0sgWr94EXaoPstu
LETNirtJ+MAwcixz8Y6XLcqHwm0BzLh0b6DTnvFiRHGk04pG2+5+9+YVbz1k4BJi+XxvKRrtR2Tq
b60f4MmZssm4YVvcn0RfEcOMOPURscqLyTLL1lpd+fmct8+ziEdUCn3Xh3Xu+/0BE0y0zaOomuNl
W7D3j6rzrilobKb01ya+yIGnCH0WM0O1NsL0b2n3u3hbhSEa1dJ+H8jF4Fopcy8NgCA9TgQV6gOx
2NmR3pOhv0NDOOEnSyVNUBH6/FvjqUqvUb2s28e5cZZnQUSCgVeMsFjXO48fOe6Vquy5wV+p40mW
JJJBTe+HSEQYoV57f3eZcKOrVZmsxVD9orx/Dcymx1YpBhFreOiZhD+Jhz4nrPt52sgmtZQ87TIu
id1jCvsel0Qz1bYWHYNF9wwZ1xxE59obNXjf12CpQI4s3JJfRFjZCwogVjhC3+Ivr6WSLhPRM6dz
Mbl5dDNc6I7o3YtbHyPNU08IhC51MOAvE+IDeBlmAPqEqeAPosR9hJPmxQUqPqbjU4EsbMzDphyq
OZ+2gRGijurLTcbuhIq5xEcFKMr/LFdQc4v95XuhaTRa8XDLPFSjg2Gf82vdso2roEZXn2e5G9sH
4iXPmpXfa0jkdCIhfQ/03TFl/U9Z314Ncu4AFTKrvWrmVJIomy82aABCoq88rJZKqij30HTFczsN
tLVKpF4kDiHGBscdxq8A5MPjlr7yqSPqq3YWZO+JzrPECGKtJ2a2sp80KDiaESDgq1NuDS4xmlX1
U4JaEt0ciW5mEMl7ganuwfGrnfBqSYJAi6dAwqmjwqQaWBfrawGBrA3lMd6DYS+ST2T/zPYm4EjO
DLZLZvTEehh/NEuwj0NdUc4GU33WrdPa+p1rJuy7IYUKQ655TUD6gG1UcnudY1EVI07O0li5dy6M
6coUbcQohpJJkoY1KjnfUw9OpNdt+NkzR5OGMOdXPKsJhgC6MO5LuwEotyBwgQ9uCPRveYVmSCUp
MZQieKVNitbIr+Z1bBXx4KCkfn8sC2UlHZ1VZgliPhSTZh1uPz+dd15B/fJyuwP2FBH/ytc2SVWi
ut8quAA4SLbw/r+b1UMsPMwfjJ9hpw0Acc22XUTcmA6NlLTEw7hM2c4fIdkn2U7Cr4eiab3Km0oQ
QSX+/YrxzdUZtCSwaDEwYs1GBlx3jUxqeqMYblZtFoK5HXaECoap73ym2VOrANx4QoAG5unWTQ66
viCYFI8xlI2GC3HMDlm5rjc+r+MQU4JU6TafJEZkWj3E9bQE7Zp+wH94o9fOiMJD1TIPfKy+jN+u
EayME4C2c/vWpEo+vVEjpJ89VugmJu7jqbdtwCTFHKxDZ346FobWJuKdNKAhidVARHKO4Je7r5bE
0kq+xGg3Gnc2E2krHHKIme6wPn14dvkTmcT28/QaN63TxO62YyNGCDlzTai2b5ADQYMwIucbtv4l
85wU9vYMKDFduQQq7w0CQupy5kZ9gYlCycJjI/+WrFZtSHmYL4V76I2ufgGK+2pvy6ZYLiUmyduh
nfKWp+yIWvo2/E5ecnwItIWvtqt0CZMuzf6/RMzp6cr2YTrVqMu38vRJ00HPQcs/H3IT7iYeyM3x
FFJCOhqIHROHoZbdlZBnx/aXQSEmzF/NaS1//wNwLZolHMclCgA/cGwUYdhiF6GE7cSRff5obgkg
ebyRVNTJEG8drhXYGOKLZ9Tl16PzHT9CpkVpF7q2ITe2kQz3IVliyJzhg19yQceST1m0Ig6Z3w4E
5DORuGWZsPI5nLdUeDQ8EvWKmZBGmgJ4unwBHwJJe3M2JuB3sDN3TmaVALsI9cocp1OfbcmLwWRN
M9eQaQG5Od4vU9lngtn/gp3Q6lf/3oLo4mzbeyq0CHQzAb6B3WvAWc4N/KImCrI2IOOo7kurCNps
SYLXm37GNLmiTLYVFHGqBxKWVoiiz9zkFTOI8AJNQ4hlwGQWU8dDeKPoS15cxfS+Dl/006YkGR50
5NKZCH5jpSmwt0gPEHKxe80eCYp4v/app/+NtJFy2VlwlZJ5IX6WSAMO4czBlM+h4Zyah5v1IGz8
i/t/9ukEOJqC9p82WTpJmyh9QExOnEguMf7VuSY7JB0y4blSTJwxXXzUu46v4hZMUSCGmrhYYfuK
nIMsx09qYCc2QdzvgeiIeqkavQakL6UPz7TZacLc/Xf8HBN/5l2yHyg+m26jwqf8iK/J5KG0W5Fx
1Hqu5sPuJsI/S9YZbzHqnl3NDlhU/G9FYmlziuOt5V8aRnN2GtZzMooQLWthQF9a1Lyg7ge2Pjas
CaTCWiTh1AJQTaIBi4KvmDBQONDQUKhevTWnSAn2zhPg0EtJG+xBXfcLB3cdbxliFmhd7F8cz1aM
0ozAbFvWk6ZM0cSlHkwzQppb+zIWKo83DhdD6KSEArX3ZOo+M5rr4UzTTO2ml6BelM6JbmjHVewb
GywGGtBK1yxjTBnRwy5LZfrfEIKjKOPXNE+hu8dj1bF8OI1gIAyTPIcn81x/Aa57GX3rvMJxeT0v
K7dpq1uq5gnWPzytLqRqYIoRnm0xelzxjw48FuawWFFGwj/85t9v2i1doa9Xwdv+W4F8nJln6NaW
ipYhlVAHaR43YmSxd7qpBqL8FuLD78UWxpirTqKHk8m+DUB/tf7EgLNnQwakzwWR78thcgRRWrM5
fVWg5Bw6iu8POT5j3rL2ff5EGLCBRFMSvSKZk9pluMF8F0cjkIXpHcSs/KShW4hdN1ORBT00IT2m
LWwXuDcNN1zuEGshbFnh4hC87nVi1rXXfVGg5Zkfq66YAT7Bgb0zDt0HgUNC4fODq0yYfi/raksM
ny3vigjx9ac3Xt6PPZX0b1PZFo1EdpHzBUc+ZuwzENg7YjcsZHaIYYqDIKBgJjQRKslNjEiWL8Rk
Uzb6i3zaYGdox1mxvc39Hw1F1ya4hp3F9yG2bUck0ehra9NUAmqhourdgO6Lvy65cT85WezXAvjn
0oSohmwUNyPriL7/OwXJjTiahj9yrpJhCoz7hPJfGkWXZGVbIvl97v+EZbqVaR6VTnQXJfql2VqB
EiubsYegKaOWkfyBLS73r+qqkXYic3XrX9i0l7AIKvXf0RgEmK+ojQf8Cqm37jDqAC7V2nytxk76
CO0sz60zEHBziZV7Ih6MpA2YCP7jVqRcqn8uJdf99WadfqoS6P6nJOIJ9ZsBbtm1pLFpaj/YfTwk
qt9KPKxttN9c8fIvOp1opNeRe5lkd4dWWTXjdzF+vPUt0dzsNPtZw3c7eITH22WE1vyziJVrpeyC
opNqyQTVaTj1PQ3PGGExDRX/tFSG/OITmlKinp509GJjr2mrnR9atTGLabcHQOkqJQMKPNZaZM2o
rpKmBJ3P+Ke5rJKfH/ebVob8KqNFExdB6N/c2BpS0BH3LKlBMiVnIouW2EfyOMCL9u/Cf3BTNd4W
x4G/zjZY/eIvcXK5TLPW3LN79tUogFX3e/MWgzsQB5PkB6pH0LmwUPmUytnb4vCceCsDji/Lcsl1
D8hIpZ0s/ZHwy7ZBsupz7ulRZx7pPW9QDPzimF99s6eDZ4+SFqDuBG8Lm4IDZcr8mW/lV0HUcHif
YosUBKWneN5NdoxxpeiTbWUXbF9W9O0Tdswh83lOLASyR/Ux2rdiPYXLC14uVHVVlnFaz512BqoF
E/HgepAwPzGrbmJj81kCAdybpGgOmeBiZLVFjfWTWT8su/ynYMIkxhjgn+a6iP2tW0IUM05Hu5u4
IGo/KBojmZN9YWVM9CUirq6sPaLF9JRZlAdr7OhLLRvWa05zM0vkgULIEoCVAq17NT7plaBUJJEP
Qcqg6mJDRZLKNjFmcDmgDP2k+g00cD5rUbQLgJJHBpxGuMrtmM7aJEccIXKfMeO5wioZclrQwBOw
GsCes8WpGa9SpWipMeDD8pAgMQLEhc93Cs9FHT2aD9s+HArb+LsSxh26wdURZBi6Yq21XuhxnjnA
+5+drYbdyu9busgPtbTQcApqmvsNJYVcmuroQMQFKuWvEVOUP4CAYmIT5vzoK9pTD7uq2axqoxTe
SahYyV7Y+SkvbuVfhCSyM8+vmN1niPGpncI5QooF3lxqovmhUqhsdpvRZNJFCDOC8TtV+5Q3Y1lV
gDkEOXOJWWeO7VsDm/NHaaWOqOgsv4vIL5F3CXuxgBRvSFHZWx6ZDyQ2IdxN71+AP/4NnY8sVVHk
8xosYvRCNjQs9UkbcTGXE0MzHwfmbCO62+OQca1v1gYCRIPIrlHPG1jdJ56fBYrBtQKWwxf+ro0X
6YXDxxZonq23MEPkz+L2JPAa0KSZeJOMJHAttP4GUnPCD/ngwStsf3idyJk4s+XkSEGS3BPHyisH
/tfTFDbvKR7HRBif1/1Led6fLVRuPHpWAfGGfWDOqB20qLToG7mjYzoSy7RqYCXkRa0xwpI4icrI
SwO4lZvr24XhlW9e6CLZWQHV98n8egom1EA1NJc0SlZj4bZP28ipiM9+3vveU8kRe2/dfyfvxyt4
D7dmsc00x4O16sZ6gKJHD1tAHQHxOgz0Frc1e7kinTUqJKQAcbYZMgJgc/tFoJFaLT1ULeXZRxRO
wtXPlX0GLeazdz4Gn/+PYFv5y7dBxroj6HXFB2/+21lmzr2fmKiYJ86IfCRW+cKEbVGzSyW2gMbi
7BCr/OzverI17Uy5rtE2fadnqOAesNIl3caT64MzMfOFjEZVr+ZGAi+LpD/QivMibEakahd0CWRW
48PasibyNHPcWYcVyCKWdcj9jSQLlVPc9IVFYndHbOINcNsrcXQkNYPB1axmFMo/TQ9VdDsspCCx
KXUqKPcFd5eHm2TAYmLtS/xueAEyt/sQE76U0hTgpZt7Z+JOfZAKFBMk02+yH68QDzy4BrOvHA8+
E4x7Rqz6b7rC1Tv+jpsWskmbCdJYrMZqhmGexgX0868u2Pv/bXlT6+SiJZNrqDIutjN8wS9FNhtr
ww1FkV7eKIXroEYfot/lPr4WfsUMduXt4rp3xrvWgK56bUHlke1ZMa+PBNbbvMS6NpHx9NFTCX7T
eStZG2AwtC+7S+0YiOwdENfB31/eBWvw3GXDkmcsUQuwARmd8TrNNpHBHMKDdFj1ChwwvjI0D0l1
GRafhXWlnONpUVm87cqpLRubC9fFgu45xhnpaudWGgyiQWu/MGov4p+sFuyozrpbN8bElP1l2f64
nJ2zEhMMT9GShazTQIUY/bO2m631NMeSdGb77gftlpdRXmoF8Z392uvcGvxjgA2pSYxx1NF/2vpr
x1VHVJuD2EpEI96pm4Ast99AZq/Gxd3tGIOHmtjKSdaUUY22Tg9i/o4M91bh7QGeLDQeEKuEJnie
2I3ZFzjdtG2fLuFvZ2DwZZf38DDwWdU2ysMZigHTjDlKy9WsIB2ACZ3KUnOLPtZ4qVpEb2oVTI8v
0xGW4FKRi2fzqZCdMjWnfHEpFRYaThoLJteO0GcZ1XhpEHKcAe796BRTGb6UoCZwpk7546zBAQCf
ceR4m5/wIsnbvJ4MscNdCebu4uv/01m3nWXcplGXz3RZqTU/iWOMGvH3cwaSLaGYUElKhjgdSOAQ
8XQXeX0ZGJPodOKlN0AAh9PI0HDIRD5uZsGVMSD/jImZGg5FP+NfT3XhDCJ7XL/YC1YAv4UkumLh
eJ0mGU+zHSUL4ble+P4B0J1M/ApO8/NOdVgXwHcBNbxJ1rcdMJ3nPYhzmt9mr3b1r5A6wk/ByJhH
B+BBqey4Swsahrc0iJmISeIZpu2antV32RLekjjCwUgW4N6YsIAR4fA6j1L/gdst27WjMZLWjLgU
+aL5Cml5mTHaI3lCV4AnLjvtVW/8yPJ81iM59aawSr9gKNNfsQwjBi1c72w+VgPsMEzva9XZH0q5
jnTZFM5EFRXoPVREhvPTGV4/a3MBkmusA5bhj1uGbq7uCQJVu3N7ZU6ky4iAX7w7YRGfL0pMboty
evRtFjoZp/QzdYw7AfZPlWWVUSelFgV7cHpo6y5CcehxnD+SQ5PjPgg8ID+MY+FzdKJxqsFlneq5
SrHuoIOdYXMui0UjgBG54nnN69Sk0BluOp7FjfG/ZdsNYHMxRX14k2lU6OO5g0PGMgYcjWfLJKih
l8FqBsie+8StuozzwFIkthBvUNpyrFEsjnkQj7rUK0U2QU67kY+KdeF0/uouOaDC5HwbLciAqJWe
lUo0M01vqC03LU97ILz80TSIkiGxubcveDDBQDTRMNz+d21UacSIohfiwdFkx1J1U83AL+eekimu
ls5TowYWXqu/41toQ8jh9xDpFLG9ikQ5B2wQ35IxTdYsZLPZD1C+oB4cL+oB2iq+zEilu9GUn0zn
/AgiUTK6Ox2whhdO+vuXepCzeaQl7pkOkp85nGSFmyBRLUoinS6j52xtt0HwbUkhdJe7i92cbrMK
/PnPppLPh/a6G1qsrJYncT2Z4SUFzbxiwake6rB3XGArMBZm8QCz7uVJGmjq6olREng5pfpjGZVe
3yhc+KxykD8vfAezA0uuNuANly6yvEcMgd6LPegPdpljeOdXUmItGi9c+12TPwscW3QqzHS6kVfC
p9i8dnHThDtmXhTw3tz5iTPE6Ba75ccrO2tyDzqn5IGNtgYy57QLTfAFwIm3nSo0wk1zqWmlgZR5
Y7lOKiG0YSb5dZ7SvNui8oR1X1NCqOGP5gIkhAZGDosffbcWtewj7CEXdRG6jXYQIFFP4I49gCrA
v9tDi85fwnPcMGyjJMMa6+OlP/XfXxDpx5FioT3A7tvk8ogwljrbc2c+/NQukqzlli+GmjDsJ325
38nay6nNoxDmi5q/0iqG5+SFzZ70/szpzPNCvLgRwmV0nNNNY5EzWXuIywaGgR2UHcsAKPdDTNLE
aCtKcqp7XVmtTKldbf/gcMVlk0ccVeSYEquBabRSw1lT2YL5+20+YdyCk6YVNmz3/MiEvPbVa2rl
y1QKfD40MUfvyUC3qailE0uOoPReJLzVH29a3AbYq1jpfD0swe3YzN/i0hSjv6bdAxjT2UVwqMUg
jFt9SQJsdyZt/4ygLCcMV08XmcJeHM+RRB1LSkxIDWM815vKjQ9N2LXfqvTyShwre3j2teBf5RRb
FDw1uuho+9kzh/M7MtdZM1SmC32FhwobKLgjPO48GeY/Cc2y0qMMboontwMr1ZnufFHV95EeityE
oZjg8lLTSz6xwghvZgPtuDtupfTEc7ofJYKwqWOs68Qt0OqsCwFMRcDCxJChApifwM4VoBgRCz9N
wfN4fI4fOOCqTnDeOxnSiKj2fLMSxcbDr7UJ1JGkcC6QMQKdDw4U6CZbE3dUklnqdUkT/2uRJQ0s
X9hTKttl4SH17NjpYzuxP418Xqk5bScv9Y5qC8icL/LLdgO02IRa6X2uvjsx3YznV0zgkdVrL+2m
3pHJMkSSHQ6tqunge+O/bbkX688tO5CfmMHSCkZ4FZswPqWXen2egvz9fPXH0/lXUam2kbkNgyiT
m+xmi3SbfYmXdhkujiNXHgR5UaUk4Nh7vXRwqUF3Kw7E9c2SvTD+1IhzqQ1aEXlISouo5/VV1iKC
QZvDjtzDDVDREX8TEvQwX8l0CnSxyfvc3GJvT30iETwnar2NReZtLQWQrYoL+875Prt2IyhJYATp
SMKW/gdl/CbjUFNRMWBeEmLpfpLag19Scv00ah0EGO2iMoSdCXoMZfzNZOyrNLXSh7YuYGRAIgLc
8Mzp4ArrwKzJSPSP6QpxF/QIz9eE9hqYn6uxEBzf+b2EU4PF5Xeo/d0O+a/7UQhYaiQOWEYMVdMA
2H5q9+T6rhVtf4ZNSh4J/KwAH0YXfVT1EMmtrvcrBVKSf1Ig6U7ZDjm6/1+dYaazsfEt7Ve0mNkh
x64VzRsKnJETpMuP7W6WSMsEaU0YxHl/de5ozBYC+Jv4mp6TIGwS07sOeagZvaYztV8gFoZFRdvq
mw7uPW+w6AjkwGKKHKgfg2J68BNhih3cmMsl4EjFq8Q16NXh7wnK+jraudiJAEHDey+FxweoJM8W
ThJOE7cModJTEdR+rA/6GtcXmS/JO3VnGczgCJW7oiRkSKyGHhr9gqOs06AkyJ7r4yPU7qi6sIN/
qmA/72uZ+cWLffWzstqz6FGTCl6W80gF02bS0FejQ8UGO2+Jerv+HgAm+CVZDs0Swe55OXrn8q4q
ymSxHlHqONd+6Ahrflk3KNPdw3JOhu+9PK4ZX3RpauQ8elrkweguuedY8aW9HIqOcXIfbIV833hw
nlrXiyC+wKCCctF2tEak2t5IHiVNtRDlv+T1bGQq7Piz/P3ZW4012vEMpYTK+sBe8kCEQ+ZvzJPW
E36MEb9itoJwWV9VJg4x1ha+i/UNws+uQ7ufUUgmCHnXgLLPfwjH9q63OKmXDJbfcd3yI4RPxiH3
YLAbRkIguNk5S5rD8S+Vu85YL9urDb38MBsoGWWCkaVu97UsLkbjL9aJwDAOIybCYlKSV7uMjt/a
2b11dC74nEJNGg2gUao3lkS+s8jzQ0AozMnovO/XjdLXMK3+m1SkqkCDcgi8LDN3wP88YeinDVhA
Un2udRMCiNegM4wzVE39WIp4dlv2XamhSApZFOmGY89M3/nvO6TKzhmbCWaitNxFvvIbHUtpVsmF
kDPj/BAGyqlR/asv54WjD1QdZRwq1P+Huz3PFbcPSWqvGYH8l4gE9ud0yK3YZvjXrX+CP+R7Dy7G
QtA6tq93v9MOzBqG6Aa/I2ccmMyWKT0moXoQxYrj8g/hxo0+27jBb1AxbgwaUxUU8Zp2sDB0Eh4f
i62tLp3sCPi49NowVnCl197mJ+YBQxBN60s4L78dxa6joClvfl7zAmnW2p1mVcOPSyS2y5A/7GOB
1+atzrrvyccHVNaTYqLMHRWpdxOwpQpjcMXp9XpUL+K3/lgyHnpdmK03l6oipBPaj4mz+2dmOur+
67dWI5NkbMrd/fgHNy+1tbmRUICfz+uKMmW+n7QHXzal+CcMvLYkZ4AxNrGN5aHEwl2jmTp8OXzI
4ucFmOeiEFLDWiNtMlSVx+XuQYwyTxKtzcCHcH3StTTJF6FEo93njxNW6J+awESx9EoH5UMTVDzd
xgogVwotn2sXrTvvw69TODtMlzEMRKZP73BeEHjAIf2yJ+dByYGo4lOytHRU3HIl9QHTS+i4Mk+S
Iv0eNPc1PMrbo8Pq1z5qc9B0uGE3a/0kWLkjoYM4FMjqvztcLxUGU5ahiIYliWlzNzSbuJvq96K2
zbB4TasIh3dk7FcJqUMbjKxs7DX4eA6XhCQEvGjZCLJKP20m6vvjP3J/LwTsKNElORlPYqbNHBMD
TpOpBPlYqhprc5UKq9um/R6pu4blLj1CQ9KAuumbL5w5ALiIXjUAUwHwqklLyFyVq3E/WCcifhQy
KHU0qw4xquWtfhDGCsJzxvTQbPdgWxO/2jbP16lenk0cq0g2j2jOY0Z3bbADSgma/uTaWYSrhRUc
uGLuRAkazHAB5aCnTjKg9EGkRSwikMWIC9QO8GTA7LUsXoEW5Do8ayDM3Eid+8grYKQxZs86Je77
9aMm7HEHFj+zVQ8c+oN+rMum79jzuAYhTENR9kfj+ggiUCVFbMKa4X5q7LB7G6pdJrmGxSI+5KZG
sCiDolYofGm6JZUqGpoijMR8q+QvcWoiW34TyTcG/iiN+9A/vmSbshuqy3pvRmVL/6hx/hn20/F5
hwtq9sGqpvaa9CtyjAb88ispSEi1F8ghU8UxCY7NBfhgvFMtoEx0XogFhGx/2rY8j93VjQXiLGvn
h6sux6Kt9i/+HmqKVs865zhYuNEej9s5Lp8Fa3chsql3/84i5hvu+1eco4dJShZmt9C7wzLSTS4q
VX1wXa2UBBcQM/2whR2WahrSnO//Y6di2Pe54qf1IjDKKf1IvwE+f9SQVZ5sQyWkmowDcIIU5sS/
2HxkqCu2PmAZrCS8hVQuGlUVu83Cp6OR/qQjdX1DT3puE5CBGHKIKbeGqQnefbKCeSJVd3GmHoNe
D1HrJYxD4QRaO8bSzLf8587V+QcKfWYdmuoFUPDyUhVYSNTD4Kg9bD5LB0Tb3aq3DjFZy4lFwLb/
CDEj43OtFvK2zw+dpFI+IYfap2uqMSWpcKFFCfUPbBq43Zc9Y9Jc31/UkRgPFSLVSMk+6mibSjra
182mdhQhgFipWHO7ZR9qVwHfSLEdM50cjfXb/LPmxnvLj6MLc1dHp+Xi920KxZJruzZI9cOrPHLW
Lfk40JAngQcnLoqZpHLDm1d4cq5HjZbKZDt5IYQrhriTsnDvz1LDYRlsiHfzhd093Wq0T/Il9L+k
zm2NFXcxuhVygqrkMh0w065BlQ6BEQ1oSO8dQAyuvx+JNLUCZQe0ZR1W2jATeGcj1mNmRWxEWRHB
JR33O9EPdDai1cUo7B0FiBN7YFfc08+qjJV5iSV0Fl2iLgVSwleWJmCgxtpnWoDkw4Xq++62ccAd
OHgRCRRrTc3nl0+/Gsw5Q2EwQDbra8xAQGb5aL59F39TWCC4Boo5IiZ3cw/wBue5FfJAaVmYHojr
i+dBm85UmnYKla6EmsDcCmkocI9Z0+XCtNj5hQmcM/N32WXb3glGDfNb6fnzyqH78DfBheX6ywu1
zwa09QYv9idiKzEdHxTMrkCdPRsYmaWk7N9ZBusez3WAjf1YCy1OrPB4a1WuDHM3D+6bIV53ltn5
PzpdygL9/lorse7/KBZLeRL+ZyalvlTgL8mX1S3zlch6sy3iNRkj1q/kQQaQbmQ3u6/amxmywEtv
FgpvMyFs/EU1Gca5qG62TO+bgu1ew6PLOysyf3aFvgJmeHSZExGmVjz3no35PXtVzJtMZ2CnWdye
iVMmSk5m8xY8WMQu6JKo4+UY7oyhQDC205TYRiqxuV8Qka6XNAT/2yWXTro0hr1Em3bV2InNJoC3
yWw/wf+XJi3uy4q3nhq+1uBtpYMRs7Zl+6F1f11bNdQxgXghjkp3cfP3YAS3zDk6NikqUaTC6px2
lEQ2RhsqO6/0Bd5DCQDg7DRyYB7xUELPwcb+niG6BE0GUtr3QG+tzDxF24EojIReMFrZnCMvQjg4
pqFYvT5dqp8SDJ5aMl2tTnR2DHJpKQVMg75q/nEAlH2YN9rE6eUjdqTsr8pHGuToQMrIKcWMmPSQ
jHPQmRwwHVdotkyTTzaQ0pbtQEnk/jHg2DeHWS53LZSyTa5eB3yUa8Jxw5R3GEJamXLeiaCNaSvz
JMx8BqCgu24INgY5BqI+EpggUP31/xHyJ5CvvKiIH2JSZTYUJttqsGESSsQ4GhRJGrXfniQ/JEJE
/uyzuyrOzDIFHw5DSdBgt8vHXs9tFRN+pfxiL5QcdYLwWIyMODt52bbevypC33rcpbIm867U/26s
DNpgAFchxc8c8KC7cu8NKfH4JyCjAbv1YWSEV+NnCYqrJUa62iXnRCPIxJBOCLWkRB8sB5L6ren7
IEmY+YzrOMQ3/RzBcHu4PDsQA706e0tZloUOkoyclG3iugrm8LFC0tj4K70LqpVxyyPo72fRXymi
NBclCwHnfBttu9hWSH+UXpuekqXyMFbhoLu1qZWM59lm3cWWYkyw3w2x359t6X5onlEb62xRHJPN
d6xbNIDTnXPb92+YT0/YdwuONoihoX6Tr1YVSRVoBhjHOkfcKDnsB7N+QQ/Vr9N1TSuj3N254xrT
2y5/QAQlJrZbI7uBJvG0GoretKlsrsZUd5HN353P6fWkOK2v3F5YpV1MsipLRDq4umJ63iCbxKik
eqaV66ZRH3xDeq1VIUPupQJUt+LngCwFmSvtov+9b77CrkZM2iiez5lmuVadg7NLGIwnxsyhj2vD
w8mCd6bdjd0r/tUFWko75AzhWleQ4M7D0VMDQ/jGY+ycH3aoIdD3mz40vfh+G4FODUHhLbxkJOpD
LfRLTR14koz7ywEHA/f8gQogakQYlYa1v/w5pKu3q3U7ddjo4nfo/PZJBNVldlO9XYJaaZXkeA6I
0Znm0agrYMnwPjnKJPXlNsgu3UZQCSryOBA9G0VRQSOcEQZuW8h+cUq3akK0VfFOUeMmS2R31sdW
qZi4s/kbKdDqaHmjoVP533pYaGzIr056cQA/HnhIxm/JNwOpK62tdwVCjZsCtjCgiilA0HwBd8x2
qs1+a6CZFXp4EL32HzqXCeSnHzTvg8toC4e9zodkaVJTJwZNjpuPC2VhItl0vk3/zm755q2DAWpo
Oxd9LE6VyPnZbdrWgtDeY32F+HYMUmTilG1XPXoLrurIZnD79ak9eiK0d9Q8GadfygHdC6SbUlvj
MM4I1Cecegd3Nrh2fHtIXXFBYPY3VSCoTEMyBCHhinkrl6Sgrb7GA0gh09ntbI1v9EoyACUwI+DQ
5w6nnESyL79JbK6e3gw7Gxxl2IepURcJR/v7pmlEQ7RLOS6yj3oialtpscatqhTS8koOjozyJ7Os
8+Mc6Ft5DnBQvsB5URAR1Ts6ilT0d0Bm4hsjTz5cgaT6FeF6znCFHrECs7Y4tMgkg7vUW2EFCH4k
G5OzyBchfs4mShMeJ8cv6YL+Ls+9owwsvGkThXQc7S750kV8K2FSLOZITPUjh6xXUwBHY0gYlVe2
obpnm6AxJ3xLKJ8RPW2mDDBun1Md6yKbb3l8+jp96nnbgX/yDUDlAabD3oziAVWbGIVJcWykHJRz
6o5cVux9iY68d7G8lmLS8oHCGSCVZ9Joq2XhS9SoEh4xVa2beuRhi0VI4lTTCanWQthE01fRmnN4
GqmhBIlvX6R66ScfGaSuRZa0bTUIgaDAGYaj221+ILmDC9s96jvVXVkwt261GqIuaLrESRsltv3M
cQpNEueE9mrVZE+6WCqVpHUYu34NlX4/RmKt2IV7GFQJS9m3cXB6gQKic/w7CupAAfHZqe2y01ye
X96AZmyXEKPj115I58THxjf4RhL6dip7v9dkmzPxiPN80y3yfdE6bxqXw7k3Vd97tj6DWS1LXSnr
vKDO7noMIJOTqAvMVYORRibgNt5XR2tGI2Xl9p3xqwzhVEuSaQ1WHoydAPuZQ2zZuMelYC8BhaAt
8w48Ig8piDXJfJFhtFUJqBoynbhOSzzscX7+Odsq5Q2NMRZj6ZTtT2F12xiKkgk0UsgnxI0es2NS
UadbIJg/RriaQEi0j3FvssiLP6XXLoQb9l+8iQ2REWyqTxoAjRVLxHllbsn+RW4ALvAw63/SFpqz
eNUaV2QwSa/HHUFQWNBGXzPpTrYWB0DOUYHHEdFL5LmUB/jp1c3eGH0j/GyFBgMUW1XbLziI1FcB
Ie/f5WKVboHrEbAAWH/w3rhI+am4TH/X760qJtmBff3BU/89Im52BpRrjsDE8q+pRPyppAO4HTei
TvsuSw50fN8t+GlkuNsOdCNoKxPTB7eLFFjmmYyfzYy29jXrlNypgh99mOOVK1kdgCLPHWg2yCH7
H+y3JRbJFrKCkAdfRf0txH4Ua5xrVDF3SuPxrT0lArgl1/5Gi7tDW46D2caf2/L/DnGcAan9W0yf
QUu+mK4uQU9Hb3kwC/W9LZIHDfwgqOJTiZHLA46Ipbsi7ja8KxZ75OUnHnf6oUQIntJf/oskxF92
g5fRi+lrypIphV7Cjs69mdbV0xNXCFonnNkXMCRNUhxCiKnwLBMU9OALYSdyv+X+8NkRF1xiNOtU
0FhZFL5zzzqiyQB4uuKAZq42kPasDhYJcvP+HCfocwlrDN6zayWKwFq6PsnDw+iAY1LFrTHW4zV6
ZqTa5jzBlTn7BW5dH1pEUWbuENLdkJszigMhZ7/nkRR9yRCTXYG9sZ72vWfn4nSIe/mCbVugj3sS
m8RLVVw452DpZtMgoqijIHsmsUpczsCkLnB3uRfgGQX6xiqrIcQf75vfNyqBv5KKMTYwrj1ko55H
31nN41JaUtKCvXI6iaLxg+5O0vFkMl35oEkmyy6+Kjd5TvA8CVPqR28uHEdMG2PuahGKk/wMVDNF
/SsrAeX6ojkj6/CTI0rAovcUeBUWksdF+TlvKdb0WROKlIBQhdRm5NAn5j8CS9pDU+MDqGN76yFU
tslAvkktvKOLiTBm3KhSljjiXD1REfGUP5gvWUjvceX7E/E58rBrYPLXWnwcbY4Jd8j857GVLgmF
YAc4d6uAEdzjWDPj+yAZUK7kpKWHuUCeqGMLM62WAT/2s3o6vXi5+8PRVombOOjslMq48+OWinOW
lF0h74nlo1EYu6cS9N9Nmj5FZkSg1rGohy110wWQ8bj77DgbG5ILfY/lljOugUPyK8PNWGQGu0KJ
ljVCllXPdWxrCm4EAKogNMMu0RBaJHA4OR9S5HG00ulUX86lF2r0tZFqm/cRiPQrwHZnFP8gVWN4
Za7kGHg9lplykRXhq5/tkXbDhtLeCArSCJv6atzzYQV3yJuEnJ0JL1F5rRaI4/hJlm59Xh/D2qRB
i07n682lFBHt3OYhZS6rQT7DJALG6cjHkq2ubfeJJVKjM9Ijuo7NgVao8QnuR9SJwGbZ5NyIrStR
uKizheAVFT2EOKVjb3F6x4skIdEA5fkDME9r5s1mixVnLbpm9mUcSgrbAjRSwNS8usOJ2K8+cdAw
0q5eCCXEdnP6qpvMK986qgv8HS7aW1Lx5YLNP+izk3DIJ80lkjXboiurt768y0JyAop6Z8ba6Mo6
Fr5fETxmW67QjpBtNcKQUnILYmWng+4FCBcCuYyoPjoG03XALf27O49ztnwXeFscZW8o4/gP46DT
nwC4sL3zehf1qEWy2Tp/+yytSREyY35HDlhgCl/JuFlX3GKh4Y4y5UoDlURDtCX96e5DC2b/Ly6z
lxnGaZ7BW5RwBDmlpx5BH4lpA/gSz5e8BCnit0qF0hu99WbTeCE683rgG/L6TekxRthTnMnkeDPM
rryDeuhwZ5u6pU+tmN330VrncXVzW9TgvdAU0DSlRXU5TzAsI33cWdYbJcV3WzFYPuL+2+pu68lR
hv1kwyaH39iZMka4iFGEOTlJLpVDrYVv1xH1MlYwRrVQE+vdqE4VAae6tS7a9eOVTPpjJrc2e4BJ
VC7YYlzrN8DULpy56Hsq0ycwT26B6Hp98ZoBw/Sipy3FInsZ9DDxx0VeU98PhPv7DhoDppo/ozd8
FMjiXN9szooLbU8Ww2VUrWx7cYsThrYVowf/8YcgMmxrZMP6oLLpyOj5XV8O4Pkv7PAWyh9Wa67s
A0nf0WvxNKCkWVn/xz2oYuvAoEnvZl9eaDGnxxF1eiegLtJK5V9L6plDfFK9l42fDE5g3GdTwOgW
i51nkiEGsRWf4shJUsgND2Ugs8y8enzV/v/gJtIEcbJmzBuDcCkz02JVGWuoqB3ouDvte94KijW0
5H4jGj2XY8YA1lea+2qcKJLW9mc7Usz0rYxP8G58k3HXLRbNo8iAX6PxvK5vx8QzT6kj6j75Tl9T
xr4ZY3Nb+eHDO6Xe+Rya4+s/TMTGbDNFK2Rz3Hn6DgDoGvppUGWOeZey8XpCyvunFyUsjO9sYaDT
ZZU1Xlju/ptfOvAgY/HC4SRIpzPfnoq4K4P6oCD54/BY+DWas9xgXnOsWaQQPwSuST+G6T9ks5CS
XWImNIrJkZEWOmhMVH1FKgcPp/J2bDQ85ULlMTChzl4nLsVwA7hQLe0UFjjUvAsQ2HK64cKZRogj
N/NKIIFkBViApDOZ1ZMLPJE6HgFIry0vptf6sAMA5OGs7qhaoCZkhzJHIF0V+IK96HC4CAo37xot
yOCkqhIQxnBgos+q9+vnednGUmwJxTb3i/FHWuWxf2lfBxBxDNzFkzfHCXIEgvNvapTsy6/q7Qfz
LXeXq7+RCfBUeGKhVfOKvdfIwiE89evwdbGp9l75EPZyD6k2/KTTrRpRNw2QSiP8qB29Pdj0OqQD
6VouWrJA57kW6s102kE5CH9wZ1RtcXl61IQ2hOoDnUnfI9NBpskqkN53lDN9QFt9c9x20dZRt8zG
NjBa3XOR2p/QLHJdZ5dl20jEELSvwbvtoTb1w/8J2ttb/4ECTb281+Z5rDTebgJMAOv3BsafkIZr
2thoOzlbKCw0+9Mmg5X7FI7zX4Ypm4g0sb5o9o6pOKK4AP1i4RCwRZIIs9RCAs4pUlBkX9NifkPl
yoKHpOnUnhJM9L5zqJ24XJ3n+jS/85jbPBJSI5TF8vre2ocTHW55eg7ENDXDqd2PwqEOXnWCrvIO
/JsMJRRF0h9Gu8blilYB+1HGa9yTGCKzzAavEEDUgn9BPrMhAF/QYMU/4emN2zOR9M4tr75qaCx8
rYonONg/MHGpjn42gAXnMfI3ASjlfwu0ho9FEIevG/AQlMJSOQqPTcQVONCWfPoLwbfEqZRChWQk
XEeuqkkGPJbmYrAQwGGL1hF8B6sFw6koTH57lw3dlFpnZ/khqFGUsb/o6YxuMxNuyb3/l6mGxuOB
wHFNrzPVT9AZyAuIjgo3s4/n0sUvuNpbploJI6aihvIqjU6m5zS7MqTd2Llt9WyQM4i+Ze8bV+4A
0HYxQRmsTMa/SL7foEnXiP/HHMrPV2Hb/8+nIVvZ9bATvRQyZZpGRuEGgNWCqkeW/7eaYEsJ+Ytb
lc8vuNWEM+O2zw+4V5NyCfGvg0Kg6EMJ8eUrAc7/TRdGxcogBRXKKmsmw1xyzEMdBbqn5VFCV7Gw
A3cIJvtKboYFEGJVGAbXXklosgn1xJremyXdHUo47Nmb3NE9ezdcemzCNnVATQI3noFh3mfSwMYf
7cLPSQpZdC7rLXaJfzeCGofJRjKzcTRDXTaWmYkK2XE6nFlWfs71BvAUdSVzMgpLGHVQkDt2frZH
/l5xa1F3M+SGCyo75k2UEz1hUqZEbEJ6ZQGvfbBGDIRX4WyL2xf+ujNEzU0YSkLyFFyg9JphhV5x
WDzcLhKE83p9Ki3vMVQN6j6SrFxshmTEjiFJU8/m4SuISQdN+Z32443A//ZPY1aPeNiEclLjD6RV
VfEr2QlRsbMDP2gRmeM5RLCL7Jl2XHbbcBzbcgMWPbbIlHDI/F5rpEjvdpIDhM5uX4DT2Bd7RgxH
TPIg+Vxm//KpkmEm0qszKNIzdVKrqFm+75AqHlYqunbiIjST4Q2qhCvtwuVSl2MZNaDpgJHwyrmQ
0KTdI3RVOOCCi3d5r48b4grupbsjhP1zFWljTKR/D3y97Ue5TtiufoFPsbq07XuemqpdDnG0AT3s
HG0I6Rp1VMeRBUkpPZN4xkirCeWLA1eI/U0YFaMbEZVOipAVrOYUAsYQDVQ9MggDdmJIx7Sy/lz5
jIRjw6gmD6tvKfmoDpLXLwCOunsTRLOjSTqAuAHYz/ewHfnjFAzdd7TeXkpXWZRNgDR/A/7XXB1U
KePkdvXxk1rWkTL2G62AxQ6tSQ1FWKUMK9jkI2n3mimig+Y3vdVnj01sRLnL/W8PHa2IXZOtTJEM
5jDlMDYuqFgw/S8f9n/GdhmoUbdc+viQ6BMyazDCxhsOKI0i1/u6DJGJaI1jlpuJSKDI24oXbboN
GzCv6VChEixrZZd28VHSH4BL2a8zKmMYYFEh5DaWPDntt5qW9O83mYVHdPhrX93MPypW7AAfwUjy
1g9yF23ztwO20p0xkp4JkAh8HXKxB6z0qPriDDk5JkI1XJuPxaKMZCgmdiT3SgB9y/x5KDPxA/Ov
C1Ro24Ovl5maXNZfc7vtgk5ye2o7oaEMUIFDlpe5576yl5bT46LjUCy3C6M7sUQ6wAw8d5gJwrer
dOEIuRzncgDE9cdOlrHYmDsxNyny4DtKzSEQq3RrBu97V/gpCGkMeHGIxgik7Hp+Fgpx0tpDBBRN
LW5c/LWrcTFAJOCeURu2seiDbHPYoeKls3Xi0ie5kbh1A5LPVFDJG2RD2Njt0f+qQ7Qicgq5jsPq
HCu+yW7ZIZeUljwl9qrzy9oR1O/PO00UETOe9IoAhSbK1IouXDLXiTAmXJKJANGWgdfcROaFNozX
B68A18l/fiexj5IhIvh3FEtJjHC04MaJOTXfGNWpNFOKIAIRlEdWPJvVGmUYgFxpBW3Qj28Awf1V
UCD5uRO0LSVDXsxIRYSWaNRRFHxRQ9vW4SaYY1xMFnMmzL8FaEpOFFjfda55KMred3SHvqzNFEUq
DrKA10iJa+VL7lRG7MwV++vk3TeYKutYtHcjDITHhEXCxZwXYtGrb1P9/DpMhJKtQVd0nCUOzc7o
sqaTJLjJy+bGVTxorkJ3aSHBROHrsyTj8z/8uSkcNoecOPpyevb0W7U2u8hFl7+d/+o4WF/A4IkT
vIM+iYTJd11pO10WK3s2WIZKKE0nQcVMrf5n0fkrf3roXSp+PDGeisN0RqwdqQNv2HT7uyDg5+oF
L7/h3urc7QRnEm03LkOY+cH6lLqsmUQ0MOAEhb487flJkitCaAXKtDt9xS6XLDEHOO9cBZJ/JJ7h
0gwzD0qNYhvJ5zIDLKZrUIEtInTJDNA4sFMoou2J4gld+kJncRPBDmRKo98n1Ip90es9imXWT8HA
jX6nQB6Tm+chf42chH9tbqddc2cqEHNkN0QJUlBuf4IPXCPFT3Mih8Gp6BORStj3WwEBE9Z7VyiN
JcgUSSl6w3cDZCCBFvQho3MAj+VyYnfPfq/atKiVaf4GkjNDiEx9bmN9AYdLu+UB+h+rj7rWb5Yv
s8cyhH/oD7ILG00Gy59GxJpsfQuOPAwU6dK8UrQriwLaTWTNUmNQhlv3zHuu+4nEdcmQUbfJ9wra
5C4/v/HWqoX2QFLmjfaa4bkYRU786xWy+CkDHDkqzcFncGpi4TeuTmWR9JGNZav7dI5MT2uTgb18
Rx8idxRh23R7uLI4PMCgIogDWeyepNBpIVZhfD6CC4RIdMLlZcd4MYOeHaa+gm3QUacrADWp1X3L
qbATg697AWNaJUIV/Ck3pxSRVb2MKoHcjwhF/UqIMHs7fPdeB2NjXS5i21sgSiksY9OQf9LmF6hZ
+3+/IVGcoC3+mdG0HUJA+2ye8TtWOebxhRZRlg/X66sgXL1PISd622ZFLc4byxz960cRBlOmEKWc
GC9EmlxDVu6Ox6rNdQQRMQtZGBbt+iqIpNHr88EkwOrRZQddHCjDMe/DSSfvZcmp0mhaFsxHol/l
uqJx2UWpqEwsRtpB/Id6r/+UyXx3DGwH7jix6jQlxMBnzHnT0yp9NnIXwPFeiIcC6ObM13PwO8aj
2+UM8aC6L/L69kDQGkQ+CZvVFflrBgmDZTy6GLLknUbo6kYZ+oyVoNWAf4YuFRFfzuEFaSjutKY2
UvQ7/h+ETfjd4+obIaGbg4htRabHRj4S7FRq6qxbviTWYchxUq/s61R5kLk2Z8GfYr67iqZNX4Ss
lsA+YE6ePiJiXiXkup065V1WfW/YwL2A7/4yxME2h8BBSN+lHgdKjUgK/6ap8B5nhSF6dBSEiJnp
7mH1FgpUhrb9R31JaD6bk1WB0AdQNU8e80RL4UPlGPquPJEgOo0uiI4dZzWagpsfGIlW/61alle2
xPU49Sl66m9w5G+Sm1MG5ORHXMD9ruQZBeP6mHKSiM1Xh5IW5ZFFe0LaWucHNtyL3qEaiyyGL4kL
2H5acB/jVu0BkE5ybtC1h6/X1SZ4uQivTcFUjgOgjbLYe9gr2hPZT40aNxrB3ZxrUrzxKT4R6iU7
0R32LmqCW9bc1shm2jcR3+NCf/KnkNGNiMrwC09utl8e9TLdwdLLZKY2dI0gDr1bDLgpvXtpMiHy
3AuMBaq/0C3rdbwO5m/WUAsbp3IZV1Lr7lX6KJqtK/RaDz36t9ujgl4zDgYKZ51CEBgxPMNRjNX3
IJt/NAF4rCKa9P/I1/ArZAWZQrD1RpC43IabVKH/espdstoE2XCyK02UlSCbR7x6QSnxbcQVnoif
C3kGbmag90uCZ3zuNfkPSPNL657HzGS+XapsE1eWqpuxWdgcl64LJTAqKEaPhWJOO/I27RJjAhDZ
WUZPc0/7yM48fHCqJXVHarMexlh7MP+U1l2Qx1HWEZIflpjw7WmVe2ySC3PBs/LSOvrAlEylSeab
uh95p1GXCBuIj5eJxbLsjraaZgKt7gIjAyiPdTaNMHETU3WhrL3nuRBEhWRS9yXaOdCVn9T62/NF
rD8i983ng4m2mz+5fWOLiEW2TX2ZTZTFRqoafg6OGA607oXigwKSr/8SfSCdIhU8FKM+WmH9cn1R
BXOEAJImK3JGGvpd2MFCTz9MGN21W7+BeU4QSY/bCF1EtlpO7xcAtnV7Pthmk4AJx+4X+G6Al09r
Sn/2+57+TdSX/xUot3GnJOA4uojA2tucIDGTI5Qi0OUHjQ1Mfx9KvpXCidZw60IP4HJYGVDzNflO
C00rvR5qIZER3Lgia7TX87ap3hXNj6bIJj5QF6CJ7j5vPk5/OKv6/J2BYZxmyvK9Q7FvgF1KNBcH
D2lOTMmUNx8hamHSokeTgJk9xxewI3GOc/kC/YoWyqCYlZ7eZiU8Yxmq2q4LgytGn7eXJSB6xTnS
L/l0IQQamFJRSe/bSCtJj3h/53DF+SP28An6kdYERshqujbLMlOYPXG0d/63nH3CxAN3nAarS8Kc
o1hB0BgxtQwrg5oznRU4u6PqWEsBF5DxKTKZXOszS4R0WmnZNAL0Vetj2x33muLIN21wAeD+WePW
Ii24mkjW9wJwrt4wEKAXGtqdkYP/yvxWaYDVKNw4t8EE7zojWcY+/VQzKdaJJ0lfduXeT2SSEywl
LKinptDIWD0HQTk0TlUDyv9huw9ijP9Bv2MP2t2J7ncLHN0luJlF4ktYoxOiNY45OzHg03woVgnv
EJJIzlpbeqQUOmrcw5NBmh0qE9F82dPZ3dglHiWscymov0LGHqD2qtiDjN0bPVBaJq67NiHEe6Od
FeGdItDAsVZqvd0b50pGvl58b12sVEv5oQhWt8s5JhrGIn1LPQ6KoAax/vVnr028RbAiJi4vMXF0
rStxO3F0nuFBFe5wJUzQPOlzB5Wl0ux41IaNKflwA2+jooJfEgigI7Z2V9E+ONAdsxOCku7jRvfU
J12fjwp366LVmiiuZsyp7lf4md9b5r0QHt2lBaKsBu3IFihVQtOxjiwlUmRE6X4LQB5btrsFN/Bm
iDYFVH3WgynNzhhk63O1levWZvV/R/nE2j92JAMYGsyyLaTFYVgw8oya30aSDYwUfARLpS0TTlnv
9MZZ8rGMXK6KJmX2gdT0wFuJpDxsxkXnlFNdEl3CECwhdGx2df8mTCsQP+HrQhk+V1Qedjz0HgCc
oeizCrNM0ns1o6Qa59RpnDGYP+EfnFmw+VWbRKNM1ClRhq3KJfu9o1MCohybm9EQdxwAnYpFOw+z
q5oxCCR4XFJA7aPOaqUVvj6ZOiGX6aPIFDLrGxAVbbPiAFoNpKbdTAdJlFoNTjD55a6esIavJvJo
j+rm4yEKsQgWzqjPfEyxnAO8qFBA1T0xA2PAolFGB43f9PZBukBKMhK0pz8GPHigoBplS8Vy4Vcn
ehl8vMB65D1rIyDIh/vDpS/8PORIveOMmYdZdIqzrTJpA+ZNRjPP5q1AaD//mxrk5BeR1TvgtofS
CcHTDsXOVIflcg1F1w8+PJ7RvjGy9s57zDjc1w4s88L/zpYUwXX80JTgvLosPVU16WKP7R8QNdqK
vL29fGVgV8tlVFX6/a2uF/bxvaUZJ66UmZWVMHHcim/PR13YcmhUqTp5GcBQrzoTkQp0F8Oo8P0j
3gHsF0rKRFysJs52P5/Y+TC6HhmhtVyNlYmEvfza92q8kBQfGH/dbSvQR6j06S+HHYMBCVTz/cjk
C9fjbJsXa106GZy7yDqQWNYNk32oonbpEkSDt9qF3aMb8+tvZaJZdi02UnMtDPh6eqfUl9gH9nIZ
06ABZnsXg92UHqbFQ7gfeml4V5mjvknqVQ/+Mg5BYimm15hiNDHOYkWp7IBVLtMEhse3eJpzw/x2
aFDsfQzarTToVb+QqNJsruFOOeyhVkpzdb9Z388ZfJZs06EfCDM6so5zUOX41PHZLqJvdyUon16J
iMdbwMVDyhqgAw/FeXZJObF609LtPpPDJKkrehnzuEV6rxUTg9/uil+llb4tA7Y962M4Tm2KBFL7
k7yyOdzGWjyNX4Mr4IXF1iBDtFzLA3UWjefokjXaXArcyEpfQM3qSpclRNWkv5a3BbKQBwbAHba+
0TLiQuGZr35bUKeNnB4oj+WURfDUXgu04G6hT/TVlN8jtterT+xAnGlYuNPFdYSMNW4SgMl5jGjg
rEji6rU78pK72R9VBFQZQuILTPzT+9nTINoMa2VWgTVzK+yJrxomvIy0g58eL9q8SNc4ALfUo+4K
IEg6bjsWSFvOqJXk4xDsI1CpSNhaRkGTOczl/Oe6uzZhrxlreYy+LJ0c1eeu0R7kTg+bKQMAyFHo
FcVZjt7u6ekJOCC2KpCSxqCPLTK4Ai+1SVwyuFv5T7AWtSs/oLHPm5oasmlKKsnTmYyoOuobNdsh
ug4wNPFBtn0adsOX9DqzzBuR2yg8EFt1GtGpmWnxr7yWeJBRsFEBIOp0hjiR79AEeR5L0OH6zgOq
IKITcIryqBJpC1R/3YCZGBeRI7sYxehfzegqQReWk4NB5QIPl264KAz98pEWbwtIDNFRo9+ZMW9k
dkfjB+9Cmcxed+tFEt4tA2RX5Tm9jmc/AdCV7J5/Zp5xjjm3IlNjqwXlFEjM6qmOmyFxdsB0/co7
msgnfuygFt81gDXts8+nne/Q1XJ/S+p4FlV8yarOsC+IpYrCz6Od9GJINXaVwERK1nIu/bi7DI/n
OIt4yckZ2xqEosYcRoMx/xMklktKWQ1eCLyvMKo3hDv+r6alc2bEzLcFhH6AR/n4Suk5ERT2LYhU
7/5X2c5DYA9QGbF0tVDSK2vuVkhks9q1XfhrzZX8BPIhdJ80WXhAJy1NgALUvjBTR8QOm8Ym6XjF
aivx6wOyo5R+lKSyiBLbuX+JRWfjab+3M00m6BkzbIITxeAb3uIdIOprZEj56OZz2S+2GHO+Rupt
9JtydrR/mW4xXYLBjA5Lb3KGZJSbuQ6Xh4umB6EMv/+MyjA7JkI4YsSnx1X7MY5qAgyIG4aODOIy
OHvTd0CfW7Gm0odlKh6TCc8V/Rm594NiChuT0Qj+33GYGgiG8nkFO7j7eJSUdOTaO8lUgmE8XhvL
BAxtsWTPqKig1P5cUQprni3hVDV68oMJGcPSeC2HiKO11n6TDgP5sjhmN+P6qRMk9FrZelwHQ4r6
HeFbZrIcY74R24EkneDxqfdzeylYAzJtp2zGn4l1hEksPe8SeJ8E3Q76cTOY5hKmd7L5c7ffRntB
iSv6jql2xfKciOgupbQ/3U355eYD6Y9nMZT1wYjDlimmcyib/uItKTwyl8yrRZFHwUPeGq7/57vv
ykS+mtbwmaL9F8Qwvw3UTTZVovlTULtTw8R2BaMk4UwDXAfEpA0nDetZiko+uISUxfjsjrdxFyXH
+CEBzUIGR/dWmnT/zIY7Xj6FSTeVFwxd9KLgpMxdD892rAzKShcDkgoBcboPwD0c6CANgcxrnigZ
zqzE+WXy7FUHmL6oEY+Rb50TyZSSZRBoIJJk9poTTj7sT2MV43U1nRGhoy9O8r5oZfJ5r1hVdxrY
wW2ZisPy9n6Kkrs7CaltWAurA4jTDxqbEmiFqYPX6xuu8Ap4qwABpg/NSHlxbLZBwyqUnUfICiyu
HXd33jic7JkGQj5l+cNgOdM/q6W70ab8VogmOp6Zd0Y/TAiXJoGdlVau4NYJylGsPm36ioHJCZf9
dvzIOaqIos4z+hJ64FuRroWMJ9qfYJr3eNub+Lwd6REC8Li/SciKltEwgk1VtqsONawzTihayjRj
ol9nk7jTWp2AE9lNqNtbjeW43ic8xUoFETOXGQBjTKdA58rGvFLsf9WmFKOPyhQrd9DS6W9fmwPb
XOlacVe6TPEBkMFZliJRqiN3uashRksJFnObLS3VQC1AELzesSSWeY7p+oT7PbVazc1tMBeXa7Oc
bpnVaStNdWa82Vmz1N/i2ZZ1S/uuLfrzp0knL8OU4DLWwtT95IKiAxPW9qMPvdqzKAHL3XwCLrAb
BVvchTr8OSrsxhOt208+qweUQUZ/FiEKusFeFZBunf3p2YPe081ngy/4OxCEsBRsOjtWm9jXC4vS
WG4QykIipeCvmtF8WXXbqFHP1iOP3iX2twp+XKv/pH3mVkod93+KRMWjES5EAfQXCv9kkrUWdAbn
NT+YmzYM4mr4FsvW8+YpXncuUEbg+LE+aRUhTfqKtJTDbZsgXyLxqNs4rjg9/rLI4ZbkyFz9cQRl
f48IdCcDzpFSeujsfSlCmI0C0p9Dq0Au+GVA3QuDKBvCq2Eq+Un8LPaLsHdw69Bwd4fzk+8U3JOq
E7As14Wyspf7kxPnuFXp9/DkqaA4egL9l1DrvlYCN00S48PJZEDUcar85Hzon3F0Bg02SvFqYvr8
Mkz+fFk4tsg0xem2jhZPkRYgzqGostoV+zULqt7YEMrtX8ytmsbOxFbsJRI0UlYp2pqXU8verUdT
asMBuFOdAAgNMzrHvooI8XiSlqXTzKSwWtNiOevFpDtQnPJNYEXyWRDNnohozw4PZ4nUg41Hp1vq
5fYpGeG5FM/MudSk7EHCK/kkt/2Xwwt3/Y5LzXNbbTT+uzWfT3BEkGAj9VSMyEROeUpkH23EETMn
Gnv2l+bDMfKo6zoFCpFERTssa9YnnxjdueMmBTi1EbEbh8UPpdw8SvId+tfs4ugB8SFixg0rXzuM
LiLG7OJq4c9J4s+ybvhfKYiKylKsoW18mkXhKZLur8DvYeFfIi+V5Vrm3fNqmq5w89gp3eQXUdY4
Jsi1XxBecagt2caP7g07EMO21KAh6euh66L0SlGdChIW0509fvTKyV3Igj65SvDOdUSaJMigfvcV
aZW5rGajRygLv9FWBh5H3cYjL418CKblkxJIov8rulbaG5o3N5foGdBGZLLzZhxLNH44gQhlmbZv
hNFxCmOlbzH2VhIn7whySWnVzRWxP7ht1D7xJ2x2LEms27v5FsfDOHrs4z0CufU1QcRF9ZjFv97+
Jua5qFQbO7f4VpXrKlg6qHwMQKVxdJZAzBLTlOxWaP1bjvzGlvi+cy7aPVRtdj6+5FHh+XHInp2T
wh83mj397RLRnkddgNB+C7+ZjdG3CaI64m36SVXqAHB1jybQD71ziEb7Asx4GLO0NhmKNvy9p2bK
MlEIEVQHCwuaqqOlC2yrVtpQyDlsdvyg37Kmu7F9eIDmmtY3a0gZF+cemUPHKPuDspFlJ5USgPC+
1SZjVnnBqxJFuzd7nbxcKLFgigVucIuN1rXNUgs8zVwHMbLXmAEr+/IvSexeztemF6q6cRX5BQrv
1HytIPSvj/sgqDcCY73QUZ9LzilAE+152gyg1af17tlYoI3syOxGqrbKpZhP/Ua6/SXnMcUdzmWd
jXQTEmED8RSvWXBCJ6e/3l7ODE7mZziVzVwbagPK5kK8+1jSUUATvY6B+s1hG5PRW+Nhi55Y5K1X
85CPiPBxKN9JrHC+1J8q+uXLfZYTf/XQLAsqGokgDXDO9wIR5GIHDcsnpqX8xGPS6V5G6qnM3eQi
SVhJmUwAnR3Kr8YR1EkoF39n+Boy4N31VogRuJEeyknBGWqqunAc0jFCJ+4TeBqgQpqHp9Tvia8I
m6yYOKCcaJkWgBI4PreykoD/fS88X3uRL9ELI6XSn7Q6aC3xRbm+W1DofOFNUsjbDpQz/zOg8G/u
lBlI4JmHZjfgmRiyq2Hwh8Yky6YBF/QezAz9ZcY2LJBVGf5uuqFGmSXiVNQDFDNn/J1kwrrlRyUX
sXm2lax7wv6ytjjqmqJuDIfCVQfsHHbeJo+22Ag5+b9YTDG10NfY35vBg+QEdYLYfE9ZeUueHT1V
6jqfNfTziGkban7e4L3zIQhZ6yJs1fjGwRd2Qepzt/C0ZQWhJckdoOD9/NTjmoblCleGKX+NrjV9
jkLIB+wBYtADXGZco89KrTe8P5wFhUZ1jCszvQw53PW0fFjaxSUzfoWhzlaNOizvYGL8exkfrbPd
3HdMWzijW1KdegROsNMatz7atwif6Ouh1yVxNxbX2vlET6mpSvITf9x7A9OFEIvuOd7c4Z+tcBLc
nCXKCS6EfH+Gs3IM6USBUD+goJGGgWGftY/bSgBIEb0Xj15cVJFN9oNGQqahmdrfqVFTAVt8kHbc
r6ISy1KjoreNK+crW5NgVVjOyZrAxK7FTNl68eowCvF8MEZIB2CX9wKpLWRxCxQWmYGG+iXIZL/6
YhNMeOGQid12ruAa9pzLllcB71/EcAadd7ujpAm/ySfX6qJ2dDtKn3DjcX0xRMLtVb3yMhYIQAu9
zk4V/iTf+1ZLgVcdGT6TD8pjhkN7BMszi47gkkyx1+MMU9BKfk5vrtMzvIU6jUp/RD3rb/vT7LV1
QDzMKpFRvOqcnavb8YOQwT/AgUJC4qYxjoN2/ir1V1wq4hl72xBkQcBlsFPYuATgGEOr+vvK/6Eq
f2dkDsCV2lbv9ALHcuNrUH5b186j79X45QQpwg4Qee8WLARQwlE5aYk+H7OHss0NTxxtz05V79sW
3KKF5jvaH4ZJwdybr+HSRf7lTrWqnKoxP+v/NpVC1skR7LAy+6iR09RTQrVIOJJmbu11tH3Hdu+T
ylVZVHhHQ2N+PmwGi0e8P7RhN3NEKiUIdAqTQnM/81V2Yq5k8u2ZWRRBVWpOxKJ003WD+M1XEILd
HPgSpGYwu6F/Xv440U7HdqQBTgegbcHqtHbe4RUSdZOFB8BfzBK47GdJWm97cgF6tafyjoXJnTFW
qc2sxTfJ/x3lWUOU7w5IwTM0Olp5n5dLcr6Rat43JfQneJ5ddFFoYTmA7v0wtfzPpMeRiaITQZlI
A3BgKjrtf3SbShC64DLqU4uXWLItlRtIQNwFbu468o/gG4mvzgHxbHAcZZQNRb5IPQffBUP3I9QW
6vOQWlis8nEk1/6qDKJ1lFKGirMxQMW1Ur1DhhLMwsDD2RwJ86iPWBWT8RyFT2075fyVz9CUl9CU
M3fn06pSj5PIMAsX4OLk9Zaeex0qV4vKlI+EFzHUnKLHjqFEpjiqVjq4GGg/0EBztBsn3ml6noim
JOb5bLWVXe5AcojDeGqw1YLA83KXHfGJpuw17Sx3nJJ4SkKoMjFstg+YXMg1CNM7Eh7QpEsC6pBM
184kzRvSKWEk6dnuPBkLOHxgsfv0m8Ib50YbZzGPsu3eR8FTSanX+1F9+yRFcd2JcfPs55xfvMwC
hDmd9pM1TlSqCFR69DK6PtHLffKym1t4sBBurrhXbjUUuIX+8Z10TTj4L08W6/fhjWEDFHlQzjXh
l3Rn+YhqpbdZdFNAQRu4ObKuCKZpNs1So8J2SJxT0ZIjEl5eRgy8IZwEDvZvZJR5L73izzWS0uCI
H2r5PppY7Ad5zqJ7LXRYi8KX4aLc888B9CuPfvB4ufWAASNokr4aahYT4ep0IiU8k7Ymqp0wP/7U
1STditF6H9gsGr5RtStkHgE4YbEbZgDtX4Jbl2LxEYt+tnwOLa2tJVgmINHSNAt8EC33Wc4dzYOx
QLmoVZBIlesix62bf7a8vKRcT865TOYHWZll7osNI+1nh+FzvG/pbOxvopqbyDBAMwYlPQIv6EN/
6+KEk/y/CDfTkueLCHqZLZqK72k+8BKsXapZM8P/Ylq4PYC/QYcSORtVOiALQM33e7Ap0W7VLa9I
XB/qyKUal3nlx8CoxfUFVEP0XmqncgTqkVZc5E/ef/ax+sfj0GT5oui/lq+TlIH4qqCQLDtXFcEw
lknowPhuEc8dNCPLo1B2Sl8cg/bm/LVsksvECjN8tOI9nbTqfc2FHL54JKOnWUqPutHlPo9rod+i
Qi1tlu1lYCnGJXutuQHuHx7ObRi82DrMlTVPFgmTBxj/8qleNWipQRacX5HhE4KDrikWvnt1sP/+
VgSby4v5nIKZY4/xpv1ffkZPM4lVIAtpt1VyUHmNIqnxcJYKCE33ac84bEyRCFYn9+wrwt8RgypZ
0FKGae+NfoDiACM12raHrs4bkLk+cwPnNft8SERUQciRG8yURXl7AP1nCT3x8e60TlzQbbTFkBW7
H4PwzDUbTTyYiqiOndeZGOANRT2Mss8cvxbtFwfr0L33Xh6xn/VuT06WhdWhqlruEhvdDcOFX211
i+WSXLpOnGBj+cqZC6U/8fWSXkM69GuPvdk8/Bhwf9vDHfbm5DwSxUdMqwQE8VWDS/NJtajMjGTN
K4BArkrqKR8KkTIDkJTNeD7orWNtqDaavT6OWwGMC4Y/wAWrY2YfVQxSB6mMGzku7ywEUmEZkPhs
HKLu7+yuwaboXK/RoAYBKMX13EDPYEdErVNiHyj2es8FtDK77ZXHy70+5gg0sC594Svb/R//7b+0
9vzbjpeBB1WX61IWCJZC7V1iJxgel5OaOldNXYqt9cMAAmGPiTXWNE0g6GVFfe1sWlw9fek6+IMK
YF76CtecQLbV5owaSVRnaaSf3yRwdFKdLx1R+gS2ux83lDA5Q3iXpdWdXvbv5YzLVJXWFiTFuPNu
sCZaPAmg9ps0lregFSNgxBF7RBk50qqP/wyymmBrzVjsGWAxIMwR5WLKnzWc2D4AxHzBwf3C/csQ
QuB+8Zt3FvuMKFi9mZDr7P6nV0wCQJxV2pgO3LS77/9DRgh2m/q+dmFpNZE+JPBYJWKG+Jaqd9TL
ByHil9yvl7c9vwa6184EgF3gO9J3WA85iT/kloID/9EecV6yIBi2r42iOc3ZT5aj1rWCtpPATOrE
AeSRLtLmXoUDcsjQM985Dxqjl9KLgToIC+6myh036jtsIorK49hU9eHmzRg4iOQlTdm71e2Vai6g
lsYTPwRXxoIf4MKEktq1rrNSPU+72O7JUFa359I8j3JuHcYzRUOQxYMamB7CKWjro0YkS4Oer1NK
M8vRhbeDK4WMSWUwTI7/UEO34QKvKtJqAcZABGcxPsXZMxiU1SdXKqMJucYbmdjnXqggjeEXNfdI
kbSDvc7JV9nujrVSzJv0oS/WFVSMGaZ73s6wIKGLbHmU0QNfXsndibnY3eo40cKSNgUwPMCROVhm
pcju6gJuwpjSVB+xIqoNJ+Qk6XtsQTV0lqkS3daBtkV2iglMGH2aT8v8aGqAeIG4RCYkEOuWH0F9
fn6yaY2fiJ0zKJpzPuzzAvrjN16zSxoyKeye/Xno51+64bW5vW+bB7Dw28TA6Tot+naYm+dcvjlK
wgJO6NxU8f7wJDmsNx+xeoM80MBefMlzaoKs3d3k5qXjXL/wscEm04keQ+zpNx7HRB7IY7Irp0mk
9lFj8uMUa3H6QtnPln4GPzKIYFy0gkR+JvqbQxSDs5j93pEAIfoGEYD+8L4RU5lhIY636q9rKyqP
pZrHXL2WHACKET/kP05+MOL4Sz36jO1Ci0/aG7bXxx0eKqrKUshyrXgrcJEJSWAgGa3/nJNUpNeA
+UJn37FWS3H6QvIqkJ4xHhVPRnf19k3bJrhIHVUYrjxFolEdaIzS69drRnsFy2wCv+9v0YbUBtTu
ejPa2qsybf/Ber96tZGF0hr7RBPrzfHktkr2XOkfzvPUsoh2OcxRB7qZu56DbfJHJ8XxV5TBLX76
BcFwCCG12QbURNwqFGblZOx4sY1VbQ0L+Y6C4d7I5qx7syNQATFDqmXT/tNdSglOsuJIDLku9G/j
sxNlqMvmiczogEPzcQVkixWmqAYE5+nI/moOvH7Zeegw8ZEi5KGV+B2vNGUyuVqi+DYjDBYKZiaD
C0cW0U4yz9jKUrW34+PfjQd84Ey0BxIPFmlSFO3WUs6FfKKUWQuqj8hSiP5YWUMut4pJN25Hv1r1
y1IzE4l65A7R0m0HcSQ9bXFSMNlE1xStzFr4oLcnmGGPpVJNpYhKDq7b7W8v/C9ce+0NSOuAkm3B
Jr8/k8fGeb1YjxuH3HrE4nIlzYtjNgeF/Nff/QJQhuzyb5NCvX2RPozp5G/axMM2KyoB9zZiwyFl
RcV/Cziv1PsqQGpeqylLzE1fHOnMZXd3s1+vffvrdu9r0R8QmL78a73E98MiBFuQnB0cohz8EysE
WFSCLnPjsSpNsjmSmSqFeuXbooqbC0hK3nev35klSruCRSoEQfaR7TpB4LreaDzptj5TrZV9Idf1
nwsMYz3ujFOaUD2t6htkA66xWt5RQJZQwRnqfEbSt5+asjDkb25cwM9Sogs30xiAuZdARzFaXdub
qXPs/Y+VfFaDjFCuPIpsPbn8UKVqHoHORIYu4wbpfW+Nx1zn4eIWFN3SRzEhX8o28dFn/9t7sh7I
Rr0b8QW7/96VrLhSwlpuRbBw/mj4fX54by8Lt7bgLACIIApS8smpfh/WjkOr+HxjEUREcKWJzaLx
NEdKwWwS3DzNGvEgo2tB8hUH4owHMJxna8qeoteFTz4LuQCXbCqvkgesjEgS1gybW2jc8cXdMFyg
Klg1DbtGwVpq79YWc4hDzsYcg9FDgTtj4yqAdh1ZHnwuVWkmbejGviSTNATQlmmcIsGIE+5oT13l
+IZ5EpgLHDrAUH4nxOxVyNQngK1U5i76y/hU7OSJBMIILwMOP6gO/Gx+lscVmu0NjWmCCuUbsT3w
e6Pef3sXESPEvh03udLDEYvVhlJ/eTHTkz3RST4t6j/jLRQZr/VPpImjwFpwIrgdyi3amuGcjLHV
DZwUMjIpYPitlquADH+G3Jg24le7ivkWlKRNQtKLd5wASPZ48KKwvAeqq857/UFW05iFlHkO22ha
TpJLaw2RBIrpinTRCeaF9qKJmrMzgGNHnAp7A549LU7kVY5y1cwomLVQ5j1zvCPDIO8KkFnZnJA9
Y7kXHXw1GWFx5bHWaT0Bn6kI3LhU0EgPjCMGusVPUhETn2rNu5FxDnmMoOkkSemsVK48Ruejf3al
ePXkyA3O2JZ82AuHliDMFAbamEZWwq4rJxnZI6X/XYflXOZUebpwax8D0TXu6Ksl5YbZOwMa5b2s
QlcLIlasJ2noXmTPKc42+TmAebTLR3im+4BHNNNgWTyUNc8jxnKdEuHWhFyHqDdFhjTo2QaxLsfs
wrg0+XlNflYRdtNWsht1dt4jcqwrOrfJtvqjw1z7AUetc8fW6aAvFglr0n9l3NEvYT27030IwL6m
/u3SLaJLLbClU+q/YaqZxJCE9FmdFXgVrRQ3ZTYWrEFyfWSSsSr672ZE18q7PUv/pn4nSB0sd9M9
QwACyETlcmrXZTU9K32iN5V46A+joUC0oR//y1Fk3wrOtRK2m5Ju2cBAS29QKLaiql/2lfWNORUC
WAyEH24HuoFp/3RkjQZYpQOR5e9Zv1hFFA5YbjtdZkQofwE6urTvVcVj+P+3JapVhqG6+c4ruPO2
kmk9owmDGvoZboSFLg8GhYAif4qPmda7ltvDlEHX+T+DlL912/1h7STLqon2A2G3B4oxl66YhsEl
jxkDpVlNWJsm8+DoTLDYRywtUSU5/unbAyfIhiIpndV7l6E0Cp2KrdAhywH3TjLGgK/PouRf9bBA
QgHE21pFBu6LhoOQEpUGkLfDbOPiZKWrelXeJAg7mN+XpoD2ROhIQgLj3hejOS8ZNSy31KPHmV9n
YCVt9VEZdTu37qqb2ei0M/MoxO63Hcxh1eOt0uxAoYOPeXOpEh1vAln9I9W+VYK6Vcyc0CsF0Q0+
HNYq4/xmuTULHEJarOrwUccMuXXYCrbS5yP+OS0p7cS7itnXNWDiTjvB/Jaf4XPDVkmoqi7akxFZ
zsR77q1Jluv6xBiTiCbTJNfYqn3KAJog7ZG6QFSq7dmOGMgzQ9Spex/CLp95ay9325S0nHljfoEF
mXJeyIJgZ2qo/FXHlOsg6wMgbd5gxAO9qTUGN0ATeZ84IWkxcHSgcrtncmvdmOmfRHfwpMPsjCFO
Or4Vqr9vYKXS5w/wP1W2YK+HlSY78GLLkBsXueILDxFthQPpc/YAsINUTIOXKe+1cWKy8G8RkoIp
OiK/zGO7gDaj5XBp5vYHm6Q+ZXPtiDRyCSfLWWAv3YlzuHEKdHuOexyH1+paKnj2TmOVPBKetHi2
kzTsj42eD8MNZvwDwWj0srZvDx1fhghlCplNYdRshWFrfzyixTxh7tZ71HLjA9vsNj46VYCfbpax
vN5tVyWczXc83y11cCrsS3kj6hZB6LYGn+ZorUPL3d5GSs/fFAETuouFXW/Ph8APefxxZO/8fmli
yZRh3AVJvlpDTCaNh0qkB5DK5+wj9/I20T2WXLMaFbCwp9AZRYNgKGoI8ltNJ2JF85Kr5LxhVE2c
12U2oRycctx2PKNV2qlsxK7wkNvQtxxF7+40Oa0VE98nuo9ET3POcCVKp0zhpqolAqLs7kLMLlyZ
BHDFcv+yz/+qcTNUReMRuzCoOnoIjdI8dTqznk4FRs0M4MVgb/8EPBVgfUE4I1HvyjNTFucmteLp
wYsmt9Xy1xxylVtcWBFYLQFhDL2ki7r0b7GZ1Yd8ATMsxi9xqJZGOrqazWaAvanUnuTV7d//f18g
yCbVxnsvakJknoAxwUfPh6di0z6kgJlkbLb9ealukmJ4kOhwysFHFpzb0dQlfSMNnBtc2C8QMs1j
MthWeHICBdBln3mBRq1TuNQg65r/ZqdUfjJgEifmSdP4rN+CzbxYZqwAGIYT9Z29a1K6tyBHuxfX
ijqg+QT44QD8Cf1ehTO3AZEOA53yXtIELT9KwXxhE7B/4DyTPC3de6SbimBdhJHIKamrVSYFJGNZ
us0OSPJF3HEe8BlB/VY53jUZHwsCJOaUYcranWAPK3wL97LZNxb4whYHxW1S8Uvt8cToFefzO1tC
7w1JJ9urSoZB4RgLBdUMYCGW1v3cdyGNNlIp73CqbWTvKFIOTE29icGzxFlaONWjC+SFkN6M2zVD
CBJeN0TUioy6v5l7VsyVC2j2nQyYGkcyZdJFcgKmEMJTEjchCLSOIm2fi+czSHvOwF4ngh9pbSv2
Hoc7iRoNj4YBA9R9a2imo6CZmWJLnGpUpT1bmKDw6koTq48qRg4Uwd9PMRGZYtvF0XdP9fYnS0nx
HIQLmWFSxR9wppJIxHyf7PXDBr8qlac1UDFX5crrnGa0V68C9rMQkaSjTt2W9mSOZ6qQrZTWKUZG
K8kVikHlU44af+zp5RpDa1AOdjlkEBj3vr0vMwwoCeWE1UApRND9W+HE466qlyYZ8p/J9TUOCTWA
eDhVeypYzW3oDfVgUsbEP9a58/gaY+C6BjMGSpP5K+icGI/KElFehpVTzCGb5NDLCsVDfnkhoI0g
lwmPd8md+2249lahtS/USsummRqFiPlgCqyqzsK5KTS1WVDqJyg0fwUUV4NRg2gzcVdn19+5vUf0
jGAjcCzsy5O0Xp4rHCAkEmBzNQzD00TLiIJS2sDeCI/l84PXgPt2PK2YMNxNJNl6YQ8p26jc/gc9
scrH4VZr6yd7/lw25+wDusAwRbId6Hwr+WAE970L8CIQW98DKfYCL/d4PYieC//4HysVLw8iWrEl
PbVQBoaeuHYJ9iYLHN4WAuQDvmdNHEl5B/2+ulrPWL9e9UE5Gid+p+VfFb5vo6G17gTQ4tAWwG1+
dGhtS7j3i44CO8/AG+wU59QwV3xpELjD2bLM+eFZM+Zc+p0NoIx2SjFgy6Bn0YpAyefEmn2Ij4Y4
S8gKTTFmOX3bBsSK1BJt6nJPDV8RbLK8crQ1dqHQTVFt8J2IJ6DdeIplDo+GCx/DG0nY6GtZ9MeF
Rca+IkClFVG+f2UyFg7E6HkXSS8IjeB5njvvlK4De3SB7bEJWnC72/qwai8Qt4E/ETIw5AylZ0c6
LhDOA15fqB/uj9dCr19HT+ZqelE5RmbiIFPgpQaVKLkVjvKxJEmxJSdRdeAiMvcB2B7KgzEHcxwg
THF4JNDW6rKKaRS/jIlothaAiHW551A+bIUF1aQ63rxykBx4Ah4yjWygGvF73PGoXz5KVAG3qf73
yqeBK90iHRZ9n3GlZKTm25BR9qdTNUfgsvmdrLwgeC3h1WaNjX+SYbX1InzTm/8SkFqk7SBSvKDk
E/r9eb5HY5DQhx4abPT2K0Z7CIvcO/N2PnomAt3XBpv8z0J/zfSjdnF7wTwBw5vL4LXUgvMbONNH
BwP05vySm+DBJfl16oPGCyjSla2ANlZP7Hz9+e0z/mL2r5tZvvQmmCshuziqFFGU89d1G0VOoqLV
i90v3v9YOhDNkV13KTpZK7g106KRiPW57S47p/WGApGTrzeknw6ChKvjaY9F5nFHYR/VVGr1HvK1
8+RfQgC/e0i922vGLI22NKV1GxZ46XjNMsMPHdfxf2DeyWJKshhPI/wsUKTkEDu5diuKHFGi3rU0
qgNUtzW8XrgtPruZpvXj8gMwkLRxzTkr/2xGDzqDDfc0TMm5bQbOHcYRARawgH/tZi4HLRWcv8Qw
pbUzoB4FsaCkFSoanY/jtFOXlSyzIoqB8KdzVorZqUSodNWxrzdVA2fV/083PgG/2ToTPlpHZW9p
FBevuTNHMVpowBfccLrq1TBXRLItcWkesLJpkNXpVwtZVIacTSWXNReT340qB2TILJQZxVGi9hoR
mtZpGVaXRulwt6nlQsKRtNUozRb6zL+ubrZRDniVdiTDwuYo9bvTLVuZVvdvGOufHvqB3frjLZzC
3nvZLCI0qzD+WkBSeGautRrINy0Iv9TsQp+itplb2zlU0wB5qgKQXY9Kg/uD1VbuY7HhrmomFa5a
XcfrmoLi68VwTUuQ5bKGPhfHOectEy53UbnAIe5Uw/C5s0c3YZugQO0vlcv5E+iA+eEn12oUyIqp
pnH3YRjGXdjz6zhD7ACoA8JLnoYeVy/Ye7JqRAWQTC9pju46ML/C5ZOmMeYc/UVgHKt+7ESKj36l
Xq9jRmNXoUXdbHHdhmCStqe04u3iT6906gsoaHXDfHWYiw47Sy+wWmP82K4KA/isXyRG0UrINl/6
Qao89Mv6Fqot6GahCY8v8SxqTi4euQwFUNlOz+lanYVghyc1H4yJ2E0uIXLVFHZEWqWuJf6B+Vem
ecvpAkGh7HX9VmSEXydtkPAyvhuYFvfLooo7T+ZXFpkTl6vFjCcDysp9/BAHDRGjtohglSBW9pSj
+872c0L8SWk7kX9JplTGL9k2THNB+cSjUOaXc89u2pxqT/6p9J3pKOYExfsYaKehCqi8mOJ1uBm+
6FvpXQH6jlKbxLBhg/yVlhUBXmSisKWJrwi3PhIraVSCcf4iY5PCxWvgwINUiv95Lw20T2ucpoAB
x6OeVtTMm/DytmkVrhUa1RVm22tXIfUExAYbOIsjpgOrdLmEijY12K0iJifo3G5QV9KG42m9P25p
cLCi+O4k0OIsTZM3sKdtA1AqX4BAVvljE9Fv5cBeKkrgqZv0tkUra0+xSjM7xFKZBXlcIsCF3jtL
RL372y8vKqroDAFZ40vTBjw2Bini+RPVYp59MSESbO/Z9XMUeNinKbMefr2BmLpAqsr7msWjiTxQ
8BymqOaNch5aXQGXWKCzrzMSfcsjm+WCn3amIt/EXpfyij5Zlr+KzFat+6JzXmCUZgn+7pApdrH/
LMgSzvEh72Gglg5Y1RvRMgbL7FMRafGb0NObWoe70SkDeItIsl33f0jd5t/tUsy7nfYpxhilBuYs
dqPpbFBk7s3Y3xhFA0b4wGmPgA+oFzNUZssrm6xI3EjGZgVHKcFakE1eOwnajM4LczkJnxJKgxeE
beFyhNmzHb0XoYz0hOSM3YfILO9fnt+DptxjxhMmARKhM83jDw3aQ0hOO9LgXmJuScO/gv+kr4qt
f21HK1/10w8zZpj2ParvmjEiqThrNJeCoX2j4b6pW7QlgHd6jzQW4p+gq10/p/OwGQssWKjX8N/1
p9hR0AXEvWKcxl7w3//jCk0KLSjWhb8TNJuOlvfxbONoAAKW0yv7PFuIqJW0l4SvNthU0/gE/XPu
Q4heBakf3KIN9FcrWfBfab8p0H89iK0sFpX7dKAzfpePjlQfGutDpV7IcufKw4/UH25VAyFqe8U/
E2TRYH+vCYARIB2ebfTRWH2pT+9Furcu5pdtoZpDRi6pBmHu6+iq1FysjztvwDP4juVFVgrYSVla
0pvhOkgBXccVu/SaQc/ocQv170ezbv0zSudOt5Xy569Mvac17jqQInkZJMMgx93/i+/axZ75RVod
UgF/lWtf81cDdgPsQPWxyTath1fgTln837dK9wr9njo0GLyfGsQ1UP6Z+lwIlRD6HE/8PM+otAWN
ykCBKMW3+lVz6HTw8RSwDUqQKsYaEC99cJPaeqO6fw1FYNMijxPdqroqTcdJ/j6J6CyWqio5pUEk
eVTaygVoJAD/gOJygvPqfj8wQ08MsgEnbsX145gagvyOGq2AoTYw+aAGvuF21FeJfyU7A34Ogxo7
zqUa5eKPG4WsVii+irWq/w55a7I2yQ+QOJbY4Rflvi5+Ers6++J8uJhLkhPchZVhH+UWn/iUPuJ5
ZgqTgY7YTRtlX7DIqoOgIEW0WwXbNmvjTx/rza7C7n2zDff049wbK6ZYwWjNbolAYMRaXvLDDaTO
/Dze8Nj7/1Y6fR2jcWq0jnN8zOH6tBzI+JIQAzr5tYwh2GOVICZYhjTjDzUNmutTICGNRzv4+Kqh
ci9DybJAGREbxL3QCXDURo8sPT87sclfyTF/nfWKExkmHZVmaWVFv0aiOp321SNWbcF1qyZv/Yom
nnDt5+++9VfRjFOCs/KpuHaFAmyFPF5gqNKH4XboB04D5srESQymEhqlJSWc6RWbAeiyp/USxN1q
Vy51D9MS814opAi4xJNGNq1N4Kq6k0J0iJ/dAj/mlawIxcw3BkRdYGezUT0E0nvFjbmVV8MxeDGm
fo/sadUbE5Sai8vHDSzw4ir4RRIXMxGO397b1rBpMNvipu7IZgcMbhOccIWQFNgd6PKcwiNVyu8e
FnrF70y8UP0DP0/k0I0AJiDJsl/wp5qvGFzv9XliyReahzlXCb/cAayIdvomIh7MC8iX4Jgu8foN
bNkLjk/VUCO8Ojd2Z4UbVlVBZJHNhtPyLql+z2Rso/DeSLqCd5gxZmBm8oztUJKR/+op0iTqF4K2
RcTxtsUv8j7l7117cmDBkXiCymoTeZ0WO24RzlWDffy9qS/Pi4p3jHSVfIamKWWGjRwjsBhj7v8T
WAnFBQljW0b2om97G6LJ4PW59NwegqQkNtiSyebOWGx9v/IsoZHWho1VPAvqgICTPHVyY3abuh40
UpyPbwfUbmgmIh/eyjQF3L6SQkFRqLXX5SE4idvBNuaUpmH2lcTNlPy7s2QXhEB88JajyQFFlH+k
RzKSAmMNWFKXQ3vTJ/mhGbiUY4wN9ikNdFTQ18vhLyQTzgu5fnrA9rNRvGTbrt97/YnlirUrhl++
/LUA7PBE/JA5y2gUjX+99eMhsY8gG4f92tpP3H/+28bvK+ezk77Grw1KrkLaMaz/8ZjUKnnQbsA5
b+Zk0ps2AdcedgmgrbTicIKmUq1q4vTBNt2CSuahY6LmpqmnUH9q8kil1VDjgqRqJfawHrv5km4U
oDIQXtV7Hpn4efsGv+LdkG/iXaYsdgKpSOh2j9iBBj5B7mu3w1wLl9qUEJS12Da90/qko5rOTqmt
zGYlcyaNVV1jYiF/JFw8rAnS/UDJz5DBLVLtlsmqUGdsCQPk8veFN5WJFKd9Y3OdIpuzR0SD2FT2
rIIaoZefUVJqwuhG7XJSMuLAMn3nafilLWHzD0KlCMWaNWA6bBvZn+Owpc5Zje9cfyJ0LuElrcxk
vtsVsTCYLts/7aH//iW1xcPHA11Gimg1IDOgLip942OESDJ5YX+ra35tLs+tdIPu0W/xPu082zcG
GWYz/tCIdgc42pavjNfhiifUa1p5cTjbT7mor94rYFmX5nd6KW28qLVunN5VTI3VborMKWcQJTxn
iY2TDgcHFu6Z5Qa0FhFoD8WPCaofO8wV8E8JUEDrtoiPbpnd7EmSMOdCUPYjYvp4pWelxJqrWWbI
/1ASXNfYd+MbhHI+/hXiyR8OTxSQfKTk1UuvFKdNd2p4nHfVRZMsFXR7DZvygU1mimvQBOv4XdRM
GUH/6TtGCizS1n7GMYxmial8EJtoUbjJWY0Y+3ly6sI3RLfgs7eUaWEskkuOWielw9wKFNOV4l9+
6+LSrge7xhKo4G+RGdmx150Dnd+kr1hQwQYcUncWJsXT849nNMHXhou7RdlviJGF5zomjYsZ/VPY
Mevl1lvZ1DgHF6cy4NUo7uD0XIAyxtiv0vLe/ZIbF5AHdirRLr9nCtpPvs6MnQaJSChu/2eBNMPA
G/B+qlkcOIW7SInmvet9oFmxdIo+5BICuvidDc4ncZVzJkuYjmpM8lHko8gGDtNopNpZB7Di4m6e
ZfsRN3TzdSsvrt/7Y25oGUk64ca2CPGaxGsjR7U5NYKQnv2Xle5fgE8W6bY96SVMiiSG1lsTPHr7
vPDmN0Epy+mFiL3pl6TF08TTTSAFBsIIRMZk0uQSNogCgp/qFraqdETkVAwxeukQQLNkrCaEyJK6
ZbqJbzbdxJbFYSRLoFy990PchW96zLl0YGUlQFApMKwigyGOq/qRT4JMU/kic4+zGZbs65Zxo+Gt
zXt+GwwbcsXt/RtM8japEQDtPrSzNzRZrIufjm116PP6kX5etri7LMk/4VrTKnwprJnZqgMxoQLl
oGuUVO4iEEv3lz51yAgp2TAdSc+I/qpF4aAPdwdF9jQOFAXfEIEt+uB/QRahPCy9/U5s0464OttQ
w4+d1v7qqWcVINNUZXcU5/UY/u805XRQpjUaTVZ/Vfj6GU/2Y0/hMnJjHFiR5zPkZAdbI/tI2vTq
nxFRgtx6tGJKNz3MCUV7wdufFyUV0z/95j1ZcdQWwgZjYWvTzt2JEveCptbkYMamnhNgHv/nvtOa
e64WF303v0a+LYMjINYgQyOTqBCTbMvlSyoxU/FCpb/2PBwjVuKN5m419DRGh70jsgaiPlDXtSMy
7YskzlE1vmrBSJ1PxfpMXJXfEoK9hCc/8VSKeqG+iNViR0Lhhrq8lapgN9kCooyoo7wVvdZwBIEX
DtMEDjp/nKG8DWTbnmHUfPSoeG6bwfJKml9Au2mZ+BpcLcjEd/pkQoOdQz0o6AIWZBwC3rBbO4af
TmTTi6o8k0xvCshSrOVP5h6hzvzD/oEFzdLvZX18mxONGzrcxxPMmidqg2gbiJhSPa5cIBqJEtOq
9DyFb4BY5awJIkrBmiZt6f4MnPy8VVvmt70gAR2ThvHEwGJQAZ1+pOkfHpk36LGbpCVImc16e2hR
gweq+AkaV5LfuumcJYWwyGmNc2uoy1gk39OJcXvmAHVDu6selDinJuY13K3Yn1A/3PO6C/lt925J
/Qrm4fdH1dHf65SmHnk9KZhXYVnHYR/NH3NMtgXQrrfUhnL6FrYKYh498H8kMZKNVKtCmW7RXcyi
x+JVjDmevNQVCEz9535vWnuTu5bIbfvt08Kjo4F0fYoWi2QWIH3K9To+Zkbho1cRuHXjx8CyRQ89
t5kDp8Np7/NiKwRgxy5a4g7S6q5sOWl5oe4F0QgmEAbQtDVYJqJ6iGGk28lyGnKlNUiUQ5W+9yx2
AB4qjNA9cg0BiMqw53ESOQFFSRxlDXhXa4KSRa/iot4aWxa4g9IwLjeGNgISg5o7VE/Q79RFC2uM
V/cZOABHuuQ8CdHEKuuNvao1qw2mqsBp8WME/Vo4KGgpKqzGzOiAFABtCdirZgtFx8/4qB7T/opx
hEQ+sMOSut94/A28Y02xvYv96TKjFczUOhmtvyb3vPAmlkffqzJGDGYLQN0nQwYjG9BOiYcba8Y0
91L8uZvlhs8XRRBJooch8UiwLZK7LZrqqrBeR2EacIYmLzCZBqxhQr4Ap3gDN+2geB4xg+YnbchH
UmX8RGsunNSedXGyoTqseCpJ4nImYk0apQQgwN8UNosexRAD7xw/EONpXa1f5ZKgKDjsY53bKIO4
C3yomuoWOppI71ZdFKhaKjzo4saLyEXaIHpKFXCjtWcscWydK/iEG7UVBDOLArsj478+VFpfs0b8
4CRjA2qqqaDynVwMZleXtTWoXZNf2SM1v7NuOWZ8b65MJsqNKlrO7PbU7o2VgrpYz9p1UU2A3lsF
Sa7B9LkmCR/gIhCVqIU9C2TeCT69xcaaAokYpVZ+Qiqb01rf6SSz8qF2PRaLzxw30/zk8sjLvyAN
/kPiRpBH9qWKDIkLBb3MMGHPNvLVLUzCZlq+DH0YQOdtD3cJM2c91ps7CIZ0RCCK8VADeujFPivW
U/9UKgMxWuLlRp07OqGTaMeCF2DUWodtUMJXIcSg3wldMlenosvCanjl6feJC1or0uvlIOQYLbpI
F4t4hbH6idHRJdqMRiq7VXXJBXSeZ+Sj4jF33ZHydZbiqnVS3FHazfgBo3F98bsl4hQM9pKcM07r
j4m8IK8i+g/6kUk1QuQTQpFB3qM3ikYJZ5vy0A+KwT+twFl2MUd9WWQnaSYJ3cOSJgSUwuD16Zya
HjanEfSQlSE6QmYf9m6egDNzz9eP14hoNpKMuHtMGfCqeNX57sZ9cmQ6lvUg+vKro/LYZjrnMS7I
csoX3fvTfRqun8xr5L2yr6+WUFNxynaGWX2nCmVk9+KfuOIJ4onZmpIrH6dUCDHm9upxD5qb4Fcn
WGaDpjSNdj0ZyHMMbKYqr9kSDmE2fHINW1DVqtjzPia9ZwXIqVTxKE9I0EaUBn7lDGaGZu1nvQ9N
QhxP0U4/K448PabEOr0QFCm8G5CcRc25Pa2KcpIPOcHtrpgeKAX5mEC41+H1MgABV6iMJmFLn4Oy
Gu1gt4fGIBZ5Mxm9SBAmu2xuxpWfpz6qt4v7l2Nesn5SxShLcQPdkRv6/X9DMuXNy47bb9dHzMjF
scknlCo3XMPfV8LPy1VyemcVp3ajsgHBB3qoMftVqqGFEPBsUaht6sBEIUQn8KI+hoFnpVnKp8GZ
pvPLR2BXluLcRosrWTLVoEjGDGFckJwEiyKC6f33GbJLPGq7b2/iH7+zm/YC3iioarmGeCoVuKFe
1+wHGlMjzueMawEAwcOqSgZGY+zbSRBHmcMcWwetpgXdfHe+24iIBRKGUfZ/DE5omXtGygCgv/6c
pInYyWlkTW4bSoIRsoDUgVnX7xZ4495tDMEcyE8HF0q6RfebgUeg4fsGk2YmTH3qrdcWzgIxJRux
HEp+NpsvG3db6siBVoccZrM9bVe2fZUoOJq2fB9hvQicKdwBiyGSr8OQBBUqlcp6K5yd2EYD+hSI
Q1JkeIp28ibJ0+ip68rEbu+OYgcY5H5hMiC073iWs0SVd4glJ4E3GZ/2cY3XMoVMbYa8b3nnGBK/
M1EtPsh5+V+l046FWznFV3gE3oJ+xjvH3qOImdnWqoM1fIgp6hB1M6W4HC5IcHnm1i6SwIpsMTEn
3aW+B9gmxfk4D8E4f0IJm5QaqeMQHL2b3wjGYp7iwrV5vu2rFOXsmTaaHwyZvhEfF3H17URxPrMz
xgxvQ98EXe96W/tzCtXW5MBumDMv2SqkYUt74wE9j8gbg59uxkHG5mKZZTOceSKsvI9439n9H7Df
nKBEE1rpKF0xhWET0BqqLd76V28mPnwcvViMX+oazX00jhR/JaiR2j4zRk2KaqQ+TBbZAHB4aztb
S+jNn1FklhLYzRMb4yOUP54PAegqOqpPKtUSEOiiV1km5LHh7ZaF9Gz3DBLrul/ZXxH62LN3lbND
PJNNQlFW0B/dfdEWCpuz4fYZgdyFaVSl6FNKk7X15Yx4aiz1Wh3pF6Tz8Zg9BSXaVgXKNQEJXZuD
H0pgeKWoN5YKHxOzvxzkrnKoBWXXnJCw9/v+CelUIAj0jZLaxZSmqB8etLYnzQEY4ttTWQ4bRj0G
qjI7CQHpxUY3PcD4CpWFrxwP43YktGYGJjGka05bzTJXPKZmdpYJoygRSBJomrMMd9CbVhm6X3zf
LBPVitwSMHcUPZ3LYhUtUGP/bYg+ulxX+Bvck4sbbgftlp+GaKoEyQh4zng0fD7slusVt3AYaoqp
fAcLn+6/+XkKyUlIshSEzpiSHuhhajXJWsPzlhohxmGlnQv8qu9mNZrOPOdWdkwZzl8hJ9LKkPJs
vARzmIe3CbmQneL3q9R56pAvlvXMkFL8EsnNFrltupLADaMo7UNJC6VJzVjHugB8eenMNANVZjdB
n+XQS1uZ7wLQTEiI9JyOQuJgtyfr+vgfmREEPSSMDidRJ45M90Rlq/v3bkEMhkOc7uwbx+UU4nzF
+apdcWrBa5IKL3QSiWFIatYcnZmYUhpnDFB4sOGpfmi0av8j1jcxO7lznB6b6xQDCIobfGAZpx0G
9ITdJueQZcQvN/ZzOBxNq/HMGUh1Y3x2k1ioEMBhMWzN9fAiQbHBeOqQOnxbsOdInIgQBE147MrZ
v+0UOS0eHa3jCtAySWzHD37TB0u0wsZ2tSViPmus+1Q6e7G5odJKY8yANZEnR6ohUQsiioOK+pZ+
cZN2hnV/LaXyxOlZCVa6zozORCL7QLMm2nM9yKGG4H6y5T2dU4elK8M8ePirsbd/nsDKLbHKhy4X
dsw5xqsXVbXNUdXOR+/dc1hgNIi9disXcia39Xt2cdFjcEWAIk4Nbn3K1S/QzS4ArKTKdrJmaOOj
H0LYCdv19BZD71Hfzwuv3SJ8Y6gxPIZ+TAmVZldwpIrEJy0+O7iRhjJrvm6IVLbeaqwUW8XCsLUf
TSeQiV7QyoecSnmdWU+GXrgJ25wqsplnDyO0bfdXYp3awXs2ue9uHVD9wsfonNiPiWD9eqZ11PdE
oQmogEsP5mVdKHbUXGNRHmIu4D6XUv7CVN5hqaj+8VeAEXqesFp3RBGVzTpQO1LoNSTkS9uZ4rHQ
vS+7bE3uKwkdccSmExyz3aS3DatYyHvyQARMkwnfLwuhzElJuNdhTSVLlYKBNFxsPb1IgL/ZsPMx
okplxMT441+M2L3SGcZNYoNqXHj/lB6dk87NTtNgtbhuztwjOKRXP6RKpIcIrfci5lbPgDasd+d9
wpsyFPeZTnqw9dARpzlBYps65DHFX9xRwD1qX91D9rQW6z+R/eKypCyS0QrLjQh8YhK6LaPwdR+O
Yaxqx9FDBoJHDMVwLKd33dEHRnbDPXTOwDeZ19fL0MPPJpTxmnQPRTVeJhic7vCD59nJFlVkkB8p
6DbRo8eRJXl3+8GRO142ojYuY2pYXBBMQsr/d9mDrhNluAU+3gHOB9ybjVjD42upCrkJJzgP6ukK
86tHlEdpz1agDv2eW5W1KjOfRGr6WS29pfZ07BppAOJr74LlDpcAGvZGDiIEzUZbAd91SSHeBzg7
xU+WvCZNSDamPOVS96Wss4xofkDa8kZaoQAOhoTMrX3wzpFSqumHH0ccKrlGLi14uyqe8bB6Rr59
+tWqYQ7JjIct3qS71fHRH6H9YnX/m0ME75YMp4Y6/ZVMjVJ67z5t+ktpWlZk9NiA5IQxPbFLi9IZ
Rd6F4n2Br91JbseD4A5Z+QOPV0bTMxUkQVVKOFer3GtOEjBU7SxsHFtiYOv5GXP9AXFnRbOHfVnQ
jjip9bPdnlHHmM13D/dOCZpjF3pC4Tk5APZOaeqLXu82dK/lfxAJd5saZDbvJu5Q78+oTv/Xqu+z
gyKvh5fLrOTITNt1Ic1vyph+Fm3XLVWvHVN6vuBT9G5JRPqKMJQZqZa+CXfg5URch8rRVchzlqXY
GfmA3ESfeaBrR6zq4KhaKwkamEumRBVBkZsmwCFCPKug84zMpm8myeRdaz9ZSosFlPF09nRiFT0B
Zh/yci6hnFBN+HG17iv7PbWPMCmguT3saxG/+gnf8YYHn5j0bk7wTukgNcVB66gQjJdv/xHcl7Cj
ZQl2ZTzdEwrpEc5P82c9uUa9jG/6KRPevhs0pvoXh7sOM66NSz5c77a/rmZtllFwNNuRZCtjb871
IebMKj+dix+8QdaWIiI1zpBZzNcLrqGPaqDoa/ydewjRRkBuHQNiUeoFetHW441UtI1t5n1uBfxR
aa1yChsmmReMcPIjhA/jKbOGOKvBR3AACuRcD6neYMkKjn4TcxNfKsmNW2HZloc5veHgc+VHVNbA
aH2GBr/gPL4WsxqN1CDufZsJanwOLHmfbXzJ59zZa/bPdycIUVb09Kr1hGdQ1Z/m91ezUelCQOF4
SQOKkxtJd9j0djMIGBCQup165OZxkP/B1MFx9Yr7cubikQqAs6aoHhveyCaettHqC3B8LiiegDFn
bUxGOi0UXRtQn/EGJv8VuxT76SkxaAEGCUjTnERcrdq58wNktFhtSff730VB1ocptuZQH7Hu8JJb
sMfURnLgnGpBjrBCSZjLGtANTJkQ+YJ29LIAAMk2iAYgEvxTQDN9qBa+LcDj6RFSjC6oQBJz0ns5
KC1BiHy+KIujO7WHR7NFnn0/n/snpd5DkHczlHi2OWzF56Gksu+k/IHD/t0HWogh4JThF0t1UaT3
9rPwi836Fflp17V91eT9qc9ab1Uw98Va4YbbKdUykUCSBCWBXS87JbHTAu4upPOwEHOnhUDZQMWF
XdTDo1/vcrBLisRSyEmLd7EktpNn13Q6ZRcOg5mkHHGkPN0w6c8QWfWjM2wquOdlWTMNY8+dJfCK
vmbjggjcmh1cB20uskzl4f5q9LmzcpvQ4y52XYw+NIWY3F0X2weQRaaQhpcUh9NRbQCTrQTqBO6Q
oD1v5KZ3qcU/Evu+nx8t0P358kIWQgmwf1tAVQLtU/aciTUb4ciGooiRk6vfbMmMHs0C0WI8aIKO
0IBQJW7vX6W+DNkal1j+JxD+eixQrgA5sijr7k9VZ99Jr843k+A8RXXxbiCvil6LSy3KPxV/1JD1
hqFhWpZ3H+w7V29Z/vqdjO+d82tzGkhuZ3azj5xtw6d/AosmmbCU0PFAIOsFjsBHGcaJgmA7dqwN
XULDaUXEDKKEzHzpKYCavMAfba0QYiXaolsJJMSuJcL57lyTMsXq0LySSN1Y4kH4kZis6WDWb5yx
BYWYiNfSVDRb5yyC9vY1b7KfR5F0TDPAuoc7y2OOG6C0r1YcdDDSgqadnoY0d28kh/Yx69SvP8Ww
IIgE+lBuqZ/E6Hp1qwuufEkgqkREBqtcPGivdETzzSyapuZ+Apf2wRTYyFu7I3cHxKQpP2+UvvD2
kWz+k6X5TEKH/sXmPfgtl+zo6B+bojupn6it4F/eK0EcBn6LDxh6kRvVuyvELx5/bILyn9iR+meE
sQwbe04m31LxXZyjiFowyn9gALNvwFW6NfawzoN7iVcgvXJJcsesKdMRZIHO8d/1nESjiIsFBYh4
I6fLmPSek26OFcj6TMg6hJvSU1k1jnw8Rs9RR/y0S+QEmczBMT6Ayaz45Sn1F+4wkosfAqfe++jA
Esnwq1mH0ZlQW6DHDZEDSMF+M5LRRUvH9ub2CldqtNdFG2o8JKvVx5kd44VhJAWNKjFgHSRPiJll
Nba+WT6BhkFXYkmY3FqktoxX3oFJ0YvnwPQYcAmiFwA4W+XNmeZgwI4NNArOvRLvwjlqeOk4N+MZ
9qYGb3ZlPOtYPCzFbXBRIH2cv7P9YYbiaU4ggcZtuVl1TetJW4hJ9rOTOGLCOpEUbDWJik2THoEQ
uzLbRd09/xC2NgCcrCTVsymD46yZahrYIwD4pRyGPJEVF9meZPHWDZL5HIy1RP4xgoD67cDd3bF7
ot68vtCmXDknF28qi3tqddDJKqgDX+lBJA7PPLmHoWuSZdkXvZprZLwR1cx7PaXa1QX4QVV+aSuZ
08OS+n2fwiYM17/h4LDUqoxI/km4r7VnYQT3fmNGeJmEWUKsk2aahtJoPIiKwpakwmzN9ckaH+eK
D8tMUUe5vz+u5cSxirKkgaC7kT5feHts2i0OZBhBYDmxoGRn0/aQT85hybBZ6PPTSh0pceCEfaAq
6gda6EqGvQ2IrCUSyi/Yh4ouHcltLw5tWw9ggNUkca72L8CdNlEZnYquQf7y8IvLYji7kiqf56QV
8oIlTbur7p7l/Vht14baplLc3oTHsvG9f6qEzJZa8fj+318oAu3b/w9u+/eGpYurqtnYqFH4lA6h
DTl2Q5M0ImYmxES0y6kpvZLaXxiKWUTd9lVi7KtVf0K/TJN1d26OF5mIxZpo10u6YgE6zvN3Cey9
Jjp0IVgjcOqUje0X2mQdzVAf79fOs3xvdwqjw3SkQDi9EB3KxC95dCwwp4JjcCBpB84q7B54GXHU
ubo63c8QobzBFZeMkqwTXA2hGZ0ZVKHiBZSvNJmdnAyudPJcYfeG3VrDVmB0FQxwpGsd+RH/zYN+
VUJWMVDDMf/1AsEfuotcuGsLm2SQ7Upm9+/j/U4XdZsi0HhbncM3y+v4emNln9TIEgKzt+UWSFgz
CsPXpnnkxL+CtbvPYvISYLSs2Hlqv1yh7nh1lEg+cq7rARFCACuAf6TtP0ou7THsI5oxrDI3scAt
dSJL/fubbR7k9qnRLvZuyk5+/RM7024K2DaRn1nuQR4ujgA/S/SCfbrmRkXBAmcZKkmqLsOLWOVJ
eOTTWJBqwPwuvbU7Nn4V+eQwol0B7OHpEY9ASZduGbNfsojN6DihEYUFJuvoO3onKfDiSWmg+A3K
PPWcYzipOfQe6CzjJxKk/0Zd5SzCZRASAM5HZ5/GCqsMuABr2/nbNZYDptRdQcjjpysiHgZ+CUSM
swfAIpt2HsKD1FHulFqEYhg4zhIb9TNKr2QE6pFF77tcXOk6AhH3aDeucfGBXBm2AYvyIDlzIAgM
FRWRdEFFb0iCx+yPnzrhSUmygQkENP4iXizRXV8DW3/oYcZbc8dwSjQvWvnC2EJ90WJE8eiPAHoo
+hlst8KlSNmPgEQmef3KJ78pCWo27Os2WyulvhyrTiOCoc+vjYCdyvouW+UZPR3/WzGLGC47YQgM
H2rWhPh6/6IiD7qV391IQdkP240zfqBtPnGnpO3QD0y5Eqqj8esGznYkLKsZb8NSJpbU6nHESonJ
FvQ43+FJnql6rAReG3wjlIwfnVFgSU6eIBYDj3xptprGiUX70dBhvyG79d5KlB/PNNjEI0F/+fuF
6xs5kBsXKkNI9GjSNser+4PefrOlhcAiVxYN0ClLnozX7IHgquoIrRKhwN+XGYrsmiZ4LBfooFgj
m63OOwO9UTzt829pQb3/QUmb62Wx5DeKTe4csHwfwJ/R2ika6hgaSmu1f2cQOE/EiENK8+8wXLxS
so/lK68EhafAlSEcZUD76e5LLSFXtHQ6qwA3XNv+0Y7XJkP8JiA5BHNdj/LtShvg7p/6BGUC2x13
eyIhDIiGfWXQDHh8X75usNLz+2nTkfCO+nRFSnTH+41mi5aS/6/qQLgKu8JEDJuK9eLlacCLjqLk
ffx52mmk3v+cdemBE4VQQnkvB8lk4wYdD+R382x76/gz2Z85Rny+lVOdui8GKBZn4PRsEd5+O8DB
rdQkNzwxzUjQMNTMWjdwT91h+wyy0DVFoMUcF26V9f+4kdeo+VEN2iiTTX6MyoAUJn1DrzOLXVID
2VdF8xZfi4kGGKB4AaCg0rbpA9NTmOvNxf4YKMb/CK6gx52UvjDtKYer9UCGTG/OHbaEd0RxDSlp
Xcn0a6fyfOR/2u1HZ4rbfSHq1w0rlNLinlh13KUYLWyu9D03wjPopuEnjDf47Ipskd0ydpSBxnms
miZGEgwWKsNGcGtpNGC3jM/dxYh6iHdb+j40BPwAP9gBcbc+1HgU1Ao6OBKAAqF8NaW9WlQzAX48
ImeDzS+EFVFrvVmFBA5zzR9rAgsDu994sGQSw03EILnQbcIoXhFBt/tYem5BR/EfhYgkvy/j/ZwZ
VqmA3+CvVFMmGnXSOa4qr/AAqjtKAj4CJGQOUawKXVRV/F+Tpg6y/t1P8jqwNwe764Dt3LFni7a6
ISqrF8MfJe+yehaGj3PFMrafDM2sGN3U+KhY74KkF0AkXfXQicJ5u9ZohOt7HqbFhKlM4eavXwU7
6XdzGrXPeHmQMoKspz3w+GGPBWN++cVBtFp008B3k4GsvS/QA9HHLBkox0f8dVv2pnvimUFo+kch
oEf0KBD6hPkeG3EaQPPonCkvDd3c5jasZNC5vNG9etPwx/qWCJLreGA0zH3HonpAh+6UirJ+zBz3
sN9ta2nS53yrU24BCHO2UAANvoPxaWqmr2I1slbqLS+kycQ5pbXsp9cPijwIiuFEFKRrDlQjsi9z
l/JDv2nL1pMYtvcHMTTyqA84voyLSnckuG3a5F4HFuO/e/TFRwowv8C2uhISkspU3YXcjC7xA/oX
jmAZDZyPxNJnlkYOcxamWWK+cGabBL4oL1qYlHofkYeStQmAWeuuAfEbfVsVAf0Y68ACqwEEB0rE
uLaAQW7+jpjbI5RXX/tewRda/F5UOjGJlD7FfQU3zpU0nZK9Ov77uZvxUuKU08m04nv6O1gKPCHN
uUdhpf67LDjkacTHkGSfKY9pnmYRQd5tkD8yaaNnWMCnUNIXYbob76LHhGlTrDJZNxZwtGCVNP14
yyiZ867HSH4QZbbgR/Fmy26Jl9RwP0Q69x65f8+6xJhDOEB5gKuRW3cBzoidSCPWidhOqk6UYyfX
4yob48gfYJNUEddOxCc2H/wVLKQOM2HeyivfyaMgOd7PbmX9lg4QY1HHKvlKlZtqThMTg1U+uaTw
wd2YhwjYqG1qPUh4+8vcLRt9Q3eNo9kyT4o5T0M0mzuz/XhWw28k6M/WcQLr7r/wqrvHcnk07Yqd
WvKlq1UvtSLP3g449AMqy69FbHWzsYvX737vus/mSThuepulTiggKIRcITxAgPfxG8fZMYuAlSFF
uJ2zG6cVNI3mg1++O7U5q+AEAmiuF1JmwyK1QCFx0fJ84dFayS9phxDQADlbFCWFZWrzFO3/DXtN
QRoHWwp/dEFPD95keqEo/xXklDNbDTfixBw8zTaJKopSomD2jibedQt8HbjWWnVaY+/eqsHKrk/x
e1Ss+7rSUGEJeqdvrVgyQ5dI2RaHZOB4Zk5M/FgeH8zKnT1cuTHlQj0U2hI4NU72zKgFkoy8q5SV
w0w9RlSQw9xMlCTOJnGGZkpBn5fEjCy61Vk+f78wUq3arbPIcOUUEqMXss6o9UT8gw8gpq96SJ7H
Zt9EQPylQ3+vSAz4w5xYN9rVNApvV7a+NsdDnKsFZM3ur8bAnXNlLMwA1bJzbGDZNWvqBGs1Qbme
M5C+YstceTAox7nD7vhUHnTSYihaDx2DXI7/7P3eHzGfHV/+2CAd5dAoBlla0sbM7vfGMv2bS+UR
zQVG39c4HiNK2Wcqibdgu8gLmfEtc/7YRxswU9XiZ5m9aU/jAdLUd+XBxgBqLeNaY7+61QiD8FUT
mcYgG7k33/P9ngNcGr0Flo4+JAgcfgzs+X5Zkx9yQfxfGH1DkSf9fl+xNPixh7attRM5qJQW16oE
HTmIqzAvE17fEmHNBCoDpO8liSG/x+hp9jLyfPp5tPMObNHZE7sFqzueWYcl87cHQDz3JKveQHoq
gbt+nG7G14B4PR6wChD6UnGtgwCGg9wfQzKFuRBFyavnqfFbEim3wkDLu6ofHOSpNwJPRfzhK8MM
4xqElH06DXnxTIE1zMjCs/Bh0oaMcTbXHkF89XDn+2qnDtTUxyoaUae7aRRWY8TI5lSREl5AaX5Q
j+9KMOJZnX6tgKaOKfkK0DYD4ka8WPmgkc48zq1UlJEJ3fGM4oL2Mgd7jgL2AfTo8Wp6P+HeoOVR
KncOy2o7q2h7/mIdthNteUcM7PzE6RwZYtAAukZ/NVeqDwcixzwS+BCRjNsPDTDEmrKvOVbgiI2L
YA06KHgdwqSCTpLF1Is6GdEKTlOvFpyXqmsm53lmZYel0KbEO595AVvJHB3wfe5QNlNz89tN4xXM
5QFAPRu2zvn4TvstLEDC85f3pinLf5bbjdDE2UUZBzSr2RigdORR53Dtuefd6MQJJfYlarQj4RKm
v6p1Zp+JjJXURTkDLIW8KWsG1yAtrOVL36ozehneOjIkUjo8swwVdxchWHhCC8bQ0mBGArCFJ/5C
FzR9zENd06vV7XAooo4apybefWkgPAWjDsKjUg9JipBKoezD5JP9Ju0FVdmYoUVPbAGeA4gk8kiU
GGdmwnWXiW52nWh9CufiPNvoOViNtvECaGmuQ6uUF8HHIxye8QGHCc4fInEhKkQ4PD6sFblvkjRf
kPg3L0ljiBmwrzQE26+6GWw7pZjfqX8wL48B+bb8ybVvy7ArsLchKQIeIGxXISHlZaEhmopxBSDe
k6kZGwrWFCkI6+fXIzKTW7+77RFJ6gvcSfaE7q9A335lpzDU/4hg/EilDdVnIw68+T9q7avHe7+v
Qc2l4KVGwHO26nvFMZOA6K/OnBMlX8o/ppBBSD9GC9OUd7wr5DB8b23+3PuO/KOE4jBvV6MtiT5s
4t6XTsiPLcaU6anyrXGO0DNg3s+eIPgdUPWJRvox+ejc8hiFdwYRnHZ1WEZF6f6NwLnDIWZ/87tZ
GZmzq5jmhRJDhKAr+8MAkzxst1SVqG2NPBx5I269xmQeZQ2ITeGdctVOG1wminjaYnbCbPHQgqtZ
/3Ve7/KELfBaN6ydmaWtBCliUom2A8Dk8/lG646+O17np6K6JgLdLqfiH7sjbzDvmXzYxyjl/JI4
lkMLsm34wWopb+BWOZT3sGBleQu/j5+O6siAUL4CfSIr8X6JXV1SlHa342xPnQR4JG5yNH3wXiwd
B1E4/vo1VP1BhZpa23HB2ghtHVMYJ5tf8uOKf1T2W1QELfrEqunRgUM6ocng4ibJ89OhXCCQwtEY
fL6PtytEeqvMnjq6fifocIFOoUp2yquwSboUOZLQosmva1jnXO18ABZmoQtVeqDNmD15KEyhg4AK
/5nN82H5bC9zv4BTSAmFWKPs4JQHQymfpwIkudQKW6oJy/bT+uFuT7kgFG5X6l9RTUW444LTTMsu
BP74UfotD9H5ytZvxHKmqdB+iaoWBBegT+3Wf6zxM4g43DIRurRkO9SLBWchDB1qKVeuD4f+O+2q
iZBbRcufI3Ea2lmLvQSwPCmJF5M42zr4wHwfKK4FwrlwaCpr+dCvXmxHHndjG9QF647b5kGrCaJA
nDifT/Ec6OJUOndbDnmz4MprvCJQEmKel8C1DO/dQwrfUWDZZH2PoDkpICFHnFl3ybZsB/8nv+kj
bm3nGXc1ZUPlSwuE8dv1+zeJ2Iv1wIGzaAuoDPHDqA6KkEjdEK8tA0EMB2MPLQQ0huLB66/xxZXU
YrK3cFLclHXOYbppmeq3K9JD6DI6VKLSTSuGvPtw375rfgW6rO9DwUpPqs1osI+Jrnsi2yK/SYJr
/Xr0/CStOo9kZl0XwfdxfS4KqjM5Jx2T2bLpSa9u2nF5ORHqVxFPgXB3IhAGF3o5f5PGLNGMNeYn
rqPNY3GuSE9f+8BPODIvUavnCWK76K2GGuMwbbRdhX8A9C6EX3VzHT64JIP0YlezExRw/G1TlUtn
7tl9WsR9ebVgAOC9DL+3yu9+V41BolmEZcdASnv3MbsIdHJh+366As5lWO7hSUpf6YHrh63ZtGAh
9j0BO+dR+SyHNtTWkLsiSquj+gXtprK5W5uyqVD2w0yarlLmUWWKbCQictAYErjQF/cDGXV9A2YL
whW1hQqxNaa/1fAxKRtQjVqNq6pyI/5oFCf8jG0aVONgvqkXioXwpgiyPZDvTVMpsu6ASBj844bx
EtFOnPcInjpCb3jgayLbY3ppe7T8LXjDfpIcgVokl59z+lRW9SvHDqdKWTqJKh25P9r9hY2ejLE6
bjJSd0fO1Oz9h8MExt1yk1BOXr4LBxAMjfj30wyrDCPODcJHGXMxOUcKgq3IuLJcQWDxyWsW9u0Y
1Vy1ulDn4cg+8v3IGfl3Rmh+p3d9KWPJYuXC8Md39Nv7s2dJm1DsLR3sXXy3YnzjrAsoPC+bifdq
V8z8d32bq5CIbcej+KGMg86AHStMEhX16Xh8grLMNIfTcZ9Kg6L0NqjD2q2+BCE4K5uMjbzP6QKv
EMhs380qrJa5Iaoxnkt21SkCkkTeITabf0J/qbQm/uhniy/KnfPxAtJnTkJQQjRv7f2yZJoOo2r9
zd9p+YZd0opxAlgslbf9YQh/HXkIMIdhN2E1ynGChOLR4w4MEYoFaoFUfL8DTho/SdYGicsJetj9
Czl/JVikMi1JL4xivP5zxJITOFvcLUtTqp47su8wE6dP7nhNUSMu2xfWiqO+ySCscfD0FQqBjjeW
cbpHx/Ztg43gJxUd1F3bHzSdgSEW6VmdO4yEuP5wdJQHdExNjdU3kWDQIRbZTUHWxg9FsLeuLpWc
M7VwSDE8yW2ZGxzc05VUeIL4aXZI86sk39+7Kq5QncCpMApGRO61qfh7tuJDR6yQMYeJj8SCtQal
bJVeWl/pCmpacWNQGDRgF1z+jseH0dbeCXvUbIpU7/EVLsNRof97+lPiAwXpzyQxchMUWhrvIHsi
5Bzdz2wEWGQOxeuh/I57hVmndJGWSFc1/OQn9fwdnGLwUEdBHiMWIbQv4+6tbSnMblpbEC3tHC6B
qZFCMPRvwO5hsnTmA3WWZ71+EtJC7RoB9NvAaXPvJtebQWDfAFv4DymlOooB0pHMthVaQqNecYxG
kx9VNE7BRHhQgtMo508rQFmBU781MgeQ6pFCL8V4YRfTMfzV8l8FrrXnS8BiwoJhB5PxsdJqchNZ
7jCezaWlvBTNXQaDGskJlqBmgWQhtmlI0AUMIt/rjwqkGWz+GxpZxbOqeqzN/UW1SrLtlPuXVUGa
11PUHx0Vl8EIXa4QYoOhcOgeufzlMx98nxlRR3G647PYEK1UW5t0063owAO/CEmZ7F13N53eZByd
kXTosGCtqs9iPOK4C8S1PGiM2kWO1rKaF9kA55qwBe5bIokPjpcAtN0R6Qc2E6Vtyq3/HYy5tFpC
wZWOHKShj2WtkSC+lmxp7CgKWX7GyxcV0F6T2I2V1e/YPN3rF+ovjvTrdrphB90FDWWNNnxeFegN
mtqYMKFYHVHZwkaQ0B4DjM5nodDQsZH0OepqPGoxXDgaVzmFLBrZ4wZan4Y+hKIMsu2/vlzqJ7f7
TEk8C527Od8AyEtknsfeY3r3kJgDEMQ14JLFrtfqbcBhRkc7O+4TIbthVxFoytcWVrOwASbhEimp
VDnngMkBjzGZ6CmzAgdVm+l6ol7ldQPUp0WEaQIoAOWfn2IOIE17hOLVF9cQcmAoHjxQjVclY21N
ca5r5eRtk5G0QJ2KmF/P9C5lJ3t4YHSoAjfW8nHzX83uQxwClipLPAyZbBMw6gquC55mv5c0jb7F
YLvnxkUETpqDMxUkl2sJVAXCidE7J0FhN8n7JCD2nMPU9Ti+3y9URp7en3yv75k1imlElLMk/4tW
mc9AoFKfje1bgp06Sg0a0Tqkjrf78pdNti4JEdGuf//ZToPopagCUMJFNznYIA0c3h6Ga3b/nvMP
Gp5V0X3ebDhee6b9qhuHmexGpPsVQxAHMMxGv/7CLfgjZsPeZUmztHWFwQ/UbP7HT8a4dBPnXEFh
wpF/iM1vAP9PeiM1RUeDELoUVGJ+HsHAo5bXL3i3VYZmQpjWQfdIlQry86/oPi3JAcHJ91Jyv6Tc
TeVC8Duf8k5APZQYuo1SBRGk0uXS+3fa2/zfVx72ZqeuLw1nl5JWPXo5gAPiBbzxb/qzlIAqQ/6F
pNxYFQP7a67GR99DEPTNENQCDliXMJQpZGM3dBseuX0/JsyrU0FlhOqfPrArQDee2BGS+FVx+N9F
965o1ityC22pP7HNPTNnSWRwPr4n1XsfWS1X0OvI/HYbDViKlJkjrlnDGIj4/3FO2kVqDcUw5bWp
d7Ii0rMZ5q/mcXCLoVQZfBvUmEfGWVoJGI8nlML4MzDgjmQiT7cJuF1QLvoDkDxhlxJRPh+uqBx7
2AgvMb1cVEXL1v15XS1ONLimGugaFQ3oHzeYUNGK+G+vw5IWjRhF1Rl0IAolgWyZYGrlqqduTsc9
XlYcx099Nlu8AXj0WnFjjWcFx4P57MxFXPh0emlJcUmH7A7e2js95oCmFkkMNlSxm2Je3cS1cKoy
IUxV5EAYXWT/azdARewYRfDEpcLejHNt5G0n8fMQ/jemCD4cTIRPh0N5ySfQ9yv1PBmMiPKfydLv
wxhdlwoClW7MXG9BYPIvOL/g8Zu2Tgs0fqRMlzMbL7qUZWo/zRn4Jp89wTieWZJOo4+fVNzAXBpj
qeOeNzSio7LC4xvETs/U728cdDoDKmTkuY5t40ogQ59XXgSKNrT6Yw2F1z7nsccbOjUSTKMDF7ZF
Xw04GhLSEE72oQecvwJ2SovMDzq03xh+LkSSzv7JaJgWBtarTHbCffyspU8vJVOe7Eh3U5HHUAlY
4pzk8VM6T7zd1WbqS9dr4WWxwiFBOtp44IrX4u7hm6j378t7jAOxRjBxBAw7/Xo+20r9fwfYlUdE
ap0ggV3h+arjijYk+pJ2rKqIkEbjhp4lx4UeAl5nhv9Tnb/Y+GmFJJ2ZvC8c/FIs3XBClSn6TTiE
xr8Dn3KNhbbsZGHDzqwgWTVlMj8vnsOLUAZ+d8ylho93FebvSglFxGsFWsDELSZpmxWDdxXi3DYS
lvrot/cpV7ifgSsWU+T8NiKUNVNz2rJhbONsEAKj/0/rVuk6eDG7AzAGL/jLtRu76rrYhtzJnoeZ
54V8doAKa5H0u/giltz+3+l7a6MQuZXs1jcRPc6kPJXixKS/y9Fx1G8WvS/m5tz6JfGDrrZ8wV4O
ezWJzZ8VYjjXVEYPt2VqZXfSEu9HnsjhLELCfAAncceIs1FAoFJ56NzuwIWLfgtaVzIOOVkYXKWt
eZI4LAGILoWqvHjAw79ifMSf+U7LgcLLcSramP7mQlnEFRPS7msolioBwLDD7cVR5FcbqgKsr6Nt
NexXbgco3ta4cbtlfDtauBu2hF0U4QPnGA0+WvmWXXTK0nV5V7kFEySe1VN7Op9m8L1wC+7n8ezP
g2ZdOgZoXkIKBOAc81PkMoGMmDcaJweySvl9jwv8+EHsl7pwD2vdnCTIFrz3aTYn2wpaMynBS0e3
rV73Wqa5aiyRZxdo7g7a5weVgH9WvNQ4jqQJOq9/dnVtqE3Z6+up6eep0kCmaRw8NrAncORVozJi
WE4i1wE5Fm0+OlCX2FahGty9pblrMU/TxFW53CyqGugv7nQ7o9MIoknbtmWaML7jxZLwM3CbE9Uy
L5YviDyZBijjU3pj9WKwY1Z7VvrOIAG+zJByrhXMXroEh3LWKD4gegSSRYXgs8u71yEV38S3qD34
7eQ2PEelQ5QglbI9NG/WFdfQD2V4p27VQDMTlPXVndPE0Lwaf+fcrcbtxrNM1g1MOGZi9yBfoL6N
A22Ovqk0Ap6KClPXeIOBMl+1QdFOBQEBtDkTb5uFUou0X/LqTjqN2EhIM75PZ1hNupwPD4fzVaPH
SieEjC2SuzARb46CHikqnNm8hE4P0M0ZhmlV7vcFBV0aQ2eaPM2169h3L1Pb7rDswlm5ZyP31E4K
7SmYYgWobB+OH5uR/GA1Jqee7DLBmW6l6VH5IXgHDPMrgxI5yjeIVHKd9nKY5239V5O5LKQlCnxm
FCGDpEDMjmytzoo2lsQ4hhK70MdX/iWmIm+HvXhWn0x2pyFU2XI3FTopp54eESgOH49WXhsjwFaV
lovMjwD4r3ff7IqsOFQ425TaCvFDiMLJ5GytSPl3TzrIx0AWXfRAzsTpbuJr5bVw0FegWJA5YNhB
QVLOFKmz0boHcKn6b5bqaZpUwOzbcCkFff+lXfMg+iVZAUGa+QuveSxtPjhe49z32Niw+izTNS5f
TkV3/Tf1UN6I7evHWYRn1wr2zub6drcKxbxl6+k3lX4VQGWCQQI0Mgefl938C6oP2qHJkDjNW2do
bMudT72zu1bUQ+hAertgJl13AgdybWp8t8h4b4EWR3r4LG8DoTx0etFDWtE8EhUaeh5Z7Bfy8jh2
wdcLkF8ZWapV7xb6dhfbrCIBu0m14Xu5Vhzgq9r3Q92nxfiYo6lTx9OdAo9uYcDAKAUHCgVZc/7Z
JhbClvQZAhw+TXDa//wCeGOJxKzZ14biPip1mU8Q5lakx8yNctHYcKqB/2vJ8Y4kjEpOr/2hA8YN
Ru1QAGRNmUrcol57MbA38TL6sGkJqbvUA8m4ppSa6QyqwRmq23KifdA54XXr1AZgZUkZHMiGZ7aJ
oCr8nfCmwtEiXFh9DCuDn809jBm5XIGHoxCurz3ypufd4N9kk5KixbU6LQjAQOdVcGE1lb6GXL8A
rP1VnoFJM5SWi7e1m0z0F4RShk0Y33P8o8e7DdJGvllCDfUgTAppIQoEjOoKcLPazHAVcqsLkn5u
ASxqH5kZVgulgq8ainYESMHJMNbSHFWbMT6rywqrkDcOi9q6oZhPqc17RVSfQV+rNeN6dqe+4Tlg
6MlxVQVplP+Nd+xTFPium2yRBAu1DaIaMnXQysssOYlrxQV7nQirRA7FmHrijAcDp/L1y3XzVZ9m
cfK8lnRMsbVcQPRbM0Rv2WmV6ruAxE82gbPlCs/TWFJnoHBxn3dsAPz8AbW2MH/T/0H6G0amNyh1
AsV0NAp0kN5QMgxh90DmRvtkA3huye7MbxIgDwVStNZgu0lhdISx3dbkgccS4WDUwjgJM8e2QkWR
9cy8tvh65zDW+u7AeKolqVCyvndCU9MNtw6Et8Dk+sVLcBPmkkk/E1jknGrgKNDvXDSwGZANgMiJ
enAUArrIQ72Y1ghv0p7PpSuStDQAFXyqrXjo1qfgsqDzeXQNNcUYVaLGj8bdZ/t0xuVU2NsfiplV
XTgPuRD0c7cGp8GI1cGcMd/oTsC/2vKOlt8KeiJ1QZ8lnsf4dcs6M6VmnoJGc+JbOXZKoQIH+2kn
ayS7T+7uWUL+Sg/DHBMq34gFbExFifwv1qAeLUbb4BPFPYa0+mPIajYUdh5CvaICx/XQqs3FcQZ6
zxZqYg/MChECcLvFonJvXYF8IYtD2EOXtZjJzAqEnqrQ7OP0yZNAOCpy9pD6P4lzI30Nx/fxeh2l
cxx4+xecRrD8pCWlQpPBRqOlzgk/emMF/8mzGSogil81JoQkqf4c8W/SvxRThBu7bL3crh8FL8ZN
XczL3qTU45+T/HTZnJtT3SO5O4j3VlvcaNYuTt9b1tZ7Wa2GOh+O6AbFUjvJZ+nNrnEyom0vEmsF
nnA6KvgNlgVVXhd5+/pQQF8HzNyWpxn83OlopwLMFB/vo2a3vTPGJgu8OHr40mwoKhkAgSZ6Fk8q
Lcc4Az5k8gLG3nQHydFjq/txZQk6IMq2RCPMbY6LC/TzfsNsLuDFXoPE+r1kXbKpXisumSzCr5qR
pM3nkpDgJIG08/9i9nWqtZIfgySD3b+fAuzkscYR+Nu4ai9vVoLEREoehce3AUardp8rcFHfo2Q/
a4ljUMCMMuwYiGBc90hx0W2nv9Kwkr6bEJcCPsWrtsJWwLynwyv93B0j9UxZgg14xFBkbF3HK5jE
B5OOTuNLxWI913tn06Rryil4dUBmixO0ya8ZSdbH44cIIHV04xUPE1x3EnJusBz6GUli9Oq33Cga
z9mRPJGtchpaN/p1OlPVs0wRK/CDkK40eFMNtZwZ/pyjuYcxvuy5iFmXeezeGNVRfP3I/ZnVwqIB
OFInIew9W0n7bnIBhJOd4g70vZGBMGSdiaWoNXYRvSPnf2jR7otQ10DpIGWyJVuY7Y1UpxB0gfkN
8x2Qe5vxl00iusC9bMQPZEZ3re7AftA5sI4QNJ+wxIMAaLle1KOXRfvwiQ+l/0cbmuztjmL2voN6
SexDy8skYbpFkQ/l0bqqMC+imvM8GmdfRHByHO17CD9fbiabtOxCqEjctdHsHhp8Z7GRQ+NOPsgf
pFzvP9gIEDWYrAS2rKOmsEXAwucipI/HIGb7vPUFwIdPsXkpDFO56pyh8HmdvQp+iQQjato+5KlD
3/gIEEo61Plja3NDc1Q1E3GQVyt6cibdmRjAMeK8qJGuDwfpFXikg1GIb70fILX+ZZWUA6X9dgvY
NucoH/ZAHV+VeNf2APITGf8iehGH9Frcmpo10H2ZdkyulaqamjjQpU4Bgfp0NM8iEw3CoLGnLkxd
kZ2R9ajFmvBQeBzbFNu7MFf5TVtqFhSM4eYrU6akiAwrNqa4aHFcf+qH2ghlfEZUgnzL8KOYcQAB
/DVwvi0utyBYw1D0X7kH97fmykw1MxdkGwvzIxraQgEjDZU9TYYCve0O9Ntv5mK71LTRX/FYl6/P
5Cu6JbuuRttVZ9Z3AayjeXScUwFZL30T0aFMy4xohAGnT4bIT5/DBNXDIaXnss10qYeo3/kUEI5S
Me/1GsLm2HBkP9GT7sLsvUvledDkb+hmKfcKUvj6B0LKZFDC5AoCTSULbBTfr6jqAXtr3BbUBsWj
SQDcWNLDA397HZRTtTb2N3lhFanI9nKxljXmbqvSZd8FVvttAvh6aaFcGkC/VKRNjk8M1R3tOUlP
k8jxrUSRhog4/0gsyafLi2pWqn9xOeMfPjbsqZIEdyMfRUM8GzH9IlPECP/4rv0DwLUzgyh38Ac3
3Jo8TyY30zO+Hk1elGgsVUcJcRwIFzBOMiDz1GJmBdk2YEETq0Kfykj+dyXMgSkr54kiH27o2+fU
sWzbpPcNcftbW809hKNp4V9XMRfUciUjB3WzHqXqncjYN+SWPi4dYJfYanMmAOXt7j+xEpJZmfjF
feB6ZWSUBs98BHxEIAtSP7uvNHqEYpct1EABlmZaSKs2PSxtgwf2o8hS4uXKIn5Q607z2omEjfJA
nh8KrU2ibTATBCrhugnQh2N/NLeKWNO0JPHsCynqlSpKZEZmhPGL7DFwHiOYbrXwLBfR1g3AmJoj
FlWjFy76IX2AiQD96TcktK5ancKh/q8q8uYucx1oZApll1RvVOyXqWqK57dRvkvB30Jb3TuI+L3t
ne5Jyybwx7oSR6Ozi1xwXOhsrLtJvHDSCteDaNaJ0CzfdL5hNBlQii7dSVRH9NgC1MwATu3/f4Q/
TNLJFGFP5KaknzrcN83hpeqiGVwsPAGqF4I1EFNSpzKyTSbLjc0DE+9uHGczenyEOzn25sVb3cCJ
rGPBT9VbrVGayzsSjYPgxylHn4PTrzlwsEAxkoW9CmqrSFsNX9xS2JBNsGTFDebGNT1eRN5709q6
lIGkq08UFAVAywNH+reDhJNu37Us9fsGu7A531KpRrcCkal366BYmlBn/fmLxdBdRaAWKp4tw2D9
/VlWFbt+005wAQUT70SyMRtXFhSZa0n8b1/XvGEuEXpqPr/EZFoFvrgwrEVaqLGXaTEjglSTG2wK
x2/3mo2PZwirldgIsJjDH8AMMYEnBF9gNUjzUyA+DQUrAhZ0Kd7domg4vihLVKSL6x7Cqqa1IHSa
iOsfI06aY0CnXkYDEW+0ETq4jF/MtUVTRuSFnGb3yADmGd+HqjaHqcwbHjJBn+ohvAfoJI8/v+4G
yVG88GFwfR5aCxXrnNe6/K7CYAj02JWZI0igbzwczkpcN/iZ7UmZ1wPE3Mu7R6qTQXpj9GYdKm6j
SF6/nRXty40wUyleTdsuY9SkK4DOZZyBDIesTIHyp9zg+GyNLNafeMl0diA4O/lsz2Lqh5FLlCzN
jICc5ORPm1CPAcR9b+OPKaDXBPcxzoRJ9latZuKhIddkpQS3sYgMj78wobVAKVbOzCVZ0MtT4iHs
RCfFwkbsgsJgA9P62DBcCzzIrxMCoNkb4X3syRRjbPxKfmoKDyH/3hFU1x//SxlkrYkKx6WJ5p5t
gYkP4PGSTwx7AtJo2ivQORs72go3Y1T7rpYV+iJ2Mb4f6Vuzaleqdh00iGT3bwi2G7zx45Psz3Iv
yMi4Sid4eklzMlCq9vYXZHznQMgxFLpzXBN9XlD71emVh4tu7x79Fho0uimLbL+6hFbr/u+Z4TtD
R3QDfcn6dCdcRuVxh2Aas+82zbx41KYhrMc0RNuYkmLSTiS9l5HsuwSwOHDoVgOZ2Vp2nhhWJ0u5
Koa65YK3IBSquNTnBSkfN8gIB4DeAWuQcJj7aboIONch1m1feNTq55Y2cGA4SBnB1X4KEFpGovP6
lOiD+sbiAgxZ6gBFtEiEJo6CnXDT0AT3o1RArJWdRL3+1QbuTGKntufYL4Ft/Ie73aKfrv9jYFrp
ZKZAvyvV9doH9knBO6twc1+5+EC4o+8FaS+tw1Pvf9OMIZ4/VVF4OjC4URkz6ESEjUewTi5qn7DB
LjzknuO21ciHMTG50T7EYUM6r8OEGHYk/rWQblVs09OUzkbS5nh0q9pI6QrWfCVGHs6f8K38xfrS
wkX0fPvDuN5YhiQ1BCJMqS1dxnCLlxV1oogdWcKtKcYQqqpKjSdNEe7WvUf8cvw7ikVw0eBB2X1v
MfGc9DzAVqOGYg9inEvsWZhORP+Cowa0G3BSKI4SQcHGfQFqGo+vXXyudTKBzR76YAJkMAWwMoX3
iJTSFzAUTPtxhceVcq54PwOCsWr0MG/TXAsDhYDIKswzayXHC73BMqb1UHCclmEx42viRtq7geyV
FL8dbQHL23ddsJsiiKadIhRzFEDc9C7/sKOoYMT5IYSyiHdHwHamOdTs+CYHUPDzFxoGpClVUgja
7XJ6yx23qo4l+mE6eXDp+wDhsErYAwv8EcA1RuSKQGqGbRU6JxjIlBWO2gy1RjtBMqKlMx21VIiZ
+isMWvxfqcw9bsSehDUAkU7xrumbmsixWu3Q4BxAzRhKDhNIoIrVeFJsvdGETH/n6NS5KtBDuaXx
yPjEdaiNveT/wyGMoSxUzltUdLvExY3DMJwcDi9O41RZwrGr2Yg3pjhOvHj44Y9WyQ7jMtN7AyA1
n9Wz9ixnPHzA0lQ1FCD+SNPGfEEC3P+W0f204qavwhKp8Y6orvWVbz7ET7aLgEs/DiQoMlYNiaDr
n7VaK7ItEn6kI06eUfj4EtjaFi7Ufs9A/SQ6E/TApQsznUEBwFxUvp4dgAP0RLm7nkNNTSKPjCZU
wPedLCDDFa4xuI4irqBmmjCOHdWMZopjQisWqKu4479nahx5DP997pItSX9nKV1NsCWRKIETVSU0
qJvgEkyXdU918CjuP1/ryHn0hSMr+jE3+Z2Thgq+hF1ZgnCujkHRjgqW5QmXxNodDrdWXNVkC1LT
mXCiHIb+6HIgN+BZ8dKInXMZAXqYg23CsYzA/eljpWsG/0UW3FcBuwpTpL/oTWrcbHj8Bgkx6Wwv
eGvP/jLUvTVhfk0rJeGe6aBLGzosNxQmtdHJj4bizK0ox130UMSR076MZm3mweUCkjeAg3kiZFtI
qRqddcPObCO2kWpRYLvQuAyUieAEDVOmNZDXIswHfI5dXYH4l/t8cNKfG98artg17jlj/9etxIFU
LK1r6Qou+HRG4h29YmKPWiSP1mCxs6Humx9DMtzsrPmnbWGLCyV7WkUn+sbZR7HZKLjuCLcTF8VD
d73aXNb6tprkTJ40R/dFRi4A8gdbmQnQANHZU3wlNXIbrcs+j5hq+FFVRugeSoa3OCw3OjpD7l0n
LrEVSLOvZ9i16QB4Qee9nw+GSmHCDAC0G9HKd5ZRmtnFSwPULTxQuspS3TZW7FBauqE9EkCz+d8K
eTKqvvXOVv8MkMKfmegcOEe16c/ZDhUzjAVNu4f8ZVSDfGg+ya/XRkpW6j1SfKl07GLHCEk7vHtj
zPaVC/htsH034YujgTybub6pbBODxc8kAGqnfdZOOEbiOnztpFtYaQXlreD3AYlfywA757YJAN4g
dQlhvUvP5Fnhqch2OAytzLQ0ODf9aqfrWuIuYjgJPjeqRSSvQv6TMBxAE1X7lsXRyaSRS7M/S+y/
//rdyPa9zBQhNx58weVm6wC9JRt92Vl4lLcPpSJs570bYkmF8jxl/DL0UbacoucU+syoH/7bjP/J
Hji4AcQvSfyNA9+Ib285mSd9lDZz1Bxu4KUegch4dItp+BcxTOFQEMwa40qIewp3+8q7Iee+/5/g
EAGnbgMQhKXKrsneJzkuqO6+ajJ8ivt/q9u1l8uAS8Y0v6mqjLXj5IilIcGPtDhj+3wZB56/NZbp
CWgfjEZt8v2RWCnMUQTEbcdQYFXT57jHHesnDGlRnAWZrgwdMZf/SVf3G7wHXlQQ7Xd3pMWUOzeH
3FWvSzcMczCJmh/YZZaJY9wK4hm+NlG6gpu8jc7aqi0GBvVjGwkGZbSLynh7kwYdjDq37ArqfBto
4RtrXAAtTyqcm7ejMIZIVNMOxGVo0LIl37WUj7MpfjkFNvvHWuJplvRVLUkFlfz6RX7R2HTS2iNy
5TSq12MTabL6x6xfxDuGwHeJ9UkB6KHRJfiSB30+ILXL4oDl2VoqF4weRT8ptEHVHRK+UGviT9mJ
VyOpn1Eu12vuxakzAavcoLJCvxfYGpNheWWeyCtrpeUC/2gfVsorpe3G1RTkzwy98/wzsvlO3aHs
px8BQRGjVPt/fy20LjTkz+KhuK6ayMdc+CHqIHufXoqEUdRW35LAPYPVgpDP1gz/eqURfFV9YUcB
oI62NACfaGMtMmE5nipfczKphq2rNoW83IrB6ScSr18TKKrob+GOtoPl6eQBl9ZOFMWXBw2mbMQg
FbYuaFhMq+eWYS4RzCT5815e70QUZem6aOig2wEm9TbNOfeGSA6heeGs3Z+94V7CSx0YuZqyU4Um
hZDP9raYeOO5i2Hx3oVJ/9cFDNWwClj8+opQrXfAH/7bBAQQvUCVp8+48LsCVHKqUpDJFQUeCfj+
2m24EU5yVm0MuOcx2TMC+ugb1CsdjcVj1yE8lJ3OU6/5hADelN9rLZXtJeYD1feYydhebnDTMpdS
0RjDclcYOBP1G1pNDQ4ZDXjD9fodMVcqf0eebs+T2Uht0FJxVJZVbkmxtF58YYR+lSBs206yK73L
SmEdvCLW/fIPMAR3ow5ZzRRVpuwujnUn4+KxWTQfiP2srxvl13RYGfS33LDgyk1z/iER71LWKK24
F9++YsWDOBayfkR1/xhpnEzWqaJY9N7LyUq5AZfzOfyj4+kWfUFyb5bgD+v7YJ/KJeU/58Ck/Rr7
568WYeXBlAQddu8Ux+zvSxVKy0ObyBvzCOh2TuAeVBGcRTWJXXiOlS9qMHuj7/L34ia3dVhsj9AB
0Q2WRMmUKwSjz/3lroKwoOSn7UgMn/fsK5xzPa40q8PuihcdxLkAezMkw6zgS2U/x1zfA04yGPIY
TpL2Fh6I/duZUddJnZYzuhdU7NtnR3RHFzmRyJ4VE3MbKQxqDAku/w4CqeITST8yCax5LW/pjEk0
T+H1SZq1gig6YyLIAG+3HxpWQJ5mpCbH3v13v8erwspxjpxqWqx4IWnngMnDqdPDC309CjsCR5r8
Kd6sfswqvxj6vVl0S5yLWd3Y7zcJw05QA+t0IDlp7n3ZkhN1WXih+ogaqA9/mdim4XoQCEgJRsX6
JcA+ADWb6G8fUIFcf880p8TITKlEnUGf24PVbFSvOlKBJAZyMRpV2ArOjjKbfeHD9Q9VHXT2aT2h
XLSdpOJF/xP9oatPDzb324Pc588IZpUcVW5HmK8oYfYhZYVrSDE/L613zgmeD3ysmnzKD/lj8k5N
o/LbiWH/7EELmejW73s2JO8ToHHhVfsztwgnGNQrZPWHFuWcLvRJD4aKBltADTUugzndyLB5mJqI
wWUnvzD7CTVPfuERg8fKqLaabtahICgVfWG26k7fbGv524H1tWrRDQqzWg/TJTXa6RrE15M71mcW
INs8HYmAN3fUZ2KrL4749GpgWLXZSXaxS5sDoY1HTDwyfJAaT911HgyQuiqeEQTenzxMEBVVRRu2
yH0B1VSuE6AxzEEWXcK88tD8JqZgWYntTYTT3QTNknGCXO36n1j5ZCoxkZP0+8wuL7SYSE+M3rDD
nijLlUiPr3DoEZHLrHpnBJ39IqM5xqvJMzhN2jIYx2xldwfpf4hOxThOfN5d/YjOU/g7h0H/iIpf
Tg4cmWmJL8Obh4fbN26sKOQuTi/fPgaO/TRcVw93RtCOMjc3HfcE6weR8FRozgRCF7LCN2f34//U
nfORZ4Ce/9XAmHYKE6DDVB9zQY0Kpci23Ac2zh0XLPCrFMVkaRpsJ4+uIaEL7CkSqItPQ+pT4r1X
VFL2iDdUxuSKpsiEzrYXEtVDpGU2VD3ejznbNySCei6hszjnYOurzPThfog2naAZV/7jClPM/HLx
a4b3mlAekQRVr8oiWKA8LYuFweCAbxI2bWTGBtcSeVJadSS/a+Z13PGMT4/m3M27D+pAPE8h1ZGI
uFslAB14N3rwiovFhVEFuCot7w/IhbjgYDvFUR1WItDIjngkyteKhIJindnT7XwEE10sfXJIFf6C
j87BvLOPATIaoZ6onPiL0BH3Jw7bEk1UqO8mGtx7Nado9H/t4FHSjSZKvnFXjWTcV2boz+ChEDk0
dznbV1+lWqxXRfOghrvqC/Uvj88FhtiQR41N+i/2NHXd/ltenCYLP3nQBG/G+UnR3toAajuW/Utu
arpSVBdXQG50tlfOzzr7iiqdS1HJ5sPYRWm4lQ8HvLswwhZg4CVWLx6CVUIxjJfhEEsPuvKqSuWe
OP6WsDiI6SsMzOWCUTs1mnVI1MkOmfbXUmAdnHopM7xRjG4Zi1LXqWJlV4+x+TS1+FWVO6DwaiOa
7VBaXNvLT7Qv/nFO+BjPcQoszja7kEXrdyPdm+UWWzywfcE1acHAua2tV2XTTewMVmkKbUue5lKs
9NkeSQq/SSaMAe2CrIHBQqSJxzc5BaziowtxOtXp6ey36f7pvxYt5b5kBTvWo/kOouySifUul6Zk
Cl95K9hFoR1XEUPZp9Zbrw9P8E52a9hJ1EhBRum/LlYX/nQoqnKdTmqGrac8M3pxCD9GCmT4ceoM
xlL5pP3jLdkujOSFEAmCrZV/CtbtZTKQA5fL/oSGbt2qAuXqXw8qnoMehC+5wvzzcj/yIe1T6TUq
6Gj2qowdKOvwoGQm3DB3mqEGRWFDy0lavYkRxo3YNOhOKHdnGosO3El87x46jq+q/D0tUj5rWYbO
QQlpKKfi2W4oPw+jNwgtL35+QVGUzlLhwe4FMyeUHZ1SJQwQMoj51LTbDDBZO+qwLukF99cczJzD
JndPx3JsEdmR/w5wbKoGXZe88KIG+DfYj5v+AyR3fkDT+DQbxUk1D9wjpTZv1FHXt/fsHyRCyTyG
ik5sPBmUWEaY69uuPMPqpv8kMsnS4P9uNkAZmAZLvNr99MAe5KKRXjbyoUmwS9Js1bz5f4SrHNTM
oZ26sURSo+FUINEh3jOhDrj4luJxhQLXBdVgcJ/vp/zMMM1fOEoNw/5Trk9TGHzolnM8nzcasQxi
v6C9UZtBxGjfpFJZAAb1TmsMBg6u51BL6atxWMT78I2II8ylhvJjngTxsMR6k865C2Eaa4LE068l
7eZYb13JukG3nb7hOFQc+QY9C5Ps6Tu6AoaoxKzZhbLjEv2o2a7UpNJpCuYtJCtZNCC4eSmvk1o8
fRqXpsMY6FxqUfaKQUM0J5iBmUZSy7Z3rvHOgRCz4f5HH8kgpzNiy50rYY3IeiuoM/NlAK1N/6/h
lcq7WsHmcXNveyQMUBuWKiWgEBQ0pF6aLztrbSeyz9DOalns4N+zypOxvaTfpFFoDNN4LUOfkCKj
vgcczyMx1gUJV5VEHcV+UjjpyBZosUHKrDJ2yT6mnklmyjlyC4GtpPfKgQ/R2IqBVME0gh2CJTxY
oEfAvErfrEEm8AYFKwAZbUqfaRgCGNFLSw+IQsR858Hpg+wzO+rmbFV30FzkR9QrSBO5yq22PfiG
aSJGgKOIQsTO8krzsQ2piXeNY2b5ltFigdXWUHtjoXlBgEP5Qm0KBG3OvTl9Kme3dXuSd6xaCrsr
vp91wvu1vmUaWkY9qn6vBG6m5IuFSFduU+5mllnpbAqPS1mV6r4H984AUN4NMHtyLHI8REwDteKD
cuidiuUOetxzy5ePXF96QunmHxPrpjtUXiV6Etrd6xaQhMeonEOjaJurqagePlxTcRh3/MXc9/0C
Bzmo/74ZDAQe8F1yvwFruqVCBeWgWtWsOjfyz0liCZMEANN7dgyVTFRD30wc/ZzMNqCWUEVBgpz4
qH2+7MIxz7beCY9MVaVY5SL9ldRxQc06gMl3+G744komQ9iTzLOeLAEps5T12wS6vRor52WQWYtW
FUIny3JxuOF+3jj4ESvjRXx8J9fmv9wWJDBo9YwBDvQjZbvi+9Wj7WgiWNLYaA6tlVfTUpgeKCuO
d+idFlpC/n/ubFAgIESyG43VtbLcLjv8r/952/wJPnb9rbGnfTRS9wavktCMkkuqs6XiFegd1Y8z
Qp2HZHmj2SLB1r/U9fVWmuC5Mzz94kTfnB4sNZVDQNUs/hR+lmwkcRbl4F7/dLWu5JzsxqqFqBcT
1NAK46BeVZoEIrfwjPm4SaxEU7IhoCWscAaU91IA4/zY7uWD8XMjeO58l5rjyTksRsTFBJBMEyhO
s1s0rY/o9R/P8ySwtPVKSkCTusDq5uKqxdR/6PFV1EjVKsey5T6colr7ITAJfQL2oeU3B0zx44RO
QpeUvcX4e1jizxV/jPoQbxi0BwmIkHcI4K1g9LuhzcOL8l4b2SfV1gE4tzvVS1NpbUbdr9JyF+B2
U/ONVBDkdxHzqxs44OS7RLutZ6awFZk6QFho6YNVnSCdvuS3lO+zm+dukCLNil/fie4OVuww5QJU
tS3SPKJFFxErPRn2SwaJWDSilosEUIIfiiOK/bKr4K23cZOlAhLX6iHNrishe6Kket4qWpYLWJYJ
391vvmdLE5PyZKcnhU61Qt3Mej1PLIWGB7yBfGFvvYEvHjNUALOHjdg4DvJnRJTtHgOMeKv7VCzf
mZXPVJYDT/qOCcVa4GX4q9RD5SiFsJD1NY13hE/B6amcrMer2n2WeQi1jflX7VC9iwY66ISMvE/D
7STT0ECAiBhsPVDr8OkQjZ3Eo/r3NcruTpGEQT3xZvt2KXX1aRNNKNla+3i4UDPKiBDGOlZAMw1g
MtXTFoWq4QUwbJsP751pH/yRtSPi4Rn9r6lNv5OCrjSvzKVKyQFFmlriaPwqVW4X5jweGOoiJyUR
yxDBL0GuFvp50jfMqzYEomY4TmN/lF3TRxEZbHnr/elv2n6b0chCh2qgsmCmaIxcESeMlL/4MAmu
mJKdE06MkZBtV5n1D6DTskUiUEAA8yEH3WFom+ypOMaHCTtWQ49OjNZ+RjySvewzR3unX41J0FAu
eOuIWwpfNisRRXCwR57E8stoAA7WJ4ur2g+wsqGnfKm1aedDysfDOE1buRGdPeL7KQGXBa2rDxgA
FjVYIm4z3eKZnabb9d/7nIdEtiDCWiTMjmKK91hoWrhXkn6VHV7Q/QTCcy1uQPQVrJuFF4MOT0NL
uNGbbhPwtshHb0iZpXhVHoUIf77S8pbSGdRHJQX50xnXvzFT50V55r7wxEreOmec576pGePbUrSP
u2lZjwOtMmRMejPzhERnDvKXb4vK0Bo3sGkTB37aAvN2atHtRgRkMguYmuNmMNFq+rFar/LjWg7y
l1GgqBafg9uTJuBRMhHC4WUlF4O7LUlOBneyl2nwARgRpR+3wEtdyus8K6PW05TiCqmIcJtUCr5h
NXAqXh03Gr85OIojjKjPsultX7RSC44HH3s4iGoWYq4bff8gLgb0E0b/KRhox7mNmFKr+TsQRkhh
q8/iD1N+Lq1ogEeqGMpEffsnbxGAJS9K2NC056YdJJ0DqBZUPCi3jKUPe90bteE9MljuBUcs70bb
zbxqzcf3eLKZqJaVtUuGe8QHrDwxCN8mWN3dgXMxd9KdeVAqsmcCi8+Stldk6fCuaBhyBC2xvJ3A
a0sDHDnSpT/HhKbmVgurZqbIkhL5M578dYNvcI/4YFt/lU5v2W9+blWWsgdqZJ2CMZWRjqRSRmYF
CPZz3x8TzLLrX0tu/fKIoR8whWnbbkSEYtZ+4GF5cuIhmHnuaNWByIzHEXaKXLstWSjvocYk5Yrv
BflTN39OLOZHj+hoJIUtStp57GXYUuBaOSFpKS6t75/R8ZamOro/QxwyucJY/AiA6t6wyj/OC4s6
o9HoNs+CX88WsEin+E/WcLAvt1UfrNrLT+GBtDQhCXlVHDe30+jkKyLSpPr7tYl4RR61qIUNMP+Z
C/HgGUgkLy7eFCmjW1EufHTJ1BWlZhFqYXGozpKe6YX7DfDxRz3BPluQNvD4YZtOitRKfrTH0B9V
0oduJ0nZcMl+gJ6C/tDPnXHes6Vcsl0V/taStrQMrye7B1+OUrdx5ogW/VwUL93PpCSNLbmz/mcQ
BLWJXoz0YJ/Nb1Hr1VAz1Guer3miUJ95d/ee2sGtfLtF3CIzKbZjph1Tta32dcS/y5OLVA6myg8P
AqLIuGCCDRPWYo5En2+0PryswTrmyHUWPsrGr2EgsJXMTxgH5YkZlL0sEBLh6CO+x0cQ2r0ClqMe
RGIzR0QXT/iMfMGuTjoyX8h/hmZIQDq8YgP4Nsr2qPGvXMayZ6o5DeZuvhdAWvQtIOTV7bqcYeEA
Uh/iongGzuBujoI38Haw83fekIC7IjCoETkcmyfthzH6BWrJPfbfhEhnSlFBewl120OfGzYh8RKu
pnKB9RtMf6C5kfW/8DbkNFKc5FrbNi2cuwGxFgL8oBkjXW+/mcOim8Cj56ffTHvPeDhAFxz0clTg
AEoGhCvlbWqswhms+jnFUggwA9VS159yzU0v49dXlE+kNcmeTf5mzpJ47/7yqShrWP4ptkDP9k3O
7tF57TPT9Y0gb8SAiRaN/9PWiPiOIuBJXesTkR17U7mYt0e2/2F1V64ugEfFKt5kQlsZkPja7LE5
fKEBf+pO+qL4ImafkPjZPPBWcFDk0YEQeNMAh+T+xVLoZ5HCTa988+CAtE7ylwOoydEjm9tWAyp5
MLj6XmHBc2Yeq/LlvVapv5lsiY3YH1gYltocacOiBQ0xycm4wqalcq11ULnv71gfHc7JF8h6XRwm
P7iP55pBotvw80ghOJ8bNKx+tlYZD/1+VwCulQ1FVGUha7pzqLF/nVkOa4m98xASZHBVVFEJDR2d
78PmuwKfAJCBVxvwpeG3fWpFMDx51xchty6nJNM8L0aihGvivSlil6I9SrgkpcyBVe21JY2VZw3w
o5rkbzCazQHPgNe7cvLVyBSW82+UopIHIxAmbJ+wThA5dehTgqbLUmNfjwRDLTcMd2/8DPVILNL9
ArirDq/IctL0FjOYvBVFataLdulJdEao+YQpjsCII458JNPMz9hTVKKKsLZTwaLZ0mS2ZA/hMyjm
8cxLjGGD314iDBRdxGv/fuettEdGtqaP5NCH70DdkV+aHxs7Je6yebc+lAb7IUx/xW5QztXQusTe
YnXxJLjfE1SxoOHAtdhjQxVjBaLMVmhE2YZjKR34BWnHnayLG39reIpzsH36Jhfgajg8DvBEjs8q
SdO6Gf9crHtqBzPs56cWPwOWnZXMkswMIorTWud9fZteQnCkN1D4/3CSTU0xywEB6dWXoWySpa8e
CU+/Mz72i4kimOoffIpM2+7rcqYOaTiqC8WB72ga/l+a/2KcdMD7fi2xeMIZmn/hITcaIt4lJsA/
0XVMeFo8+qR6CFPyTsei0tL5knSyBl2ujZs8odGzLwiMf63Sa0DqOVv1RhKFK5Zjpws8Ka5wRLBP
KuV+M1iTf1bLpsBDf6bO+2ZlpIpgxpSDChUeTigfXYaDa323bBTjdqxGTnoC5J2ssOsREu4lZ1x5
m1Ve+0nEiVs+8KfyfiM2SoLbo/cmW+RowmCXVY9nNyWuZ6L7HhXtpTLORC7Uq4olfeXvJ8n29Fzz
rRtrzOx1Ra1swrTLGyzmYWQLLO01NqkK61Knw7gMDsB/0L0ta9inLSxb5fUvWxPhKN5JxF6bEJEk
qpRU/Qh7ve60f4mfBBBr8IJiNwe0FUouu7KR4/EA4R5/1NCjwdKUBLv3JOohhCO69tDFptIx8wuv
9/g8RX1gmfAylKTf9YDarhkKEuhFpnR3suKpR2sN9GJXl3cntUguT/g65kTjFhQmdlZNCPgF0cAv
A/XETxf+a+YQH+ygIM9qOBf06RN7NfxxWz1g1AZ7HLVPtDRoNF7UsFPhbLeWWershdOAg4mwlYgH
XnUl+VGmr8ghjsNyRyJtIktt/7jnRGMBTLyBLORksXC3IYa69V9MlniPPQ/spLiGC/aiHJ/jmI2z
XuN0CpsApKbqpADqmV5rwfrL9p3ogUJheSiWEyM9kA9DO8ymD+q6lDfTPHRgWk+bS16Eg0KfHBqW
jf2hUqL8GEzqB0RJxhEkq1aUVUa9g00XNDoi/+V5qU8p+aKmy1g2tE1RTy274FeWOiKtfjXqsY+v
HsINwQNkxGnEhEz4zwkJ4IDdbm6WdM7X/TOnsfani6jdk/BrHNAVHay6Q5r2X9mGlKxU6I+cYeYF
DuVz50vZ6YoyszZrfys62WFF2f8ol8Ql59W7bjSwH36fby5/JI50fs9Gl5QS1imYpNOj8CWKyngS
12QH1LPmZadfWTDfMTwmY228Q/ikXHcvz1LFwYJaf6k111SoN8fzbO44XgRUnz4BentB0syIRPLE
hwgXQq7PzhVboeZuq5/Ph00v5gL5OvmGtioQ63ZC5sjNeIelwEXDcpawWSesWdDjtqZhCYQgKkFf
GOL30+Bg6GLiGkNGRAAHIOH+hdf3QNhBNb0N0354HTq9SbsL5MqNonU9icXlujI4s5QJF9xSIASO
6MndDcO59JanvMkZ+7Qelk8aTkeNIGN0mJWM7rkHGaeksnN35OFFiP6F5s98kujUPu4MX1NLMQ6B
BOHerUEBwC4rIB5kLBcFK6Z0I9DyI1WjB3IHZTp0N4ZZ4kZyx2WlXLUQqrcciXDvfzGseF3Xx/oW
QGDNzgv5mnc1UTj4ufFlAyUBpIBURM4XwKS0xbD4DxB/LTf37T8iHPgMOIC7BrYJeyx/j/kaAP9Q
JcNQlhzIo6NmTrm5GrDqDAPKiAAVMWA9NIb3TqUVQf/9+XQ8LF6fKl6paw/hYzeU6OYpdL43kK83
4iCcmHDeCFtJLOomTJ3gjpJCbOGxMCjnkfNvRt8/7VOuGX5EDctraBnRfJfqhEb/sGjwgoqajAYX
6TqMNcctVNRr8gJFawWjPCHKElpMA/M0WdCIOYfkig7rIUG7jJQXHLwVTd38NnaJ2JPqD/mNhTSX
PhAkY02wyYXLCxTQFftlkWWIywCBu2lBHMpRcx95RpDah2xdApEpO29b81Byu7PDZIqYfHXd4O1J
toT3ELat2Q2M0ENfpy/9XMjRqgfBG3dOXM1X/tUU/ASYew9ccIEOzu4mC1IFA8CSXpWT7/O0e75r
K3zmYf7Cl/0Dk9lCbhMCPaYaQW1vfgvgZt+FpasNRJJs/7F+XY2m3Ddblx8U0of6b57TrGWJ4NRm
zkFNX407xftJuBYq5TX/rJDd3E6+djgRUOApaEo1YSngobjtRzNy7SWIzzimiXk7/Qivj0/m7VTT
mEhLgum6OeDLZPTaIaucHL2xD3L58IrAbJSVKRRQg89rTuilNXkDr53MjQ7gMVWQwrSU4Kr5cYQR
D96SgbCZJu1FDvGR+dERWt4FeZKA2WIKL7xFbLKiVXMx9EMSidDx932ArbxMU4PuNz9FDqj1b/TV
dBbkws5aUSxht2MJXgFHwCTDCe4nHo/+Mc3auPaqNnYhM7tkQE4G1eJwEggKnSD+5nQeAAInDdku
6m8mo0he9AT8zgZuK/Y5EkvdzSHsTyWM4B7TWYUf0bM01+7PSDncVs/J0AbJ5GJWqNfv8UnU72hE
LYwRjUy3KvtbUEh/lwHfMEatjikaofhHV/95tHotAGt0z4rMz1zlY3vNqM5mqmR0I2+WNCW9QYuT
H2gID5WpPnD8VMED6KnnxUe5fw/ujpenUT7p3CHLd3cV/X/mgzasy9lBEVf4/x8aqNTVS6yPpMfQ
Kx3maXjqhIR3MfVyKgDau+Rlk0Y9kAXFEjfqcEqWst+rN0u62HaUhfC6kvx+M6LGatcKsQR+6s9u
uxfeZbBpm4vzgeNpYr2rRViPXCCh9GsPW65LI7JrDnsPubWnodn7YUHtoVEnOfhKPvLq1utC8zXb
XqGS+YdmtpJx5Cn+NCyw4aCAOjMgFafqItUScBKQl7GgUq8usWF6qGayAClUo71eGbkEQLDsQ17O
2gBJsuzESgkkio0LgBYU5vwaU8O18BppxRkxDrwFtZRMB/cF/zURkYViDgqjk/+Q3HppXqkmzAGQ
z0QQYJsI4McHp3x+IIt/Et4f9RAbJC89ldjK4m0+mAgsR9TGA1kNQkl5xSCKg91gLxYT4ds/RQPN
pFMdN4LaTiwfjuDmqzOcDcZkh1x6ReWFm+NqNE6/Rz0BlL1EQjNq30f+5m6GFlBo5ecWBaVgd+RF
O01gntej6BW8jgAS4cpArTFJ+CimuuAdd4U55FWoGQzHqXSQhSMio6AiXYA/6ospGHQjLLCQVXPB
6Ma6fZVmcXYpF+JDJaqui2iy5p9pbYNRpYcMrScDqOL2G+hmGZlTaOmeEen4RjfOLqNaKPz+Fis/
w9wnOmZe1kjKYmf/RJFkFwYMKa0xMhLr2kSL/VGHBbwXlOH8xzYiSHXTK9yoq8DXWwMjZrbinMia
b6EgU5VXseRC8X8TXHn6PFxeNJ4gBCctGQmDrPXnf7Du5xB4XyxNsJAezimwtwg1Jw/Ug/6XnGe9
LwhCmh2KvJFsiY+aYMn3ovr4ZbhSGd19nfSFn4t2vnBxKzXUlQW7prGS5KrKOor1bNmrzjpnXCJ6
6wRSK6eEffNcYrDb688/ThtMJyEZvbysSmB9GEs/O286Qn0eb+vR1y+uLdvFjpIDLhJBPinIvNEw
+/Biy8FC8NVgn8dwLX0+Jo98sgss5vYqVoiTdlsKExMY60F7dSJTOYTAfcBG75Mo0UwF1Gsy8tac
f0aVZ+a1qLscYYI8NPh4MHrZhUoVgN0ss7+C62OgaRIgMxBuWx77KUcWPtiDMASS5zmm7JHUyQwb
QkiEv137rT5gN4Z6lUeYmsyUviFwaqSXmeMleKnvciPZsOswIOQuaUUTwle+s0pRVd2h8eHXBB9l
fLAgGMitj4P2OFiT/ifdUr0aICdmJAKYWbYPKKJD/R88gGYhZj1RB6K10Huf6D683oudZp87P6Od
LiGd13TWJvoZayh1owyF7+uSqMpVvNtFeR1GNKWPirNXIfmthli6OmhEI/LlKxOnmWv5iwsclTPL
Drdt3q2BvtLWja74kiA98KMDa9bT6teisvUMAxszqSJvenucdzhslHBqqHKEKLr5qcwi8Ovt9OTP
CjZXD4cF03OIt083GFBxvz5+dH3bbgKlyOuWYY8CkqR/ZPZ55X13AeN1dkVmUX4tS9ivKnjmw/BK
LbOHCLTksN1DrSsAWGgNNiuM2x7urEa3Ov0NnGHwRRx7SxnulxL/rgPopReC2QBWoFt/VWobreQs
j0QaeSuAFuVWyHQmc2UZilx7o6uQ5qiEKvFCPYPjZSgY3453Hp/i0ttb/BWdG75tXvaMRRUEwFhV
LlrU7lHJYCkT8cZDku57no9/GIdpgMw56QDAQf/rWn84mqclAxiUM7/PVE/xhTrgwOxadjaeggPJ
xCyj2X8zdv4K1yHWLS4YIeRmef6tKN5+5LEWAEDzpL/UQrvMAAkF/OBbG8+hLS9oFATqN+eKuyGn
le5IvBDkkoh1pFNFqrO37MI1zGPn1aSEwlyM1O4NfHAWKV0DYKTS/PHM583iy7NEj9Nkxxs2s6j5
EqMulGX4dc6EeaC6T4EelBqbEVGinu17wVLySnCbPyV64a+AfnFlQKnEq7RUQ2dUc32+60V+QpmI
bh4KSYgv065BJeqJLz3+67/gul0B/y0ymcaod4VmCxGmr9m/V5YOFe15yrPty3MaapX3oYymp/MK
0AvvMlvPErWtYQIYAn0Px2/yOnDhvok7knJTjKfqneyYA/TkV9wY412sRCCah3e5yi9jr6t7IEyv
wGr8plm/pDAfu9HEPF37wNYul/VN2tOw+FYIUz+Am/nyFXgK014QmyrRsSVzhXoVLUGYQ6Z18r+D
Ty3XP1RtaR4mkN/U+xR8MD67w2H4RgiMnFTlq5iELG2Pm7WfH3TWB39soYZAs1RU8rBLYaMkYU8X
kjqoPFhr3yKeaNuXDaSemm5ClltTdrbA4Eom5j9gvfkN+1WFfrGAmR5Np7t6lL+Ta4w3DDOBDmec
wwIWmU7Gv2WkpIYZdcOH4cJx7pQ9JQovuLTLXr+S9xHtTM2wSU/HZXooTaxqrKqa+nK/yJTirm26
fW9QSTZIqt01Voiurvs0MoVwJif92kkEgm0X3lRFrG2FmwFBRbYKEf66WK9y5Bxh8ZpknJ1Q8o8D
5Oq/kIMv0X170aVHudcPq7a783BbOB5O9Nyb+WYcGk0uZwGXC5fEheH46cjqLJqrkJYcTLjsJm6T
JVdfIp3YGbIRLBUhQxM253H7Zc6BQUAkUas61LHOSN7SBpo/l1Nrpvgi0vD8FLdniZ4/KP+gFhkY
Q/6O+ILzTl/hVo0n8Sh2GeRUvzcJ8B5inDz6xWDWw0TXZJwf08BcFfmW/56aXlddG8E9WVEiwmIW
RVQL/88LnUpBfB8ZYdlVxPs6jzIOjxNTsTAg+RV1MTkPEh6KPyI3wfoee9R4IQsShP7O1kC87eqT
Mial4EcEeVB8gfJjvCnubMDqL7fZwpR6OwN+Z13tBs5HkXO9nrUnqnNUgqH7V+6BsAPS1qY8LulR
tCt0ycxDrcVmOdYBaX0ngrul6fl7znOA3mDeotwmtEXmCl9fOnrCAiYgmvRITNkE7tFrJ1X54Vwu
FHP8+H25GvDPq0Xma8SYlDimN6aMc9CQFCQpw3YjFB3H9SxmbKgm94C4CKcKsryRJNjQE9krmdN0
1+C9UsLmPCtwhojj/asdQQyDj6iiyE4UWlbFUbFYVbD1WgMJ3TTCBbFR6uIY76+zQGDRN/eBAgqf
8Xye8UhY4U9Ki+WyUQaC1VGi7KVW3bOG4VPvII3B4DyBrGSzC0qa20rHp8Uk9OtjHlwqjkbJuKWe
TrQ5/KIvS/M26Lxca/D1Twn1yG/kmYXx0WS+Us62WFvAxJgARZeOFK9JkfVRkkZbwPRjV3M8oyu5
9J1Kjp/ZxqJzIuPp0H5aktJHvun95h7f2h131kIuzGQ5iu1NHrndp++u3eQRXs+mvEFiFFai/HKk
rqH44Kqsv71ZH5KGNb3I5KRe1fDTTGtl0nOWD+nKpaLlHncEpu1g+UJtBfGXw1ZsUoyftHWxdAAt
U3IpHxoMpIz3gjky1l8FgGG1MsLwNIW7FBfj6GxzQGqdXfj5JdocvUQu/em8yWcNGCoMTwyJ3sEP
SbWBgdnpicRZJknpUps7QYErZwdZWnc2Uja9P8nzHGrGHteOy2z0/F8rnw+z/7EixjUICXYlDdq2
TZta1X5d+TBT0NzAAsCvRegjttXv2nDInWaGg30uZjqHACj2TRrc/6zwhu7T6QbOH9Bz51/Wu40X
ScFwDKy6vEf4pPijmYhCn8NqWfeObTbxd5iRico82Vb61lfPCb+GVQpAIAjwLbnrIA3tvHal2det
o6oTxt8tujhYK0uIjMVgyvzxs4Fttm8ZHC2Dbvdgi6qn9I8WAKNANAEF/oAkh3tzRoxD1A/EeDl4
ZSRwSKUk/HaHU0uWhYWLZmqkaHuE7f1t9ovxl/m3QcjeBcIJRKmB01UzRExFK7KrBqR8gY9VULd7
02NMgshg44C51Xme2fQwODz94Ot1ZiUjAQiTIHFfQeHC6Nrr+2VnEA3j7QrxJUNhVXG3prZB8K4U
ikbIu6To2axR7EudNnj30hgi/UKbR9DP7IrBRmeJbGM84CITsDYE51tqf0VbnvMgnSyW25P+haVr
xEUkt8dv2TURC0YTpvOgCJ7t8pbkm15/Y1wElJscycNrqcuibAPoecJq4NibTz7XuAMatSnzDpw9
/dNIqcBhGDPgHPWdaWKr6kFuv037pz1GtmxOgpIhtUVaf/uZWad//AFtG6l6TUsWMl5uL6E2sicb
yTtwd/v49RaNGuo0JcJCdhjNs2nWFOQmPq/ZD2qxGpwOQpr/T+W6ZIYYU4477n2vSPVM1ya7Uvxm
iYXVDwYrYdQxaCcoKd2vzmTTPRBDUmejbu+CMBHZj7J+bEkzj0RukW1CLuyM1jFuSVzvosSk+NMK
nunLlYcXxTPzBblhwM4ujontzYLQxWeqdyXA4ZcRO93KzonTRB0fsKXC6K17QfaCoLZgDc1m8t2B
bDctI35DFZ+AWnrxtD1I9JFd41J8L2OydfpDIdF+RW6cGISzzAnnDihiVyxAeqM2xuI17SDZUVTn
K6xIycXCz0pmBRCuo5MKEezXlolyHU4R048VK1qIp1yMkVecBknNjjTDJZEFDzg9WmX20KDLGcDI
ibAfreEvT75XdNm2RXRTF8VUr/7qfblP39cB9WbNXI1zhQ/CIJixhNMnI9HtQhuu9g1QQp1zgXVG
o/hOh6zxIsUWn+xXUMdXmSmEhds92xzc4US5q9hhCJOVhbKBFG9YY78vCk6yTZGafTdwZExQMNzT
YTiHwrvTXGGdYSPgEsK2Xf2ZNqNUcuALaqlqPH0AYx8h9RGkDSsVPdqsG10BF0geB1qKkBss6mH6
FYzW1QYZ/Qo6Dyj8WJUW9qdXfBjGorOzwL6rGAqNU/yAqcqp3aXPyq6cOaMNBKrxXUxhVIRL3vbw
Av5k9PJFjSz/u/bZejOavZ0oy+1oc1GaKm53OJL2DwvdL32mLOVxtWT4d8zajVNmO6QlRGUoAUM4
ySQVZXpA0kbe0BQnTZh9e7cM4PyNiK9f1xNqUpZJ+ZP3DmPxpzsUAMCTlXhCyY/PWaJvoh3TR9vp
zB88munylhQ35Tzf5mny+BnKLvNYYdeiGI8nu/8vsJ6AgX/xrJRI1XO9dLq8sWe64UMJW+j6G2EN
qiAXKbOT/BD+U+RaLc/U6hANdribmp/TkYEjjmFVgbHwMJl73vqpVJRXi7il7xGWFVFk0Y4FJkxa
1ATqJ5beHxxm2p6K+8mQ3tIm1YYz8RCmKF1OU44JXmh2dEx2P5ZgDAnig6HZX59bzzTqBoy1ibwy
Q7yPQjBV0irN0GG00Gm/g18fNj8qq6bdr9vm/0HiUO4CP5bz9I17US/r/WJy1UVhJ0TnUmvZbauW
FIkneqsw8DueWyJRk2kWmkFwD+7jsI/refF9nOA8J/91K7oh1Ez5ZDjg8XFoo1GckIoQTpwiOYWI
k9xuEA//qZZ8lY+IP7T4Yqn8UjZB1FpYtWzHacVvbFHLgu7tvYktiHkwaLEF/khaPvCZom3Xf57S
k2YhyKTOFG4WtT8mkZx0W3LU71EPbQmewvL2ZSqw7RPmxWbskla24+atLfLSXEj7htJDZI4EFgCn
T2fLRmMvTLykCqtBajLLUcf0nm1vH/A05rqC2WXTRiEuKN671ZtoG6vJMsZBEU+5Ko9EN/yOY5Jf
JFuDobGX6uWEyhb277KxG/jBaB94AcL4aSDEIWytN3mQOs7QpMOMbBNEvNzmZktgb7PfXQ/GFAMv
y63RxGlD88iaK5RWiDUYIHBtCDSxp+INJyfRn4MDMVKTqDLMrpG+rFm+vpf2wTITCafGRQQHuWZd
tLklKEUMSm8+GYPAfynh9qk6EGU9ufJgokg7Xe/aQh2W3HyBGWfpdylsvfUw0dA7xVKgbS3uAWcV
osN0HIMgi0XDxsNTxW9fAFRwgOO3x0Eke596u5FVwVvYVw5Zv1+Nggdo5w7t6LDpXIcJ3SqpvkLe
Vxlp844I3AUuBCpOdcV4qG8H4IQU0gGjWgeAxxR4ELoY+I6yo3bzf9ofjCi/ejR4g+deMSBFFcPc
cTXWI7suATFkPiW3LT6crpqZKmSq6UCY2gaNWbMoYgGERgqN5b9+JIiC71B5/pVD/lPXxXVuG+Yg
PlZVXmk0gi67vNaFWqlXMhfrunqv6oA7GFoLzSN5ZaPL6kr/anEkzxrM9UJT1RsmO+XF9BAtq2RL
mQiszK/xKfG0IlxzeWsbr/yI02Ygctw8E+n3c8mZNb76xq1UgPvgub24+o7SvQjb2kHNkwPhSgVu
Ugixl935WwJRgZIByivTuIpVumslupf0CWHy9gsNA96UuSmT/Oxdt8m8aox+lilOJJ7ZmedhY5Bm
acoUwzhEseWCdzjmgbqgQJRjYE/+K//NuFFl/03LxO+HPTR/0RXsldRX1KagaAEDR+cS6z2E1mqW
idFQLRLpKimbGR0hAeYgJNw49eKB1HzqPn+utGG6NNeB7lo4gjoyt8JTk6hHzmcRL7Fnwxyk6Nu3
ICGfCi7oq5IM/g3arjXJ8KRHwy2AgBtCl1z5igY22izLrnSGY7XD+tAgbsMwEsAyAG0gp3ZiRFgs
IFSkPLAeXaO/hTAU9AMH5vPFAdFdGiMgWiMQHKd2f60yuEIndkYBbRuBcbKnafmVSkUrkDAPWOC7
a+tjG9fn0uRqWtcndBXIsVl5oACx26bFBWGGdNMBvJHrO55R2oYJkWNk8pZ3LNj2r25+7L0s7ohF
XVc8BwhmzhQ3WG/O/+mTaNUxoQHcyaGJLMEajGcSjW8RM8tiU5QwPkvAl2xpthtZzLWrmJqNS+ut
ZuSg6pjP8dY+cMw8v5cI93ssnxlWypr/5htqeFojccSGdeKMcj22uRJC7X+xSwA7QRaGy6BT7pNQ
lg7hCP+jW1Sy1aWr4M4/ZfnKidBsER3NfblZkcye2HZuv2VHPnWZfISY0qoXIASUmuyXBpk3zmjv
56tU1CardtUx+TbG7uK0n/e8AimUd5vqeMcaJ7hhPvuZTuYu1EL4Wi/3K+72OxFfnGKylQa/NKFr
9MXZTecBHVJwXc1lBOwzdH9kAzqpzHmyUvVfDJgIheCHfFmZm7rlo8nuli6t1f4I0+T4jsb0ys78
AMW75afyJ2Sf937NZQ7xs2pLT+9MigEmu6xZ40W63qV8emGQ1d2ZwciEDHs0/Hj1zRmb68IF6BHW
nD9Prn15EaA93lMHPLGYPUMXi+TUjv7uMrJksv53UMQ12aiPpCVZ8d/A8md7J8/HURowy+Kfa7lE
thc7mxjP9cMpPc4HVIUeEQI8Hc6vVYot0DYte12CiThaDk0Ksh/Op991in6iLO5XDT0x6Drx6YP4
fO9yoJtbBOljHwE20COU/Ooot9fmdGEgNCEE/+s7ql3p59rz0KBbJsFHmXuV/78zn4Xm9ptAhdU4
RN9lWfAUwslRxwq6rMPMOsJJqeGoXRTgQdSYr8IMZuoL25ExyqdHS588a7mha7pT7MSbabjCI/lC
94VKjFOScBT9UNwbuMWpjpewOfuo1XksLYmLziN9bpkWa+QmFV3eCERxVzDXzKXgkikEfIhoOPDW
um2D/bCPFOhDy8p0oWkWdGWOWY0OF8wnC4Nq3Bgz7iRJrL4aetArvoqqYniwHDwtmeyKjI52LGEF
rBK2Zm+1LHVQX3a4r5DvKnIsN5AyP6vdDfEsLZz7Q+QubeKM+mRrEdTcYZYgikwMwg2ObUfLmrQX
rRHddPYbBTr34bKdj4JNVZbI89ifJ1abOoe2VMRVJ6h4Hs5nYBE2E9NQNfCxGYjlt8Fz8WW9kpyK
F8CKmVyLpjutoLRPhMJTV5tuo7YxDJ0QURvLkq3F1IjO+r8y+T38utcALUjENJsAOsXLf5xJpKHU
cp3Ea0nAf1giCD/F0wR2b/KJqQtHdpSN7YIE8NAtHwyDatqpaFkjvFvTpfP1R/0WZslbQRu6pksn
LnjHEPfgNsc7xmPd7xMvDL4i+fDENr4yxq5v9lB5q/KvGX4Q8WQEOYX67uAwqlPn974YPpvkVX78
7sC/8Z7yt/I2buRScKE9qJk9OQ9OSRcYftc53xAjsMid5QyUybUmBEtddphCU1br1dBAHL4BVCdb
PoAi6idTDIi3FN09bcIzAMiDGLnobvnHVNTCOBDh5xkCxSgMyEhv7nAkE4SFuGueh8GcIShaGs+M
m65Hqv5f1Rdh3PrUeBSRdr3O4C8qmU+WR9ECRQ4ATPs7DYg8YoqFJb7hylhB1C9JHNtduwOlmm1s
2aJJozeOGHSECL+mdddQ/rDdg+7JBAZrY6i6uhhTgTJd8BBUaVFlQsM0IoONUkh2zDne1lUA+NzV
3JlFAZ/pne6pRqje1Tn2P9XWFzqT5iTyXYWD67LWgjHBFru+ZRjFVB1SqpQlpu6bUNXeXDNxE8iJ
7dbcqKp1ENjmTM6R2EW7dO9A+blaaOk0OlxntOYubR4l+bbK++hBo3FrX9JBQO9TxrKyl/Zo2YJb
8C5RFVFlz57K+GZQLS0K8Pm0mQa3X/tkP3Jc3G32xUw3ElOCQE07o9XAHTszD+h0XjpwkKgYDEmJ
GAw/LbQdZAMt25PKBVauWBksv0fYPwSS4Dai5L7A6ANTzRWqQb9yEdSgy68qvIRVw7Ckl1YMPTV3
GFswHac3sG9VG8Zagi+fH3eUdBoERVqyR9ebN5Lz3jMY+FUCNuRsJbi/cFPd0miSf5H8sPMaS7p+
kB/ygBvCkKVFcgG4QCcxUmUW7i4wvpAyjUYwMDI4UBA2d2AY3Y+Ld+LQvbr8wbqmevAy+a3GV8cU
eXwbx1VrCXwzUcf7v88fHXjvjVNABYZGNGpnWnJY7O6LDTyU0nuUM+QRp0veaqeo232FBtJFVZe6
yVpdGXwa4Trq3Muj/EIeD39WwKNTCSCspyNI6wgDwUxU32gmEDicBev/ADAH2uzgr6HNRuxM5yeF
PJviaTldoeqU4VkIU940/hxKhA1jVYbzeCOJ/17LMn8QD/uFYZFUcYF2rUU8pTzkFCzaYkZABhbr
yyVROehyrYAXtOaIeD/+ThGJXGPrE+pLSl9EG7WvpAVuoB+fZm+/cu1vSSNaRZmKHLK1JUaG4Czq
qch2zqy8cm5X8aqoFa/cFvSk3c1XjUP+GTn8QVMKSXGUg7XDC7CTCZtb7ofyr7GyQTbF4a2S42dy
Ft7Gd2CcESH8JOUi9jinWxnX3Le+NK6rWYQ3Vox5wOCR4PHYHTe5jFYTWbQxVcl5lEnH/YNZzPIP
82wGSb34Asi8rW2MVPwldpFvwep2Q+0MpZH+xVc1+CcWQLqnnJ/Ao8fhRyWug424UycWN2h5dBg+
OLw4F7qdMO+vmDai61B8LwIHlC6hPF2TXjHI/1HjhBXHSxslof/U16p4SfLiGW/kpcncBtVHgZMP
GfgHjffJNFHM105a8aOh90jQC6DOMp9XGTqte1jAq8bulrihStG3BWm81maRtLE+L44dcxqbAByf
Wlu1T73rpDTACaxwlgQ5keVaWwbbj1w2/mr+sODHQBLWKI+2zN+oN9JNn/+xyPKrqU66B0+D//Wb
qYbafO5iNoyHAD3NYF0oIh5ptGkBKRxragFm3PXWPMD40qi9kRiSf3ez0bTwM5yjPOLx27fk5Tzb
K+xJRxSHru6dIhxON9ESLWfZ0nelMeTUxQGNK1dZjrJwy+5NodBz3D/PB3zqt8T7m4a1pqrXBdXt
wGMQo4ZH6rfs6IGLycBr51y5ubiQKr/JIIdsEEae7uuDoQzdJ++4G+47z2Dw5T7FlTgQpzV/y9Ok
LKcSvQwpbJIbMaXHBuw93BV6Su/PWoTB8q/JwZjO57HPykq90g3xjMN0EdmiOJzUOW6Jbw5ROnnb
+R+sNr0bHcQHKu710jQWkI7kaAKThw0WjTZmGq9vNrpKqlXn62iHcCTpxNdLABtTGeYEqaIlCIha
1U/XVWIS9c5CpBDr+C0po3P/xUXusnuUk/k/C4l4wvn8+qeFyvqrfKuFcHMdHHDCFLIipcmBruBK
a1ce4Yw0rAQYqkNF05CXC8QeQVrB8bTQqhZ9dC8EmljOobqUmHekfK1URow9hDSzFoL1O/PuATSd
u0YMr5HuXr0SqEhCp3vQWKVb1P80iDkaF4wAtZeTpsoBwJptZ8tDXIRtHB+sb+F4hEAJCCCyVXqO
9/f12kK8X2n7lvXCaBAryFfaMpwGF95ciiG/GFrBQHJO9xZ2nAAWadYQoNIFkZA0v4+kBGtemdrI
brDYjX1ym0XTjM/BnScag9K5AHivJnYYLf0cbzGSBrPOqS/VI13vU7ymFIjy24ycFoQIYtOya8QE
JjtAZRWLkE9QcHwpkq33Ha801G2QgHSYw4Df/GG4WVi8R+qFHu9VZ5KogDlySOO9/B1xBHmqQk2d
gDQIBuhkM1+i6RqQJEfHdaKboKgChPV4RkqqgmxSsCMclvIMEgmBPqk3phICGEzML8FxzoBaeHgL
Ufk298/9XG2VT6zV2evGJxmaAKgqUeuDLrRqdS/NzpxpYyJPZzg+kW8JcHQJgT6DqCWUISyOhuk8
MQmhoC/2YIcWZxFbk1AvKI2EflwRZk2ayGi6Ihds1h8Id0weKjnWlKL+dpiHU8gMiFK97p45x1WV
yB8f8XfvRdsF7BmbiAOxVsLXbJncOaNt81g95b9RYQRe60RguHng9vwCM5PJ9obN3NCOp+ZOQn5/
gKi9D6st0WtsicadGmRvPWybt0WodQVZPimoXxJg03+lEUF5YCTHuAAUBSB3cx0BvyWHZMYKYi6l
T39CfgXSwcfz1Q3guWcV0TyuuM/AwbqBUyhlNYngad3EKFwAOZD4Hhy5dR02kL+yrRzqsHAThMhQ
CZ2qs79kBI/EInbxdJf7MLmvyN9oMInjoxHHG1gcH6yZR+gMRBIJi8T0Nnijh5RMLTsLryWxU+Du
CQGIIv5AAGh/JwTgI0xr6Q2A6G4Gesnwk1hmoJFovGnRLiwzyT5BAR/+v6FfzYtiaq4n0Wnwa66S
+J6RhUTxDRIMh7HcMkMk06W2RtaYYqDpSYJwY43A6NsHD2fBUKEObh07XGd4DHzKNnv0yCtnkAY0
H/IazH6ci2/hoT37sopTkI4FzqwxBcdVg7nysWjDjOtbxJ60hzoROgaybdHk3rWkXxfEq9nU7KZq
RrX3qF8elJDApEJCHQ3u6V917hJK5lSzluy/4eRvF1beW43rd8X1CYSs+zAAT6+nUlPRiQqBPsxR
IzSB1N7zJBXszRha8+mWPPiKkfwVi65BPZWwcS3dNY0Czy/6jjA7yZgXsNjhnG7tBV3NFQFQuKZw
+mYGC3Th2A8M+vIm/lvLI3EvEbVfHXZE9IQ/Ty9VsZfyJPMPWSHL4mqGTzK4ckw9Bw+kW9Ad8ieU
eSYlIaJh7TxHak3+TrON4baknoph1vmpNH6zwK6Zh/6xMxiEotbpo5sJ2V/M2Fzof71V0rJsnsGR
bVvmPdCEUbl2QNEs9Y7pRHQbyQthwtKaWpG4eSng/zJUnWC+V37ynMKVmdp7epOSIxzbAPj9bod5
D7xPYe7FVcH4tgHach/jO7v3z7tYHwewP+lWjzHbx8xmSOBF31ZS1H/+5SoBs6o4sSGEWvrRH4s1
M69O63yc3dKUrSC3MBvwP67iDwE750TupNEa4qyAYjCimiTl3nl/vTSytKAA57YMzOFdEosjop7d
jnYZr1USFughZ7zW7sp/woVCfzIbH5gize1Ql92vqt+8PwX+QUQRSKdTDb9ElMBdosrvpW5Zqs3k
XcCBIyY4sCHpvkTEs1Bm77szAsMg9krpCJ6UpL6yu/pBs82JFuTfpLZ/YtznqiHwcgQSHAoyoMIB
sTGJNT+3RTWabRQmTY6dbCmejo0LxQ0D/7WFvh3zpJ8RAzKnbk8z5rylUhYy8P5dElZe5z61OC8E
Zn51Nz4D0+2mSQjSF8eStTiEfgNDu03NyRvPGBePB5CfSJlxeW/zT3CSSl5DsBDVSXq42mNEy/ji
dSIk5sQyH++4Pnk8qnjOlnKGyDvI9SiwLAZTlI7fUiedCyAtNDslTbPa2OlABtvAsGIGCtPkuTtc
7mdqsIlEWWun0Zlid07NloJcZskkEmCZ1AhHCbINhExeNTj3JcscYj5ZF2x60n/1zQKa/KeQ7hqQ
JrY+LsrGsrY6TGF3LrRVWKQIT4HMURkKnrEai+9mhab6a2Dc05uWwwHHbHMLTLPJTkwI3Bb8j1hP
3cpJfJ5BDCLHztUb5y4J7fGB6WqwZXG3n9h1kl+E8jIEZ1+WO/+adJM6uIMlAXl8t/IQuIlnY7WR
NhMru0NrDzlv2H6pbCJQhHYVk0fT1lMk8Nto8Zq1j1/EMlkZGt3hanw3nDzknmZDyf1E5thWVcW5
x5lAsMqfQ+yyQ/+krFYVnV21SvkuFKB/X5p0+p44wOIwdo8z+tFbyKCxbedxJg7ijxZGD7lvSPBE
yq4Th93pFEwMd7E4/2jtCS6Sd1NY1wGSxwU1WSpvVl7RYOBL7GAdU3WdrhEb1r5hgtVMhQm/rxPz
BNfy5XK/IeXYfGdqnN+HxOMpxSG3vMgRXqqkgJo/4zXvPo/+2McM/wLWPuBYg2ZLfXJgd0WoneBG
3AtJM6oaTPmO3e5nCAvc4tDnrCWO4e4u/BJRHr8szeW7Zq/QUrmGOKRLQk89BYKHVg5QgKXQc782
to95xQA9hJfmNX8uB4z2eha2Sh22hK4ZQyDV1sWkNO4HM3OAIkcdBlil/hk/z70bs8sRqCe3yt8V
8z7IaUDh/ckv/I4D6HgJrhjQUU0ctbtnqT+LkLzcAXyS+zjhLBxsiIRKe7Im8m0N4seoc2N3VUci
xyxn0Y+9PPWhDGtejiMpmAyKs2+yh7Z3qwz24k09IR+FwyZxp/AhAsDNx7f/kCeJroI2OTBFe/s0
t5+NCpEhUTuQCShMcrxhp7JzohhRrku4/e1NLnQCmptGQJMqtITVqK/MM6pzRFiwbrjrZD4yMaUS
vN8ePQjjAn7t/rOs6vZk4uX5CVo0EjRVtVBdIPKpaq8v30xY/toZPecf7mosJiIPOxQ7SI73pRQx
FwndK8s+FUrGWsz0BCa/RjZAOTAZl1AhxyFuLj5DCaf/rEJPE+dZK0CTKbSkYk6yOVU6O4ixbS4i
xk5+K+oBKZjozSk29nemh65Zqob38UMIEYl+hiQwlmX+NBYtwzTEFi/UnN53enB7eb7OOxtH6T63
eUYFaylSVObp8CZzt+9i3MIh1v8XNZvuqDSZVBJ8OCCpvTDEultqqNEcLx48kHwr1vl8WkK1Y5fO
I9QQOoWJvD97kG4k1C778K0upe/dZ1m8sFKP98mXCjWg1icOWmLGKTw44mjbIuRh0tZvYevK3jjz
BsZrQPcGeMYL/pd9PdmCAp4L0VCezIkz+Jh7WxctAhTWNaOK6ZKnx5SMR72sowCvi9VnYg5ksXaj
B4bFqwhJJTMAKkK2hd1md1DlLKf/cBhgQdfAYB0/mlGqBDQegK0sU2BqpSrUgKjKJtZrDCt9AHOG
PTqvhacE0KNXK0a/DtjNARlNlPNOLoyAZpsNfi4M8VfcsnM0c3T2BwMns5HHsBTsAUFtZyBHtx1N
s/NANNqHTrsXGAmHzqcqFU32QlEBsWIaRTjRY1ea07B2fVCC6D41m2RaLDEEOPSyqW5QdlfVvmWU
kgSBgZu5YfIBhDVqvy3UGSls7kgpHkDtdlzD5emR/Ar/vB+raZYUA/TFaOYBP4A52Po7dSLRujK8
1jRCF9AfF+m3KP4AIM9Jh1+3ae0JuX1tqvmIFQkSC2X3gU+uyZbP8p7PJf3AKccYdfiXPSCWmilh
9SmDsU6DlTxSQ1AdFLkWYGBOmRxXXVh8JH34dJyRgasaIsGHCUZcgjBlROac0k5ReVH4Lw1ruy5P
XAH3qio4z+IFZTpQxOO2bX0+fuZsrK1njYF3VRWD7xCv67+tPxC2kHxLPdJlcLSIUmYhK8mmpj2l
1RyX7eVGE1ccjESFbsDbTp+mklVGaA1PAeSgTR+NbtVGmnWb2FlPMB1uSplSftF1RYXJsWzYSeLG
2ERAMAntncGsn+GoIRseAODXQJUXOVC33zYu+humfP2xCLGSr15+GjxETQRaRhZpfll1qGUjZhdd
Gw8xA6KtnbbJDegeRLkkV2aPT8hSiCvJvRtnwHMWomE4mvfNCPK/cedSptsEEaY1dvOBwsF+Hh4/
o4DB423gJrLfrq0NwZAkN+/aEd1BRScHg5DTKWvyLRoUAsABnO6XdYM0vGRwH2DWYVIUrsdx3uUt
6ji6TdbYP+x+A0mEjHZUtiJsr0r4XcCwOhTDsy92Vn1dhQXjHK+MLVEO79uvQinlxI4yveJmIG2z
8lyKefygYOWARnJGe3VyoK+cZ9fIWRy93amPBslGKTNqoDpAMcTV+8mq/LomJWk+YUL5jeLokZI5
k6/PK8p4Ah4L+V00RcGjjOm+se5qll6CqETjI6kmgV7AR+YR1e0EQm7IYcyX3tYoUM+ZI1OP8HQ6
AAhF7vRf0JaKPMna8dCCwZIiUIrLNxm3axMuLfQCiy+8RhVf9Z9mkK4Pe06GE9OdB/Qbg20iGisw
RqlzgQK8Fto+SbYHVZx6hGjqljQi9abhY7m35Wwjp0ixUsj/cS6t88sgadB3o+SbrTzUDJd/GXOu
IGnAB778p8Yxvyck0cGC+T6B+78aVeaWx/XOSPN4i4x9JhkTIVlz4nETFYLzZToZZphwvv1ha9g1
xR0d7g2FWsLYQC9Gdn2JF6gkZeRWgFrFeZ6g1OHvViSeIhckFflmCSPkqjS4bPuzX6JengNYpYqG
v1Wf5Oo6cHoHDnLcKlLe8j2DESydd04akz2q8nFzz7L0ITm2OHLA5G8H+eltQlaFMHArDdaBWMBI
j/ckLDTBekDHb3PR2/cHoshpHHuiQ/8EhatjKBxBlFuso3A4GWrB+f/2kb63BLBSKvaTd4gATtmY
kY1PPK6fM14ek4BcHveLEkXCo0JWzthjNCTRfUawHPiYH1zGEGtcfQQah+zKBel0gTJqANJiR8Ey
7H+dHtpYiFmF8ZycBqd9BLc4oVJ6zcZqNcNI+gwwjyJQmc/6U6jqXuD1hiBzB7irdKgicz+12Fl5
E2VvdLob4iyFfSIWNpaXmTujc24i0Z+jLVel5jkKWDFcVaw1E5LrAkYtQmfpsU9Ph5V3IxVez0zl
iW3zqoRaEiJCaW/YNKGxc8g0wY/klH+9vqGNtmXt2bAzGc/qDhbCBB/RjvryleTm5SSG/6H2jstH
+D/LikIuSBPTm9W35QHRyvg2Z03her5u2DiYUxPSzcpW1CIpIokSlQG6iTuzFMC6smlj0O6IzZ2I
dfdDMhZQk4olz8JBzcGXtSJ0gFg9GRv1CIUQCVi7jNS8+RraSgviS/h3vlr0PB9eYGXIrpTnWzsV
ynBUu4oFEV2nAaASDNHyUKNhCil9XHz2biD8UUENgaoOf/mojxpjFnXA2Dyye+EGiCHV00+Odug4
ycIq0auDh44g/KpHH3nNFDEJmVGRyglFPhgwXE8OmI40osA7wp8BvlZ1K1r0NZz/SXBglCGRVJn8
clQIDKP3kG2Tw7mJ+PACEwCQ0wlci/LYhshHHNlMrjmON/lBBTXLCVxuw5phl9QyUTxnYcKB0cit
a+xlGjCmpXIEqPINWPfY4bHO+pxwq+KNwCXYLQkxuntMSNzszxQkGBBf/1BPLiWDMuXnTtI4ZjRC
mNV9NrzHzj/GnuXPrvgTmY6Ol0fCV/weQYMQEaPulz1AvAdaJ5pQMaT47d1xTO5pe0Z0uqXK7Izj
/80eUysOiwdhBldb/jYzud0cgnYQoukk/IKj928GD9iTIMehdsOOWNLDZpJExM+hmZSa88sQWVLh
E1IsTL9Hs6uqc+yy6/WQzUvwsXsbaVr1CMVJCPagc98UujuK5hyurvkP4t4Q0OFGDZjbrSv81iT5
vhs/kJMLkTW2ZjYnGpPffQkuDDPrKa6CmwHxi6Hb5/aLM3ejqgrFfQ75+R59DxajwQbw+CpFsKaR
QoNba78r54BM1L13lQCo0pFi6b8475MBxv7uQnyYGtH/rpZmvJ+nrzPbmmU8d4R1+g5PTamqGg8I
KYZapg3aeCy3Ttvtq6U3LifuzRUrfe/ZBk15kVwd8DgogdmGPmQtaKz4PLUXt3loQnyCyJEJyTWU
Mb6B3xAH8AGOchjUmCLAQ6uw0+FpDS/UVeFbyQ0/S26XfPX10LJBaZ0ESbGEiE2BM7ig5xHeoiad
3AEex0xC1R5KIiw9HmSI28VbcE5CjAYaWyEs8MISNCPpUBbaGYBl6APff0DpDypZrCz97JPLbiLS
TttAV+HC0bWw3qzDoj751q6niF0GbtQNdxYvIl3eUTnXVZ3y0bkRooIzlHB4fxM1b/UkQ8D8Z9OH
25AK0pelh/aqJmlBjNSTy+wsi4K/XOFoRTAKr9kVH6RlxUxlCkfzuR4q2lvdwiSAUFIKpdj9w48C
gCzeTBrTw4C2oeDj6zQODwR6Fo/dCpSRj/6zWfT0nMzVf2WIBVorheFFKDYvYnm9bM7pao8oxM2M
67CQtoKL0pk0QngrKOH6EpR++uLQTN4JVo8xArjYySHhIq90qmPTyX5Cm8+W7mLZrEALONtO+pbW
zhFA45sS5QY+jkGEPsDIIzHEavUhIRP7EfuM5tdgOXH8T/E+Vpeyiy872yKXqn0mTQEor7GGlAMv
7BBQ/8d1pnRTmLQ0a09eRn14wrgka/XMYz6HnLW4dvt33YKjXxfT/uKngdYtWmsQjwhEJbD+nodu
1tGeZJH+34CAZUZH7fBoO9uC9MOnfqWSDqgPjhZRi2OQfTeIY40umOinPSKFW+Y7UmoVo9gDiYv4
xy3taDttNgDDIKDF+tCvL2ukW96OsQJqD9iEJATObtCKb3OAkrDnvF2pg/8Jdw2Lh9m0MBpCu/89
GLxjp0EvRWHIhfwZNn2SR9yHj0kmm9csBe5JaAMBpLsf+/yShfMo30Oz8x+Q4cxk0c1dQ2bO+T05
a14y9XyUtFycukbHnogS6P3qiK0wRSPlhYzdXOSQpD5nOmcyli2H9qMP/Z1ikR5C+pmjygIPmGCw
+fWt9ucj10DWXE3ZYNz9ojyI63w97/HlBSBYyhyzBqEuDZS2wnFaInQhvyST/FdK2vuC574aLtej
1Ew207fQYF/U4bfgO4DyGeyb3HpdZf+KCSuPHnYObp1dfdoh7Ps87n555E7AAyVPVK7rYsHNBAYg
0SHMm+LZaQ+dtI2NYZCi1H7CEu5gwoZ4cRHPx3KE4QcHvv2FmJjrnJIqz9+QlRSbXawr3w7Obv2I
wqSYWni9e1E9zeLpeyyv5fINnVOud6FdXxLEJAcgDw60IkjJeLtnGKohuxebnn5WD+X2hUUrVKV8
V2E2+RgGG15O7utuGdpGGHU3P6nwlcg0aR16Rsvfp9MKgnQ8Ta9/ONQawZXv9ZLxmkbzI186kYmU
hTDBvrA6eMl6qW8c1O/AmYY8aDnCTXsfAalGgT3J/GHzR/6xC/qCSR8lz7TOvGMpqxESsahS7QXA
3SL+LfhcX+7zz5DwYv/lf4ls9ic9aqkfAEBg5+WiIXnzOcpBhO+wuKDUy6Hlc4NeiH9YDDNKo7J2
gyw0/ifL6M2aRDIijTSFupIWSant9bQICiT1hSYlzGxTYVx8NLXd2rVjZf6sG5+uuJFkcyckofeM
RqdzflewwgV6hIxIADFqNHogDDFL08RKL5FNjXKMl9Z315W1U+oXpE7zHyNbGqDYKt1HpHBT9mbt
XPVO2a79uByN6VZ4CXhILbkGVK0C4H+vDGwzt9f8fI/5CYfu7f4Io36hySRv6s7+ALHuqQjeNpDO
W0JVl7rmwRzB9tyXsuf3gV3OcHmi6mucJ4w2J7JY4zb3e25ZSZkOwq6yuZ9ZrdBhlSDwZcKX31ag
XOhDmE5AfYNwnAzoo/V4rP5/ZIzcsKRwhvKgGhPg3uy/V58efXZZ7gJXC10bHiVdABdHSEO2Dcwb
EE+h6y7POLUtGD68Sf89KR2NgQ+Ktt4NSAQ4ztdT/nGdE0aejGDKoI+czoDrd2xvZLeU/b1UQHb6
Ury4h2DV9WjWv7LlKVxhP50GLwnCuZwcuZipap+d7dwD826ctfVn1PSxrYw4awwYb6epFKJJl5w0
hSDR6x4O+M3jMkid/yViYQbrCpVonrqhyYiPFn3NqFsrPijN71zyDuhPps/jh19iq71MThHhMuHl
o3iQSKmGuSS3+RnYXsa19NVTl8ZiNQ4bzunMjQMs3MyGQCwtUIasZSPjusEx3fpuchuagVUdrLYg
cN0IwuLyillp9SsK5PLq8Fq0W7XsfFAzcrDl+/gV2Ti8Gp0BK25ztS9CEVHEXoh67RwFBC78oGQN
BbwCmMSdfCkobuf+9Tbe4qmj0Gf2oDKSta4QXt1NKdrFZmh5dtTM60f+F0OsTULzLAPP+yk56vnF
6KDzpYbMEZ0w5foxsf/LVUumZwpug3X80v/c+jfzweR0gwbF/31hZqWbAPWjgS5gBk/eNj00tnDi
jCkxrJjTQlNQF/QmOKQNMZb+iGlHRZFpgKZ4+71nzT6Rgp90T6hBOGgnLWZY9KJxfq7H83qvbo0Q
MKWB1jMzIbnsXGt5iXTqCrjuH/hI4BKqpPpclYy8oDFAUFbAqyDC+p7fOqfDnI/MycM449rw/PHX
wAH0wmvjS+Pik4Qp7VVKrKyfRLRZonvFTl9IzjiwQOxFT3FL7e8E9l0HoR90Od7LyxLxQbQxQpQl
aHgE1KgUigvWB5fSC/UluyLQhjKcn1fJQ2vuCzSGAfFPOijc7a5dFaqD1XLAi8LEDrzbBDs3vG6d
57QOglX2z+OzT5mG2GE6jxaEwVv0ObjET4he5bfArGm+IAiLMSfYvW25lBpzE5rB2vibrd0vMz+A
CMiHz00DZ6LQCNTTVeibalBEE8zQPDjkbqeSwllmP6C38cRVWdXcznG1C8DilQqIZGrxrxeZaN6y
aYEzQ2inNqdHsIAyokvqShzThtHv+Nt+zc5hyXxHmYqYBiwSJt0T4tQ9htrhg2iVN+TOLITkPp/Z
1d9lFaAlul/acL7kkzEpQNBM1Nj3WjMm62xCPdTRnqQ2DXs1cJaUwBPK3ROrJGuZg1fM7lp24zjk
unUenIcQ2Cwq4bYyjC2ctk17P8um/z/gfKZYkC7AMrYa/hOE4dU5PLcKb0tBuiFQcjoAn9XIKfXt
az9RrALUlc9/YMscyf+A4BtIP48qhMCGxpcKnmVnX52k1KbiU1IQ/+yH5qFlq/d4+82xVooXtsik
WL/HMSfmEx0Qf9kHVePwCn1Q7k1zwvdb/MbEDS+xeATnOtKBEcYvcc9WdZirS+bUIQC+FlOY4PQN
kUDKPW6zUQJ+v8dTG6mwwfauf/6VJH8MVkOVVGHMm7mioQYPuB1IkB5P6/wD3nsv/LtpRVonTIw0
5vQKlfQzX/7P3Z1ifU1afQLCX+4KhDAIXHG4GgSaH42/uT2J7Sa4ZVqc2AIeESAlFHTKg/btz2V2
ba0VFdYZoTbWA7QbY/zh4olwHy/4UXmUjyPrJ6KhfzEtJ2Rx0WaBoXocAdEBryKJF2+8FwrmfSzb
sI/XE8DXGuNmyhQfPhuEvX4MST5/SxbDrgLBz7JGmEIMkYBr4T5ACPR1jxtzG3JqMqlp2Qc0L/b9
67ziCYwGZHPBqmYMk1H77SuQWruQm6NS/LqD1Fh6VFsSLq0ZEAHY8r1ZSzjhRyQ7Cvo9EctaQwpK
xO4/7kMzEzvQIR91IPds+Ne0kiWLKlDK21iwlXThcYbeu1iELSlOsTi7fk5N4h4STiGmF4jq+e4O
bUiDSBza2LgcYSf5L5DAX+eQbWjRiG8oBS/Q6y3XtMOJlHOiqXYujRHYTt47dG1IMI0EoOYy8gJp
yiKraOT+iiHuKc4aT7OnOfyHjnL6xI4bNVlNkxrGy2TsWEhG2JUJsFG3Xm5Kn/FqCcUq3TZZsryy
lxoa7+ruqb3qMMK3CQAcOl1sKLRhsznu0qklXbLIRErKvYO02FTgiEVeHg4Xb5MfrWkssXWx5D1w
3U4mDnW6bmS050cL8B59uf+nhCZUkYdSM3/Oy81e0gzG9nJ11/uKPrWAk6Gtv3c6PaH1d0DImO0e
1gXO54/xAWYxA7iZapjHVVyjrHRtBPg8r0uBihVw6cxyeXGrSSwNxbNJ7bRgxE+hPhyCLrgAWpk0
zqUsN73fCS4FZH9ZFN56DfmnUKF913wc41p0UHc+ZmEes+oaOTx5lsF08e62RgfZPQ8B4YeCSRjK
+biTbrJQGYrt5lUQk5VS2OVI7JYPxqom64ViuMSziqbq13dyJIC7j/1ri8CtoWBSB/abNMcogUYq
evhJ5sBuUNdfjNOXHB/74XecLtax4sJVrM1n5u/v8Nb8u5Zo4qAiSEQjurwIyxOF5IQuifEtcrc+
D4n0mRCLa7HcqFjmjNT39p9XtRlrflas61m1XHBD63pn3nriMN+voobv7aRBdH61Wu/X3KjCEUd/
ojF0f2WEYr3s0wuBpyODhsfAWgweUgfI+wLx3aKVBbAG7WhyZ3BOu2wUEgppD5wzdkvZBSnej2cJ
xqH4N3bJ90B8ZYrqaYxFe9kHFyA5My6Vv9sV4qgjyA7VuW0RBHtTOeoNJKRhKrEOslJD4Ug4u5w6
kg3lwZaPXr1TtaNWsdqk1wPc5vAlcFzHyZ/1giZ0wFTif5OHqnCHPvpmdWFtLeBsKuCHm8vWaDYD
MZXy5Ck80rR5tnaBi2PCCiB1sn03j/ex9K5U+uFUL/wR7AX2MH5wYkeoUb31y6V5l3zNnhf2+Kb6
Qf715oUEZ73ZGtTny0VAV7rC7scWMNRBvaSR+kR2CQMyBj9hXkcpK51GcBRYcQsWd1uKd1vKJ1HG
c/Vb1z9trmpYOVVlZWv+UrgiBVTTSejS0UrqeiuATVlXVH5iLWMXQ3LQ5PAXQ2/mslonFMO8sedG
G35NGKh7HJDV5u1hM4n4LL3mjSPCLy58YstnXmtYJibL468p1Z0dE0GbaNfM2EaiTduEZV0vqTm7
zfq6LbYhgqUcOLwxhLXwWpNKIPFw9pYn1O4AsOiUS47r0aBo21JXv98V0WFfTpGR0uwp1omyAh2X
cO9/0kE5dWkzwzqFk4ldhVB0KjHxoawBZclR3Iy45+YNQqnEerTnSsmOnv6H4o3DB2wugpL0lViG
Wy37AOt8jCQraKbsSs8cd9Fdk8T4TtlioB6sJYlBAd3tZvyqHImq8m3GlHx+RVe3JHooRikdzlbq
m1/1oPRM5G05C5O/8h0IFCrPtK7mUVl64npb+1nHy+wmYJxsIMY/chjkIeHF96k7YD5AM0hmp8X3
ukydRfEUQPRpoOjuCGkH17E4pp/L5dRxHdlW7omI/XKra+T9NHaq8cx/USxgkvT1B4V3zsOZstHr
y1f4Oa1wEQKemB3HxjeBX2GVyrBkdTnOuYWCyZTcbcQfkKfqSiAsyVXEdlJiXj9D9ZzxAx/Pz9js
yfFPCblr3PB6+UqbfOo1YAm65S92kCLpSaFmJco6qRtzSG8SiP+/vwOXZapdH4lDF2jXvRI5oOQD
CKFc55qawheUFw9yz3Ib1GsTfzzj1F9QkVZOoPin4qm9NyilqKBdWtuzekRZXGzXec6uu5MzqHsz
A3Nj/0m946fljJIFmMuTHDnNc34VqFvuVQ14uXmFqPakyt8Ebj9fhcsM1nGEiSzPSO3mRlxY73yy
eio1Jn7WtWeSJoQCNnKbKUJE89gO5AFLjlVmr745c19/WfYMHiguUjwmROmFRQmzsLJL6EHXGkRG
2iVak5a1ZNd2xLp7g51E859YpA3G2ahNDscsRmfvDaTD+Vv6DleROw20iqstdq9u8tEoRlJvZxSL
g4r5hgirwaATfvcb1EZY2lO5ZQV2eGp7EmRnZHeTZvTRpnIkQ8tJy/5kzVxd7NecLz3m22sDiEMV
/eI1wZvOR2td2I4TO95Jn5Q/U064NI7eeZy6hYnz3sjsy8riLQxCILV616owHLHNHycYuBqFoU6I
NCmxbIZtlP0MQygo+V3Tehf91pVVTRAh0X2pFN5/dG2xQZdoEOrJ+i5NeVl6jkoa0Cslb6/b8ZvE
PJc+wzEwUj2b7juWdg8BEJVxRTvcgZjfag0aecSwwM0t5UN6DiyAYG1514fKMVtiDHg87jkJ1VXV
RezKVgdM8FliT4GxhtJktewwDiSfsfhg6SAfRRw+gjxnmRNKN+1E6QKvTQQqTHru01Z7N/VBD5Me
/gQCuEnjQx0hSN5WEEwuhzSckdF3KwQTi1o28/lOuTZ4kRiNVclPvO1SeWY+yCynbI1lWLzsa9NI
+u9/Xnbxe/UEmLvL0HySqRN7d0CpX4PImEXZRAewfJtBeXkSttS1K+0NrOBBHtPodrYJGnaB1i5S
7tSimO52i+Mvg2VE32EQ42WHWgO3O0jj87KS3Kc4xWCvXtjMQodPHnjE5MvtWoKr8DTiBErV6xwO
eiUPfUi8Z4Zxbx7Pd4AGDPDc0xg+FdoX5bPrd2GyNb4EKMTpkNMQ1++IU6YTV1zwpfr+dg8kcZPn
lAo7EaO7ISffxLW58voprIUJuZ/hYj8Zbaqh/iJ6lD/RjThvCNRsvep7pzj6ckAiWzuMUjW4oq6W
UTOM5Occ+jnDFfzyMl91nTbVmdfqgH/EDAmVpT1eyaHf1cvFxiEisTtdn00gxzDcDhzta1WFHoAN
hq9KRmUbF0LtuECWExLPfnPtc4eukomr9d1AXHigGYPbqxcTV0xlT/hWITE9z81ftEjGapkYbaD7
pzV2lCfGff0k5mZak21RP9ZcT/aOVQ7fXXKjMvXLEF8BPudxq0kWFLKQN5C5gR79laR/21eA5Fvi
V/qSskUE73BeTRN3HBhvnTXER+j4eG6ga61gcZafhcA7C458kFBtaQq//yT9wihFnQIw6B/Qcq5l
BHZeJpVGIH74zrmukKtCr0K/IekDNYOLDJudLFyl03nx4wZObZhMO90X0W/n8wdvS3WkUbRyPnEc
tyl+lsNfhMersIDTbaQB9eD8gCdRvGB+Hvl0XsBT//0xOKsUUzfiaJbu2ilj8GINbg94os5C2K51
CGaROC/MJhyTznV+fKDADvYlCLPq9gwUdVsWgCI0T0y8e4XvyALtErT3VHarUALOSP+OhmNP7AxW
/miK/kANO56/ZhDdyjpDatVH4fDYsTlcC9iNcZFk08GwCg7Otlq8YxYfXE5wcr8p1bcxyYbHYSYl
XflYKm8SKxzfvmuWDJEEf5dMeeyG9w+qpmuiPlSvYVLjRIKJyaAcJsKuRSw6bPNNwzjqqOr3b1/v
ZgrDQb4cXt4KujQAzseEhpiW8zlOuCOA2FhPCWAy83BNQZ1dZ2283pvbY9Wg/zVzRDHRPtW1b9ul
EZjh03bYeMZMHTVIGwop7t0JGUADHAGi0zIV0ri8QaQ4eV2Z8D8x+P/W2VHAeR89MTQRyBUq+TMA
VhbkqSvZrCVrrmr4wCiUhzmyoxVdwLZ/K3PT0wVc5fMnqdP5j79oqSGt67ZWx7IhhZtVz+/wjBSZ
iuF8jZuMicxZdgxUV3hiaVFA4cAjQ+1X+2RXSrCIvVPwSR+u7xjm+iBOviYQVCkBkN7/FhrrnTbq
KDdAlH620SUtD8/Slpro0yTwyNdDleApGsMdSb49cNeZQipm1HxKW3oT4uZpaRgFYvpJ0Mh30fM9
FQ/rI1zbjIZsKnCVH3EZhcnE3Gf96YAxVUei8/Ev+r291m7sd7G3t0CYhLnxciveStib+seRBRJ2
xeujq6D2x8YtTIFbNq+BPgweQYLMaXMF7X8eovGr3hakYN7REKV83eM7DaqoZFi/AnlOWh+68gtr
MI8lTcCmzmn7WQ1Ny+sGULRjMo1ly5Ebwejn7wQuI58THiQgU5HgVbEm/uZY6F9YMz3W832BrxdQ
P2IBdTRSOvuG/R0OBWRQVK03ksgPeMh/XTPuQZeQ32UozSBz+fwXdwgb7/vtq2/GDaG8LMiPZT4g
u3HfmJncOC12LwWoo56jTzthIYvqJgjh3hrf4L8ZCefjXfekqE3zHfMGNEmPQVeLUp6l76kw97ch
6n1xS2nPhGkNJbZW4t4XHDMuL2wLbsLoY775BKSeuxAQm1alRtZOblI3/7HLKXtmyBdduKcfH5jy
7VfNBF/D8tHVvxtVlpmI6dwnFHpXAmSH1M7TebjnLIFrw+LEdV6Inewy4FYDb5EhSg0+gw9cXe9t
nwfqlPCg74ThuVPmmkV2tO3JVIjLnr+fiFGQJ5TubvGIpD2FLMMkDRhuNm7nKcERkeeCyI8yrQP4
EZ13Hjs0xEZJRHzl1BhAAmeE3VXBi2avLq+BnSTrRx+1FtFF0A2GmY+IvcAM6KuxIkVO3Hws4UPD
hs1tpbdQPf0jLpy2HqoohDTSvZdR0mnrENhMaRdMXUj3Cd+S9fg0Rb41W7J/TFkQzz5vsOGvU7Fh
FegSSbGJHIO/URlyMhU1HvzxBFep2fPETaCTbOwv2z4KjdUBf7ubF0zXQEi6+qQr1yE49gPxMCIv
HBadcEEwfVmzzi0poYLgAEWaoLjbYJmTjPaXDOW7oSUnCSImjKoz4WimDYI16GpzB7QQWAtbjq0q
1OKWfHhmQoIzOAP/pMXTFVZ1Py6I7kk14Uar2fC91iM6l9UpenpJ1wgkkHGqRh9LLHVghGLspFPC
cPHMuu/ugMTRsn490MbmqiJhDiqAHFUwyUWtHpEF0PGGLUny32P7y2XY16fyl82qCn3HE3gxyNle
VdJPOkf4mAHs4d4DrAYyblCWkpHTFsg+e44NcA2LS2io183aGEMrDEtY/RYobVzbmO9ilU+FOk6I
rG+2kuen0letUjhf7RO1dwkiRQdKq/maXKW+OnP+kosCX1s512jIdOB6T35AT8bhE6RpEJe25uBF
d3mPYjPYGDvu6sB9h5FJBJT51w9hWgnRwCfZxbdI/zV6NYS2wg9IroJvMLePLJEnYoFCQaaA7fzY
Z6ycAg1nTCzXsta5IhMHVypaKn0Bj5Qo5Xo/l7mMV99STdX1xSGaa1iTADDhcHDvGxnJXXdXYX4u
EQnZaEXcknQnnY4vL8XPr0v6DU7XbSn6/IFE/O/l52ZCaQGkuXGMuinw6fhAyXvsP2TLpNLtlmYX
YxdF8flCzjf9k1tXh1j2201Grw8l2d9YA7pyFF8BB68UmbgxPwJj7JsLNTyhSl/ddpA1fwfi9eZ7
GITkqm8WyA6W2m7BFeevPT0+eIAJKxh71LmT9ONSJEq6OPW85Qzu1AuqD0CSXIFGW97hO7FGmCeV
0MKIpXp3KBZICVbj44P8aQQ0vvpUgKI5gRSU66mEzJ8hbUOJjMG68byKqqBSse1fVCAjH2awKzQM
MRu5KPN9EbjIBgdi2IWWeCj+yrPwWmA8c3eItVHOKIuUtDeCw2tyVha9KwCYJ9T96nOO5iwtMCmv
oMdWTyxDUbKdKejqMfyFXN2++F10swFAf0dnXe33U9xZpA9HMIpcxMhn/uttB/RkEFCZsG63ywF9
HxxyWuO/WqltY9oOBCb+1Z7vMNlegnqoAjJWer7nYO4JdnUKS1X4JhHI7ktvDUPBkkqaibEiiVOL
Hmdj9RA82NmMhpPgIqaAUDMOwTlXHb2G/ISQQrqpmsCSe1tuyhiLPYCLe27bX8piu/+ihmJqoQ6c
bzFqdatuBU2Z+RtL9tuVgNqZUbaMYbz16iwUpJqF0bLgE+NxlTaeBP1LMWXheSD8T0q/Bfleh2wV
eJbAQzcXzklQD88c/XkLCJ05MqPFssT8M+T6y+lATBcfLYDZMqsipRvKgADfTlN5hanzVnuKjkz2
n4dCTB+852Ao0NV/k1Uy7kAK0s3+t8712Aw1WOAvZvp6XNKe/msf4p+jPyi72WBTteHwgL8Tw85K
VIsJnwOFmnNG1UuvK/NXJF2M2WyqjMhrE12CTuUAX1zWryd7zKBANgBbkiWptN0dy+3UpzyFQn82
8stb4OuKTpCHXrMXVO6WQL9zhf2YywbnSYBnrAgHu+lcdCXwH1RCTiTy92vs3NMEmjwgYPHCjXyh
TmGV3KnPUreTD01Z0r4YT1yRJsd3XqkYKTPms2lpURaHE0tK3w1Pd75y0TdBNvi323kVP0BUFGKP
egX8tQ5SF2/cRMPCSTjRKETeWnHlT22i9eY0p15U+aaP8upJfrkfSjhbiHQTWaP+vbZcmasr4Ce7
eWWHPaOXM6VfKy1AgWMwcMfLSW+TusCFq1rkBo62F36aqCbHRtfJygAYuRX7SihYo0t9j9knG7b6
yh8ZoyciYfyzjpwMLhLFrmw/JAPbVtIM1E6vMPeoqD7hgnwelkKU/PCSfrk81NBo499lBvvowReo
c+niS6RNz1kzqoWCBdLp/M+KXPHnJL7p8PzV/MXr00+Ht2M3i4Ah9zc1mnZqi7p2WBBz42+3ITog
9K6P55Ubph5jcs4auP4KHJUpJN1BgEtj2K/Lyu+js2IvGnQB+OL708zA94jc6vKwHNhpcaMtZR4t
oYjfGh52mtEkH19p1j8CFhx+FFBKmwToxaTAv6xOG2R4zmGJOeJTDi/gy/R50sOY83i1wUHGuAve
vGccDzb9Pa0DnXba3l7JBZRhS18QU0eVPRmLe5O+F8H1I8SiJEK6s6bv4lhupPZOR8EvyAY96wuZ
e5nl5Xjp4QYWAtk5+FG+IKdau4wR8bZJlvYjldF9ohUjbSMF5jXN6pasrAkYpGx8ucZuhSVhF6tD
6n+ocnFVZPXMW5nGMEIT2hF/zKTZoRyD5gbdaNhN7AjFG21IC36V1AEU9tta4R8/DY09a5YsBASl
mb2tuR90FhCNurfm1ctsODg7odyg/87uEZOpS/+cn81ib4pYbZFfNxC3L06ZYICyz4ohaWBloY0H
vrjcihNuuVk8gJe8+Kkfx5qB2bqhCj8zGAm7kB1UpH44Y+XINU78A9OpL2z+/Oiusjqf6Rm6P6EO
InJiLaPu2/DtdVhwnTI7oU0N492MGmTgVkePPjyJqLYhapIkOMsYQQjjLWvMELs+002vJKPHzYRj
lGfS1O/M84CeFw+CLTPgrBhdhvFoIynpLiWN/upRGQ2eQP1wt61EDu6s6ykmCoeDFVXbe4LzIm9q
yuiWMnXMlAxURb2XAa+1SPMmREH8P+8kmZfGT0V/QlFHb90M39zBsVeOKqq7WGmnrZQ6/pX00dJV
OwrCrhnYxLAvbngGpt6IjTQimcAOCygGl3JlS/tclVcr6DHaN9b4MKszPDLkAivFSZioxLLOXJA/
HYocDIXwTlzcdfarU46WW/5autfNUbBhDhhIbtbeSx8YoPPF7ZNMs3SPEpmN5Vn2xgXR1D/kbAJd
zbus/RulPbAsyOS+WqZpSOwNOKdMq1wkusg0kw8f6JlHIHkmX66U7VloyMdSE24CH6kxamNSHLDv
IHucNdWj5M2t4cW2o2FZy0sSuUptvbkjcpTYyq0qKTdF4eoK3QmVe4UEd46ywTRhGlK1XNVUHy4K
4pS7bwphLXHUxhBsdSQZwwx8uHEXiXFL7kGE4cEF7lQBBmo7MJtT9Rx0v72xOv5lwyq4DhBbw0te
j79NEInVHRH3Xl5up/FbakZAv+10iPHIaZEUx/JJgEBrRdQxcAl1nGF44NTliezOP4T9LITxUOfL
7J162EvRgjb2juZqSDD4Y/c5ugfBW0yuaRYby9VzSKVs+TAA/t+ecsB07CIQYi5sioneMrIxZqEl
Kr9AIRV8Gsyh5PwU5/zq2Hkq0HXJ2BszqFhQFLSRRiZ5jn3OKlzo0C06VgJvbnW1ET73aTwbh+XG
6xUC3sA1EYFU2Ok246L+ZuGc/Mz/JI+SoUS8gICT2OIuQAfj1QeNRLL5A139xe54/GMlaq1ZX2yR
xWWe3Xakyn4ZQn35Ma0zytbE7Du/ff83dwQekxspoJrDZQCY+mWp0aEPV0MhePV0UutZqEXrFn4Y
Dj/PFeC9W3E3M2agfCuFNRFSOPamGttL/3ucsYH47bhHDtcGeEulj655BPdaPh7n8DtxTEMDkXGn
6ET7X1WJIt2i5Yq9jfcY/IiDdYbowurZn9TDEIaZxqWVHhDQ+kWfeNLht8cjp71VVZ32kEW2W10n
lqufiVyvVT7dgLzXgpnGpQ/qUHw/73Zxs0G4VIk8r2vUEXHKJQcxsuhAuFAi08urp+oloXwn4s6X
22W5qq3wlIXggeOPTOEnkdHI2XP8zbxZ5WGaZAQkOwcjLrZu+oPIhHQSd6ri9RzUc1BYesBSMsof
cyN/jCp64UqfzqMvkP6iWfYLjnah9jTxQp35P7JJ1Z3NT20SzkEVrveOKc1LpnvF7Gm3/29WpfyK
+ZKp114HzuTaaOisWKE3qlJnzCLZl69uXhRXw8GOVKMIqX/Z2ue7eSgGS8E+gf333aJdgU45cHA5
S73mZU3geKYTDRRI0f4jEa1aGqnACu5Wh3L5v+s4DwY4fiee0EuaTMsE3KN8H6seOKZtcFzrbkM4
Rh9xZ7pBnUyoJ1NpGiTLOUG2/t63gwW1fGXJAZ48gsBczasN4oTjpvvvtE7uf5WhRQ5hQoN/sYyf
G+HJS2lcE3iaOHjATpMb1yLXJMFr0/Q5MMewDcGpdtlVfrFhkZDsYkCH+nAEN/OABBF+YaMvOjfB
YqAgXGd7ggDnZCBh+bRLcC+BwcdV5LnHKjzAcG1LE2viT4tGMtkSZeyQ097FrwJEjReUkUKqtrNH
ICD0FDBaWrhhLUuxV+ylA9kUl+21A2ud6c+sU86RV7eFHrzOVkMmF90e0GgqfTrY3R2rBfUNhVV2
4/SeGxgvRdaTd7rDdmZ0/pmXMZlU2cFzrg95CQl3Y6Gh43IsZizNi1oGaOIcpiapGt0uNS2f21bH
75lF19Chp2ouwPtGRDmdo5MvzMu+ljN8u+eArfDyLgsnK8p+V9YhgZvilQb6BITqdST+/GDxT1dE
8mwLvR2kKbphF/XzYyhyhPE/X0RyMcUAVrsPwPJkFQECj4B4xCCeHeLh/h0g0EargWfrvZNluODc
AhzSn3yKR916lwW9ybc2+2NYX3JS1LP2qrVv1dt8F1rWbby/YZGADaUpg1ISlDrV4Nz8VGbzrByf
L/wwFc8tlD6YTE/nfcMWFfTSXHZ8QrAOeAuag9bEXHSJkv35PN54QDRR+RY9+woI9+Mip4N8tphD
Fe8ddFNDlt9GHdLMlQ3DUkMROOQlGXmjyBrC9HlOUr62jx4ANPK4kZWUWy6HtmBCC97zKXakxSEQ
e5VtALavA41BTjDqIloWELFRw3Vss8ql1rAGvedWNQQfe7MZWup6Qcde41IIiKftwUQ+4OAuHuUB
R1XusrBlTv9iLdDCje4J6wgMGjEFoRkeoT3Tk6XuxXHloSlKEWnrGBzhmRMqUPBIlCXunkuyAiXH
s6PZIqO6hXVP4JUIhjN9vCF8kyDIcHSn1HwPT3Yc4VBea6KHpKri1If6NyF8tJSvhu4uDwI+cVyv
doIyHVuzzwAJ6zfZl3cFh6fJmuvgSPwORGk/LqpeWCLeJNQFVACWH/QjZsoWxNBmOAs7rFkidn6F
ZIKNYW86N07kVBIuamCimurXuLUe3DWiMCi1vdO/R5zXwrcjc8j5pXmIDF/LU+yRQufLtv0yBq8X
wy/ldp8Q1VhlZbYyz8coJyqlS30rAnTwAV90HK/AXFbkZmm8PQvbXf5YEk0UvsdWwqMh7efIvWd3
jPcu3Kbd+OXmYIfRtD1z095kT3/JlUOVnaeLG9H8uiw1KrUDGxm6vw8OsDVUgqLamCj/uoeYsfe7
cBuiPZYFoA9K/BlKBTnKwsZmgwRGt9eP1PmXsQpxauW5nbE1Ha8PUGp+f3WLLNFtz4HiL7GXeEzq
o9F6qasZyU3IS1H8biibkRD3pmsXRXWp/wtqlsUBFkOC8vaUP8ttoTDf97Z7s/DjMm+nGhMkcjBV
shMNvvsmtFamqxFlzv8PD9betol1BodG1mCbiFML+qIVQpF5pdPe+Ec+wWCPDBJWHzKkQuf9GJqM
FuJ48e+EoKnoRy3r9F1mter0ijrtgAQZ8roYmg+5uAsIT7DInPAjJbhEVuILwMFFjrmf8aO2UIkC
MxSeh2z4zfeRobE1sur6lEFE4iDW7FdaFzZfKV0SRCRxp/diW6zPFaswy1osRfDidhyD1ZaClEzw
+BufdhjNuzp3Z8dCy6ese+/0FVsiQ2sP5vF/CzMuL1aaKDIFjblkeKtup/HCv3QBjeyhT/x3yQfZ
0H5+80CBW/Bqw0EjYEFJWrakJXhvyQnsqaIrvxLtWGWlxsJgSEtxhK/rW/zEjxNvkMeT+U+w9k/B
xcTnzuzEfpb1e/DNHan0lc3A17DSM9xOnCknfA1EypFW7MWFsAc1kvRHznPMEUheFprQopcQ90zq
SfjKakSR73I9Fi1jovWItLHoeJFrqPZnFVd1SwZbcUxTyZAFG2lwHYhLcx8VnjuGyp4zT1pengIF
yLZNgFLp+udi5gJiR6hSFBRLxPqbkb69/5/HOi1+NREvDlBaRmnddC3KB40w4vLKAUhB2vlylLDO
dmz35K6l+TCHlwfCwDtG8gm8A0i4UHhrd99SrNgojKqCy0METpbKqnLiCF6wQySmzZzfrusz03tK
bswcHsGOBlj/i1coRBmTNOdseFF7TJmlBEMOuiVDcDFdNGj1WcXzUVT1H3ImhEl3OD7tGdOZXy/0
LRVCiCxbsKWwY3J1g07ql/K1PMax/g2kPAn5zd6rjpWDMnkLNHgYDlphqs5grFQxu2InMWy/NsuQ
2clNEtGFagaUDDr/uBXuTJRhNnsJNmj/F6dkMDAFqW76vtl93r6zmNk8ikP70q7JF+/UHArm2ND7
csVG0u2F12iVxhvb48BpCxmH+Af1JRS+5w++XMsVTRe1fCBTc9GWzO02BgvX8Nrtic5IZiuHPhWS
J4SroPU8lgZUL87OBXOl5I65phLqFFiWtZBKXyORyp9m48dpPxs98XtKirp7z8OoS/xL6r3TMuTJ
u4Ye7w1LZKJRuQXV/Iodo9X74FwfpSmsw/m2+9imvV9mlAYAMJqjv+3ZmXg1jGYAte/nyunlVJXy
TK1RTiNjHvYaYapL8/QvA6TFNoPScoF08zgkw59KSZyWE0U3k+A5uYljPVZgW6w7mpvRK3Ry4Sv/
2mXPhnttiRsOjwAU7PZzuL5z8ft9TV74jkd/bhkd7xzNSsg4LQbFmZZ5WXfXNAfPvCJhKfiq7vpC
1LtFkAM02kLI4ukXQVKNVNiJhemJEgmb2We8JfLWdYYnytiWT0BprsslaiqhT4R7dAkhMxgUvSRj
9mnVUTLNZLtV7x7tto3LnZRQsYFAWk7XIi3LMHjtrjbFIY957hEBSBinlRsGyuKTJwYOWmkzr0Ds
wmHP/UJAd9KJC2Mt2Pktf/o2c+d8w1dkWy4T3/4JICndx0GBysXetKbt8b8GhPI70wxuHVsWVDqH
pyTf6oamq6vur4ZhkwMN25/+Onjb5BlKY3vJE8avfx8u0rilq60G8PWRPJ+BcYcfkWhSQVRytBG7
OcZgz5GE9Q+QJNS2fbXhQ9t73+4caVZFq1sSk2ft1uKfGpq4vNJmI4d6GGRoOAk+N5NBRdrGt73X
Bw+xHSbWWgUDCK6TarZl+P/I0xKVNZ5an+dkmPUTEM0GrXtkd8LftfZDxbQPXF1fI7Cd/mzWjSx3
tmo5dI0xTC3G9pNVeh+eJVoUJkidFofptlWc/QZqilLsIJnCT8ZCRioZeAh3e4/Hx9HJ5EvSuFlG
J80w/riKxH71tLRFjvt9x7kgSv1znUZCsZNVgsr0mwpKIYq9JY4MPxX9X5EsICmn49X6Mnx1ffdj
xIQvI3tjYYl3u7ikZ9FPZETZe6E9RbbIlJsDr+fFqDsuKXAg6+9vcMHU+0apymNXJ71PiiTdEAX7
nwRlQktBYstSdsIk3IMVnyr3gqp59qlr6UK3hF5HHrFfkQiOIX0cZrSEUoASA5liQlI/hke7ZmGF
WECdyxNNrmIr2TN5rKidYmyPi9l1s4MpmkJzCQaFZoG9IxVCtheaRm5Iwi75MNR8Lk38eN4hh1uX
TuyluBScVNigf6shlh2TdNnUgaEv1zrv3EcYuZFwGJgBRT1IRRGHocVLkC6jUPqF6h54V7ajxFz5
JgrKNWnLeX35pzXCQ8/xOKSBYWe42nH77qTeCeASfL1cin6Ryluw97AMozqJFmZcHN1rxIbrAOlh
wsXRIewIc8UrVbpnV6Hd/1I831ULiXldWltJiMYXtOR1ek/YysG72l1Jz5N9loSJPKh7vTzvJGM7
hgCW7oRIi+C+QgOi9InCbpLE6b027OOwEdmF8HAhan+g1F4Ohsn14EhQClrltqqsSD8M7/c5dwC6
DmP+T7wTrv3paGEfsJ2oyIOM7LsOJKVrwxYnt88gVnK4guPv5tllvkND1H3Kony8GhVtHCMP63wh
fk7lIoYkoQrac31jjmWSI3YUMWayupVqI32uRK1K8f9+d6+0ly2aseMoiFY6dV/StrdVDVTQsVnL
D8PJ1uvSODhabBDYZPDHa5AWS7/1EWEF2ZmBQU/XfQHixMQnwJZfJUvIgfd7G8aIA2xymcwYtxPD
mqLaSlK6Cn73IHFlhZSkKm2HT+kFGe24VQd/t8EAlG8YGBTY6sTk/7Bt/pPtBxH807zohiyVN4sQ
N8n0iHO3LumiM+UjvN0mm5hKnZiE8Xy7iFKPqJhgJs4pYuEfP2E55wYlb0YBkd+9aorMOr4uJp+c
xqAs8swhfDhCC5vyI8A2ronPNQamJdivnSmodKqZaJlNlDV8PNt0K2Y4Z5tu41zc/CSN84vv+qTR
Aw76i6gsAoYFWtZbwN/BWbV7ZQENAgxKEikYawjh/cjHxiaZiEnkwfTVM0uMIisKTuXtm7NQc7k0
1dFx1qPE93EeP4DtbW5naJNzK1oITwH8uh+B/ctU1ckDC9EKnGqrUP6JwLv1HLaNAW0JrGlIFOk/
RCbDjPxCdVqzb+9kioTKZ3ll5sjuZyS5PEh9vNxJvk7a6ZnJ/y9LJxL0uaTOq4zwAoZC7/a1ntWH
VqSRvCws8Nhax1aWKv6eBAKEQd3rgrlHBfceE5uEsi5foaZA0TmZjqoWxLjMyz95YQAWVYc1cCbX
rjxGD7prDdn0ARni62/xpWTr5uhJc0XYkLSvbHECotAj9mDr7pjt77V4GfA7232lBzTXEJwKK1Z0
QC52rynx0RNMA9zuU3KiePLe/FSwhQb6SkaPnyPip0FKRe5vEEOioe1zwIdHky7O4N7m07nhNhFI
zSNj6BCX908PBiJQ0SpgBEfONAE/Br9o1JS8isx6n6nzSUZA84IPcC7jns5+Cha3PhTPU0WZ0B/p
Q0wOJXI/zVd7OlVnUuXj2Dv9gqJV1uO1ryOwAkDR1aCQspKU6CQ6ozQq2iUCEhkGPaCqRS9b4a87
S4TzjytyMMSqw1kZljJqoeNCCQyk8Jo6PlZHpHiNYoaopc4oKGBRPmfTJDEaT4HOkMrv4L5YZ5tq
S6JGTTyb7W192OzixUFkTrqXZlwgscKslVQflwEM8fimqMfY/soIATkIdv8algv6vL7rL5PRFkfW
vK2+pNXFBGagsM2axBNkJp6kGoInSwOkjl8nw6pqO9Hfw92ehh0CLGjoaKlzoJMgWYSAjLBFpufK
wnaZtwFFzhwRSqeCwsXEpWRvsBOVOFB39WsVPAXiyC+Erp9i/rmiuRJko29k8CexwsCqeL8VrkVb
MHNMOiEXtb498oIWKOLhRxbe7DCQyWPcREBSdlUMM13FoKM06xkXbf7Zogt08TLSbNPDN/Pzywsi
ZbaxkGkgHVrzyrkcMk9A2Tdjbr5xQrY1op09dVNqTVzyBECTdbPxi5z+n6Gu5wcNDIcK2LNG1XGW
108a1nGTIengaOr4EvADW4h4eTlSQ57LRkltSAk2FgRy1+xgeWWivS5/4sROS0h/38GPiXaof5oW
YbA3NRcBsJ1imV4gR6zOlGzayJsS9gbWIDEj3MWn9vZjDzeZa2uz5SrllqHMT/uuu42DDahHOEK/
pbPp+FYFwABjrBDuHIPFBgxOn8mfo0WUvIGbuitSPfQkED9P8q3s4GSxCtrjnB7Y1cI7hN+LwdK2
eF/YvT0MgxPGfwad+gvYlf2ggeTK6hsAh8YJzzMxS4qPmAZrdSURE7ap0NA2m9HdmzyztgqDZRo1
g97SI1K05KzYSVc+HRtIGkmmBoaiCj2y4V6rYfT6Yf06o/rO1T8cqnbssIBwJkneHkEMpRZRL1LL
KRz2MoZuNGxf/7+TkCnvP4rxTOgCRdbyolved6Z9pmxE+SDQIUGUxSE8JkBoGr9jVlNioTOHhkaC
1Od6gt9WlOWHDIxmOIlSq8kqwV1/lxBLBpnrczTNTMhAmSBGH8ngc3PD1VNIfamry6pE1vqzNtsh
QDOwAca8I+g/2jHJpGAQTWxBljp/p1R2SHSOG6Br9S6xTLvW1mkQgI/zfhq83Rz7IRbP+CrVI4pg
d8762R4G5CN1779iluHF1Gyvin5jOUmy0o2ufavGunj7YUj/lUZKNpEU5MmgL8PbVu6KcpJMBMIT
8bJMEHGupSAtYeYoBrSATDbOMgftj4JvdFeSy9CUZE5hCCrK+g/IAoUramJ8DK3LMiCZ6dc1mOLx
xy1dhOasRQOn3pDeRf3e1oGbcO5Gt7dur67H3bfsBqLj4lE/XGuW4D0koEeHtQ/by9G4BgEDPsBH
UQXR28Wx3OaS1sY7sff9bPg6KepRYcQFxTdrIOqFkPLxPA6esxyh3tOhyCGS1bJbw+CPNqvlrmCK
ajDnrDbO7zWsR78pLELI6vE4yzKCVVXhhqV9yWAQCnEpu9QQzSM821erazlRE4l8YWzQv/dcsqPD
eJAEA6ItNstcTV+j0LNKajekNcqzPXSDd4IX2Op9GKf3tU3Y1V3Zs3yH6ueLQ55DITGo4HZlZra4
L80IdB/qPRz/aztAw7Nn0SP9oKKlPSZ/GNabQUOOyJQGWF5A0Up5ZzP9mGlFnD5Tv8C+9EHMMv0R
cFV9Gw3ROUlbYZ72zy3E+BMOaQLkas5ws+e3nSYqCGq1LqfSSCAVGrnfacjd/QctZKl6T3I1eTqr
pbBZVA/WUhSaqkTch4E5hfFN/ZnQh1l/E8v4bCVZabpN+haZsBvJ39DwWE/3fGdx/oEMf0dFthkJ
QgUIDxtZOyYSOYksrr0xWVT4iOUUKYh/ugIPTZ6o3AMGjXCi9B7S3IrNByIYXqoOoBAZj14g5YFJ
XQ5IAaSBajxtdT73B0qEFeVAEXAX8683LQNPEZlr60F223Ov8v176feY6x9fk6PBzbbFJJZ9DBr6
iWqcWXlM3aaFif9WkMAiokEiJ+ZEAmOOv7ceCPH6HOFv6Osykio+NAS0uMBnWZpCic+Yro6xzlY2
aJCh6f0gwb7cp/6GcC7JB2yl1lG9fa3F2xCOR5tkoczTjvX+shsjKBFQjS4+KMddwKHiQH2xcaah
YwDMpFsPKbeNdARF0ZiiJaF5jMU3pkxMRorYSmYJj9EwPpACbL+v+KNqicgDc/3zAK+b2e6gnPOi
N1RTmmP6xlWOJQhPrvwDBLwu1CiplW9tBP0QBRYcb+AxhAz9wqiOfWOYh+ZXMtpEAiSzv+8NE1lH
03HEyKHJI40WaMSH94ktBWUrvOJh4LX+bT4jzTYIvR5b2hU1ofBK2KsUKrzfIlac0gYzIAN859ra
FGbpUa9JTAYb3HzTk2jrtY152/ZE7Sytv3RR2Y1XJvOvJpm2+1GwehmyOyxUPZzHAape4Zawl4hH
rTfQkm3D8HxMAk/Rl2VVCiYSmvoBGDSR8cy2sC+6TQQduKQUEhrVX/QrLxTBin+XZEAxlytN3Cnl
xnubmChiKgPMkohfI8zC50VPlaSznZ9tlwPPLoNlr9anfotHAc57/9yGe7KLY647KUcmAi39SSOO
GznCApTEp3suduO1oIWbM8S1Rb5qhDpl+TadmFRWE7e9nhlBjMYtEYp0EoW1jATUoursu5TAg0KK
/6Cfhf/MJ6zLAy8zpYa/XX7u3qGdFt8fyLDhAfSa3vOj3OjwdAE/sjUEJwthyQeUS1iufSOa6xFk
+NyimYXgzTsgKjgE0Ok6d97/nI/quaE461hH2WCkJqeUXhYFNIuyA5OfDl9JdsmemVgu3IJoDEMU
U6iw/l6gzuXEGO+hORddfSwfG0B3AaNAT7aCvYT4c3b8bXa+JaEr2w3FkU8fGU0LVxY3N8AqtHPh
rbGVIMZmDsIiHJ7O9wYiipM4T2wY4whQoHOc2l+AQwrtFJ8tB40/3FafOWjfMueY86fzQBf7bdGe
u2OeXJ3sKzHCFBG83ut48wOabaBNJuKAyEkcyUN6rIJiMJ3IXPUCWRgoMueQiF+ASDFm4VTHEc2k
NIBPoZT+PJeF8GoqwXwjsPWmvLKezzhSb9MJafgwBBP7SYap66T8D1J88qs0zvuwAbiY5VYI7gyb
FLtppxEYMukMqU8TEQERjoyAZTvwMyOoDZ00vuVola+8ag1A7xUjTUdDPUce9G7B5cxKWKLCGCbe
iXaHuFeq9jy6/NXx/MsZOeqRsNiFFu6dIOr0r1R8YTc+xrZU/hGOMacezohNAI0uV6lJgZma+/lf
Gt7k1nkkcMjkLCyN2svd06qM8zu5HxHhr9feVkz1rDFVQgtIaHkkRuO2EO6OLUh4jDX0gA6vSdIW
1tTig8/UxRtxn4erXhQTrGZrOrAHdUFFGubqLceQ7xPU9FP/bTt+DFY/xcXid+gJM//enbTSfehg
17Zwm/JFP4eVRyo9cu3alZI7E8p2OtQyhPuj5oAjSrZ9gPULJ/6HLs0u22uwJ5rsWU+RlGM8qnRR
ApBPTvwt6oHl6Vo4MjC+mREYUS25DJ78bK0GkhNzwppzCb8PTo2lAZbcp+TUwgf6jrJ9t00cKJvc
Y0798Bb4/HmKRGKainslfqu4QUNWvE5bwmdPrKk/WjtIursfnhYL2SflAbYAAbnpNPIaCj2/l/sO
eIx5sQki6yNgcy+PBADJZFI4wCntqR5054v6siwzPvJ6WQyqQNRqgKZwBZPR+2TeUD5gzFEfZnze
Z2CmF6rvyZ9MG4snfTXyIhYQUE3L0elGj8SCOR/A/FglqEkA3yVSmaIfPehkHgpPockuDycJ/Gk6
fWxrV/WvipygZ4RLTzVDsB3Nf4Um8gYD+TzLoKq4RypYu3vJvch8X5sB2sAO/JcbxABOVU/EprVw
t/2+0VXUUARaO+l94mCSoTmZnEbk0vNXrIVsECxhYrIUIV2ta113N2G8Ng5L9P20yfRxCO0LMhIf
5Ba0sVra0ufdsYhmSUJJwt2nnzgEcyKJkoXpPuUVOLiCK43B5Hug7KOK0/Ce/NB3NqAkecNLyzBA
+v98E/FOB6Y0Sy+hraLmGkdnKiX48XJRV1s8AB5TE8fBzxpcn/t97Oa+L1HwwBUegBqm0bzBgkkc
TItmnNiY0N/eV3UvA/Yg/UD23yqOff89wtQ087e0UyYfkBX9T+wcXH7mQ2DakVFNUnVffPW56rI7
SYCTp3/CbYnCv2+0T28CY/iTJSXHmWcnN51iWS51VS04wHYzv19mjLuHRVAAGhsbVr+j4xE1njeZ
YpD6aIHJSlz2y2qIxSa5plIch/PEgW12Um9p35eNMiijqZt2h+/lVXaTKnNivzezw7MjQckqhHkd
tDeuBDSC3PDDbYe1ohBpCihKVpSFgSQg/n9ylnWmtrksNQEgoN2z+hR2JMAhndNvK5HMX7yCclCM
Hhs4FV9rAwVlne27fJ97gQmv0UVuW0UQJhAsQ022fRoBOHaX7NrBnMLfv5kfsCPDLLDwGVgG4lgQ
C0dh4sEWXQSOkSF7tRDBzlHfLAbqniVcXlf4+v/HLddjV/zx/uzENGT4mUFyF+At15EMifJIIl+A
XUeVzip1fua+ttHXYWueVBbTTO282mr6XDDliiJORG3f9Kk+jVRTQW6MRQOTcM6xtqpxuxB5wp4Q
+v4hPIvCOff89JtFXgzjYO/LcC1T4O0qoU6PkHPVwx4qi/Z8Gj6GeXat1nrO4ZEkaDCcVdB2YiwS
CB01GJuhWYLGXB5OCsd35nwRAC/6F8uA0QdnGAu7BFgzMmzeLVqI6eYz8MiWZykA3lEUPCyK0ycw
yLProQhgSE0RVW5XFY/RP8OTgvYl0gdd5oOu77NefX5qd84gpBs+hRLPIUnPT3lhfhIRs+K3kVeO
qF1HlMp7/tXaIk2ylLf0X04DSYsVOLEmfelE4KHn1OjFbJlbtlxu7iRT3upT30DuyavionU09Sdk
u0/pIf+G73ccsoppJupz/8qcjY8Ngb5+TP/zqyQElVesXIin7xRLGYc+4l9iJmwhc3Oto4FxqIgi
7VIyXg/dwqj7/2WnWEMK/VZqxVLvf5/eJBCf1RvOD28KAwrfSe76CyzYBL4s3jmGU8xWEfUvwQM1
z8QCLeVK0lws8eAugLwFv0KtHrlwY4peA5Mm/DgmOUHya5XBzhGEXFE2Pd9tr/qXomPCgtd/Dt2+
K4UC+8Al2nG1w2CBf6d5LOzrRk6CMdLcA2lks+u8vcwjZjt834ZdPneFIokMpV+DTH0tr8VpN5R2
Rqe5TjzONOfhGoDthS+5AicNoXOaXvqvzrKJq20x8MDZ2C+3x+i4VVTAnCJBGEQwm+3bEQkdVFSm
KNHxByZJ59zrCF8oY5OYuJDalFFIeixpf2LjYLWjUFR8QwuISybi5OIKhnnZI0NesWexwAXJt10I
ktuoEhpLlI+Gq1yjLrPtI6EusQuR5IG/WH4v7/rKVmWeKfKvDewhsYLkMEPxaDPhxGNVBlhHPVfW
Kbed17+vHfB+hYc0xwbf79LvYNJWgAxO+Q16lQB6kW4ljdQDrpZG0X0pp0sE6ZR9qlaT1SH3uSBd
e1+1gCoJiO93ieEyufzjiLrasvBHdJ2CADo71mQpG2QRzpBmSQwsI9nSD1PqinXh5RQXYorF8FZI
oDWK38zPGQSYpTwVupP5pGxznZhALAvrSy6TwNFgj0Zho9nobcAZAAm06hZ+WN2ULoLN62K9DlpQ
cPgeQE2wXbs2pzwbfKHJYF+9P3q4CPzS65wQA5ubH0JkGqQH1OsKIi7d4p/BoiRPUTj2ymTk4NTE
tujrTlrBVdfhqzcwYTDVrQQ+/I7EyVrwo30N4CfELAVjlHqqi+9LOiZ//Kkduq4I+C/hR3wVemYY
XmjS9iozNyuGCwdax+gioiK1Ehl7KU/m/T2IEc/Pl6yFqYNQt4rCIDdItAjouHVKmZA7moXWnxef
hQ4C4rkLtUjZ4qOzAw6q3IaAfpI0j7JtFv6AR8ozH36lGQd3v+lqO9cCgU2CVTWnW67P6uw8dyVs
TCqByafKxHjq1d2VsLTcAQGmVTS/+ao+ZsH0/oPfip3ABOfGlKRv4I2lsIhjYVoVwOdmVLLNiklQ
h/OrXGvxavj6fV5ZDM6BEnS7q19ENJ3Z7xK5FWPKLhpzXZbmZC3Tuupbj5AkL+YaQ00prsThUZev
jRpFdduWsQypXGs8xBpooGEffUQpwzhBg8gZqmDDjcTickNl3FA5nONQdGPrPPsfWfxTv9FOJxiH
cdu7CFP7Wv8NIW/u9VG1WZA78kDT++mzoceRH7YvUJVz0VD10Ouy8+QvfdOJQdzZtPcnXdEylYx1
51vJ7xqGyEceIUBiLc4H4AZmCQoOsreE38uyxqhzN6CbjnCxfuzito91BdUDvdUCBkag3u7HzjDn
zO/ZGDUjIb87AeYctU+t5aavnAcyMHT05LASQiBygpCrnjlUNQAqatzn06rQaEpROSNQ1clYVdY9
YXO1G22baXw1SfQfv10X8jWcaWgrAPiyUZewXEh2LLG8PFdS+5SOwuTZBM22ZGFHYA/6uQSsb+G/
lmy0B9sInLefHIOPN4in1Yq4u1+6ADl3ezMy9sURToGEIhgJXmtp3KBfHSVgrY9GwdPGJPrTPdfR
cZSHHGMxbrR97x0nEeUOsKEhznU+DFIppjYv8AZCU6s3WVZQYjhevqZEljSf5BH+OvDZ3xY4FsA3
Jhc6ICUZGEmVyECKII2IWca2Sz32Ir3a1dMxU0dvO7E875HQROX/+0rOMGXesvL+K5fHHv6WjkJn
wSAqO9Kzq/YWW6WPBtARO4T1v473g/pucxOj1+SKmswpS7bjPBdzoZmtHOotK24fDgaSyM1CrkeK
ktSjJ+h2J10nzdkmgAYR8wre0AiKa/iH7Wi9nompDW2f386rPDCq2CKYet52XVmfTuCjxUdES69i
TLkX1AdcLifzPMKuNThXBnyBtIbKkAXvORCQ7Bi/5kAhgDDGeoDZjQnov5azL6wA8UwFjUBPyhHV
QTj/5c6TyYmB3OpJY0x07vDqNZWs1EetUbZl3qLhfV8N/0vx5YtakigrDi///u/p9wsP+2OsZpF5
C0VoQs9vmamQPTldk4mVCCA2uJyESLZ4oTd7z6shfceBVsC4p8SdhbQAKA2EnNyIuj4F2+uZhJWF
aJH/uD0WYrP//Sa3QNoHo9QJctvdtIB4INrhVukMhEd+hLbd0i91y3MDtEHlgxDEBEOSgDV8sKKo
GW+9w3Xnkav5hTSOuuAacB57yg1ysI8fj5gqibG96PD9hbatv5gqXncWNmRO+JMD5V+kuXUwF6Bi
W3B6oEwo7gWEPfhSfkHSHrm4Y1isNJG9LfTBBdPd1JgHqmxGul4AgJYjpEpw7OUyusdsNdz+1ENA
a0U/ERBXFHeKXrWFnBX/cpOsdJWADo72ySqGOCMueXkBs56KJtQsK0/8n1W9g0lMra0VdJDaE1vT
zSA4+LAWuz9U1WJRe4353K5OsmxqHNr3MRHpFFRDkbD7ORNdHZeNmLjZdVBAMMQseqSRXVpv3kXh
v172U3SNoMtO5a+z/VLnif6leZHpnjfhr2/2W24czYOEDK21nUUBm+CN+O+PS1RbGr1vBFOUGTXs
erSeNIjwjsyb84TTKUEPyDNy00EHx4uD1utuGepZ/I607fzXY+eqH/WptyL20scrdcua0x8hUYDU
yRJjanawTKyGzdy965N6OMVg3xqKhG5mrGGnF/IckbdotwToijLY0rWEfm5P1gbFtpot/c8+/IO+
qzf+rbPGBsgCz6NvtqHOQ7PNgXKDHucnlgEf7FpikJls2JvoFX7huPhEo9ARA64GarOBQ7P11Jih
9z94Jnsn3bzJgMtS6UrxuKHxBFzGlXGa96H310sA6kCbYgwKJ+zRK+p+L6x7UUPwUG0eZxBNaeAa
0OWqDDoDNowmQpQhy1uVk9cS8XtvEhJxO8fE5ye8LXn6Gvei/FbK7AIBkZg2AY7X2jYwkEvpf8uc
BNpkPjNzSULq2NDQy3mgvOG3uI2jIuizcOO/9aQdbWor3hu/LdQ9wKR7wYUzK4AoBhgT2jqGN86l
8+4xFg8lsEpGfqFWAMZzorKpJFHos0Uk5lqU+Nf75p0TcphFsOo3avIDPfXVv4WY1YZ0lM7YkiVw
bHtEc7BVezj7J3QX97E3qCY0cSF2+/AAtZuBn6hSPYSpGZO2uzjq8O27oAMvA0rlejNZlOJ/kACp
lQrgt56LGg/GPAnOh7qgGNxahUh29e/ZTOuCAbmmH+sabfNdS59mC+kBLZPIzxSwsV1vhjvsUpSx
ECP+6AMldxmlPYLOG/hDWTH+cw3CWOWHqjutYiZDeI14TUxSHHGMmi65APDyovuJsnUvMjVsVFow
0UWcbUFlYnCFbBDNfW6Zfs7eLIIRHjWKRwYv8JB/ZIpdUQUIoFJk5G647FdqKbBJ5dBQkx+LS/+q
9/c6f/zdDAxe4oMHe/aL6r4YB2iiZfFNsJnc3N9C6nqLlfU3sRojkpC+8tHhw97iew6CNG8S+LLN
kkYhcAekF9MyhV0cMNyF51uvKYQSIcLRERzzu5cQBgVY10cKJDIfAdQlEu1maxOPjsEd3Q37WLUw
R6iAb9B8rMBCBzgFGjm8SIzCRr95NBROy7q5ChIV7daM/RP5LLrU8iLoGyqton5F9wrbbeDOn/39
yLyPXq0PzuslfrBddHnF+OUqY5z9dkSBCx5MliFWRf53D74FbO1elbin/tB+/QH5JJPAqxTgdduV
ir91JqJO+hEikQd+4ql4odyHYy+o+0WFb7LCCEd4JgA8wjHhvDUajVD0ze1njiYgt+NF0cO79boY
b+zhuMtpVdwUUqww4tqoMFPZLaseA4YiZu2jVphX3vhagApEE3ddrHCkJmp2BjxuccF3IbT8Tqv0
lwjldDsvk/u05INEbWEWRCF9Za4fjMS3pmgSRmg16p3qJnj1yuLBu6FZifjtORexuUBzhFJXg/o6
pUKfnreg6rNn+amvW7vRi4KJdW8RvSImyc/aD4pB6SnAlm6TK4XD6pt5hkg73beq2AWoetZhASno
wBCpmxNPVZvHMfLLn3Lzg9jGwBqQ39+Lox5NKiCTcJMg3+xo2PscJB4wphsqXydQgc6FVRXLGFX8
HEFapze1C00MkyogbEmfsBiV45VbbC+DnI8BJS7CPPI6f/pnq9ctSzAhKuGQV/Fx4iCJx2NFw2nn
p3EQ4iduUC2lsjZPS85EqwGUQPwFiDAzcbViAz1Sxw4d54iD/pa1cQ83nwP1vAzS5axASIZelSVD
54Jm3iGAzXVz/uFR6FVijqwOQB8YByYSHqrhZJOKCzgLjc9Zk1K9MBlNIOY/goLP/ZFjSDbAAT4D
8ARVkBG7/2w7yIC9wdrBF1ld/blKDy/iHBS4TcPjqjM3kJSOsdIPCIwzHUL2XpaPgimP8yuSWQDD
VqdSkT7LuxwMDZmaliOTxCcmpWf/MDrp1M9PRfr1cTM63ag72WYlZ2l4x1DMtPYJRSdnQYAmggB0
kXMQgiaIqu1CaSbhkV3FfwGsrrd3+pfT6Jwo16FIQOtEYhAAyz7eNDXi4EXUfXxfbBKrtuTYyyna
zI3eMTLNftEd1zQRbf5YIpwE1FgaMfiRaKXCdsv41OlXWs/7ospKl8j36w1XgtjcjDST0KL5W+B7
r/jI3Rpfwg872zFnPut+bkP5qvsKLej8CEfR/qsbG91qZGJHipBsYIEeEnt+ztEXn3IYgebegx0o
9M0l3eawdnJyeQ0tczXsnNZAFD6tP/jG/PfcVeyT2P2l6KBGW3O3G2gUAD1jIsPoyPBKWkv6XLqc
ekkRKN3HEMdhUzj6pm98pS3lrpmd2EnJFHsPxr05CVdicLx1Xtz4Y1fYcz7LiRCkquvsd+4xzGcF
LI//GP/2yVThpf4FKAVw3fW0RfurW85sKT4RKDlFU7nJ6Ibd41nBoqjFCrW+M+cairpsbCjROMx0
yfX4TNu0PXQytLAv3RqZXbZTLKkKH7YS2+Uiqoq3uv889rh4+pb0UDPxkMmU70xnh3HPKF7/ywuc
KZhE81IgVc8IW2Y7Q9S4iahBky4Anq5pv0ycFyzBxccZ3qeZgdDM7nbCQx8Et+0MHbJU5VXxo1ZE
iUJDefLOtHUwEuVHpzxACMT1xSNKaWZyoh7B6q9bjt94o/M33y1oB/pq6O/2S+RWB64omA/qRWuD
zpgsK0uGe2a20AZlNTlh/60b8cVv0n19a8CrQ2IQ7r45PH5axSH2g8GvVRFIfCU9fg3Fv2NdeKa3
3rWULGeC2WtRlSFs61JfyPS9+lhvPoOLSJ2cpiVft9qN/DulwKuM55dQEzZrMHhupnZ3HAkOxzA0
3htdTXI9OXl0pGtCcZ9Cppg+wh/xmk8o8s7tWFerdrloTV+ef9P9B7URD9uNuRC7Pc/QGvuXiEUA
B3Mf/keta6LPoVNSRsnyYTwn3i/BnM2NXT5/oedG2et2g6PoGxwwGJUgj6gCmun/v7Z526G+vYCj
neNQ1sm/lS9S43UT5Nsmh+dgsJhwc1OjxkFvHANCi/5DjuvVx+1N8zMSRBz5ud7Hw6Acbg2nqkvp
XR8MVuUbcTsdLmnv8FpvQlYpg/7p1VAobNYCLdBGoF2dxAkVKC11+/s2qeQEFtetL8tLMAWccL1X
VrWZpd7DdRuvBRpDk38sHey3kNVwhU9snWUa//miOJg2ywnqBenpjIdxfeMBdIRmAXjE13lORepl
41WvAyZ4h0dzVVtphGityRQzQKpEGf+WAZ8dF8zpO0MHYkR2Xq2Gf9Jx6Iz04vk/OzqGJAZqXs+C
gNh45qVeVdZQpmeOn0LBWYD/5UdZZkxVr2ao/blao2/UCiGqaqVmSCpnsyrjIpnnT/7mJjXLwWWW
fg0I8S7GO2gWX9Wm/mvQygZCyBeIRmC9cA5taraBTUMfwSG8c9yOY0m/TbTibdaZUNJ6qbnTJUgD
ymhEg7fGRn1yON2lkXhKh86iyqtANcYZBI6rRMR+wFvviIkZEXvpEh+GS12S11ASnINhRqVGHDf3
d5Ud906W6gsOQQ80AB0YXnMcsYOwQqvMMBQqtisHnNp2oDTYBo1B54whMNknis51uETkuvaKhfmw
5QnAybgNf9xRVbEdN4DDLql5dq9pa3VIfJPMvXRKZ5U5uq0HBGd5rFQ7ylt/bIu6TRqLOMV3f5qm
2Gznm7foy/rUI8rFH9nUwD0nhuUeAvWjdFu8TmijfVNcWgZmrVAlDEOltmm/vbtx3Qh49r229mh7
WDUWADt1Luo2oAlEWz0W8iRBTXBU9C3d1fV+7Hu0Oh1Vr+Z1pw/XoHvx2l63LtU78B4RwQrLV00l
kRK7QmEywsP0BvJ5WYhZQ2ZynIZQDKZY4BX0djkKoRu9jqlZY1acj4JjhHxdEmW+sw6RKkpMmSN0
qZ+gmk6NC9GRneN9ce/UvM6dHxcqFIs9kn/yYeVwJ2gIYShNtECOSOt4jTwhsx1CIm6Vr9+zjMA7
0IyOSf+0XYJ2VnBpgWNpO+9m17Dc15tLn8Dc9L670xjNERfyi3Mgy5Kjbys5VtP4al30bfTP4MMA
qQowLwrBhejnCDhDjcgoCiwFoo4srrt5uLxQF2cRJQZkJHAH4gDIqRJnZ/YqEsGpPB/muyE4JCpZ
PUI4dcuTdlK0zNKLWHu9POphiBnSE1GASbRodCSCAI38AcEnVa3fGZoV6np1OVOI5IkNq+nhW9Rv
gt9NkMDClrBposwWib+tlMezU2n+1H9nHx6DKrR4hOfrjkUGK45YdvEwTEtUTC7WN8mGMnj+k8n2
4ykWlasnnWEF25sVxofOCGM9nGylkGe4FMrxWHtljjfeLvKLYr1Ses3LUo2Q0fW9gido2gEccuWE
rhInWUx6/UZ7u7eoVCr/og0ADrdJzxwTHvDW6VJQdJXt7aS3IsT8eY0RhIgMS7i5B9bvqr34p1+H
m4YYJKZ0zJ2o1MuXfETFHIg2G8fkfE9KEHMk/w4pEFmp+IV6CZprTYW8FgtEUH8YWrpDqfetmApu
JnrIapj7n+MPdpsFlQ/4cWmztIaNxO84sBmF8rRLsX+nuuKmqROObxbiqddKCMwU4ClIMcO1OUoE
SLMXUthzv2swCgICh3HbUbWgdwy7XkV3Ee2qkY1wB9FpUCACtM0PsAN/KwZ/kFY4USMTQjmDKH8p
cVi9NxhpokXRHdan6LY29migmc+rSPwRT2yW4RchTqyqkqeAEwOJ/Jg7AH36id2UrQoXsxfwSxlR
ZwOoQdmKxBQ5O3ap+f3Kj2jtYLZfL/FCe9qSKNd3/O5IN4gAp0nYpgQJlwYo+H4FyL3xVlSdwc12
TyjlHcDQxnqxBZ8m20y2hGcRnkkMIcKY655hEQ8RKbygujzHAv4OrIFl7860BCeCwR81oMTF7wBF
NTK4bz5U0PUKBK/vUUi30UZTwWp2Ulw45ikSIZTRLPEtIrlBYT4GYgLOXf16t6WjX44JW64bgRjR
lhUVQiiS0uZ974ePGFBOaoZ+aPoiAVphSXGa0SPGhSQov/PCFiGoN7ofmNjE4zp65cZyGBerqek7
RnJiFP6b7GhG5PDW3Wnha5A8c1W9NYz0fIYWYRcYAOfyq/UQkpGAA9MOwHgf3xO7MCLWHZTXKnus
vg9oUeAvo98zX9VQ3BPxrKhkrDHHCSuL2ipenQIAeM7U4rcDTlE5I7FSDXSU/24ZVqrQYX5/TAxa
76kQdoqdmKsS2XHv+G4tWbILno9a+2MUNmUFPF6NQJmy0cfUxCGjQSsDRqJti10yZEgQVuXbg0e2
GM/9ulv4KIyTxikO2X06yaSFPySWKi8vJ8Yuqloq/it4f865oIopbAuiheSfzy72OJDGgPVSogJf
dzQC3PpdyYJu31l0YNR4CnpSu+K2aoQekvwi0ABL9LT5g3L8u3kPiEJhjobWsC0kurFQydoYhv7q
3OAEtQ2N359M27NhsBsYEDbMDlYPt3U6q5D3IWvs3TFhvJJyHnGRzwSF2PnchB0xRsuL1SA7ZLON
9l7WXhHSKbGLRaf7/0+42ha4+UewjnnNUhBefKwaifzGpKq2JeviLuHNTlItjXV2NmpQwN2gtvao
lNzT3JEi2gbqNtVKYzLHAxqk+qfABkx0HivdYcrwUh04fMXQteL56RiyKfxSLDWDDOnTOLWHXQGp
/NSHJSuRsJD9LLhY53wFQeks0tNkc2lw/L22G6+nshfMkQO2sCX4+6EmB8/HlZiel9Zn9ccRfSIk
LUgoMG5gQdbRlpHIwcuNJRsCZmNVdFLIXORb2eKz3jdzvGRAf2VibLpgoUVMQM5MnbYuHZMKmC3z
h2f51vTHeRprutJuw18gvEs7LwhzORF0p6gtzsq6Hj2nau3FTO4pclZDK1fOG0zjX/fbk7WWJdcF
wApfUMth8M+gq/EGNgMQrARZ11cxNvhHFDp40gBSR7uJMIIxhifwZbZpZ2vnH47d+JEzdPrV0qg4
9hoPXuESpRecw1mxspGXhBW+6WjzlCVQuErJu0viNdFpznzbwCnzfi4Qv6YetYWpAUIMUmSPCHxP
BAJExTT1aiTQqh+Zw3mCJtOT8YOUqdka5IwzsmbRiK/XSIxpLGc6vgkA0rabfeyIIfjhSXQlZqiu
ZoWrfo+PYVw5rN/1ZxNDACkfhmS9P9WXKLWzMTHR6pKO1ezwj2InxgAObIm3JbXN0R/p4vg/sT5Q
kaLitAt3AwmmIqfhK6a83dOCPsj1TiWQvPXnmRQK04ryAUUGUQ+sVlfihzOGdU5n0fULgePVVaaY
bwUU94TChOip0PdXCtevpgRumq1t3RIKFbV2Yq3H6KQiGJM4b3W1HR1cRc0F/ddkTBBhEkDgofBL
8kUgOC293yCCadLozn8BIp2ocu8NVTEOhJE0jSfZ10cBsd4fUH8H9wCYTNXT4aKrbloZaS6wb+LO
cbyhux05K8/O8QVsb92a+5DmYELt/H5F7jTwBJKlxn4x9601tFatoQwKr5VkiPuMr3drW/nlZiyr
Gjy4SuikNmKNf7qsEo1lkIt73Eebo2D81sEwm5GnT/fmGHYkWKgdz3nKoWmWw4fQphDe0LmiHJow
M3R5hYyfuKBUSsBunY0XbHta/nGkyhre4CbVzb2J6cfn1w4O29HCoFK2p+M3pnssUMkjoImsHqdr
URPilhfVQCAp10t7+DaVf6kKsSlX/8DA3qtf0p1/B3hKIjocII4J49DMHk+Xs7fha5UdZZs14fiW
Oypf81ujdyoqmEwOLshWu+EzBlBgML7BBAT479DcOAXt3LK5eJOFf2EgHGIo2MTD8t9H5233kWwY
1AqYYkLdyzewII9+xwwsazyikGHp0T1F2zDNKpLvXpu4BoYTIUVlyVWN/Pz1UPpCv7zWajkxs9Ln
n11oZZKBmVsb0Y8POCaZ3d5kZFEeXatD00Wo6ME1k23W/ER8yNdR3iCRN/GVw2oq0cIKCVSYYykR
3E8nVlNItn78rnOVIAqxEzBlVyLGyt12kZ3Db+crHoI8IImviCu60qYfb7jYK37Vl/VYZXiMLcw7
a2OQ/ExS0EGjy8ASvj2yXh7OuZI/oAQ5cQNXCblmX7/sMvb7GbubuVxQdnn590/4OxD3i58P7olG
Q1kbNvqawm5MmJA4MVYH/tCAfFHaxXQluhOJyqKuaJ6yziElep+r985naWo+1sKMQd+Alocc/dvE
oK+g/jlrkYp7Q4+RcYOluVLB4CXqEOk5hwdsidYmW0HvpAl0X8yrFY9uZOX7iYqHetaZ9tg5zmXT
pfSTwooLcViIaEsYUFZNsMBiAyMe8INt753Aq8f2m9pxt+QPRkGq7aVHICR8heBo28nZ59tz1qF5
EeHPZWrcn6TYxbq/QZHVkATWy1Gc11WnBpg8PViHnu8L2lB3kr9P0YBuCZPBNnCimKwsxLzCwDvm
yLAtF+lRT0N4k2l+vIEV7P+k7wPU2XERDnSKNwlc7T1QofZr+rVrBIvN/au67UTipqW9e+TZb3tl
WPuCsWYKApZwormTHbtlnvzpCOMn90oshxeUrESQZrGcja/idVMfbpcwaPPUqqQLmabC+9FUSXTS
3OTL+/8gBmygPyNIqjyovAuy//RWpBP2y4K5z9jYW4tt6tf1weNrgrLLlldryIkUQregEgyKDweY
F+ubMX+RenmI5iZue4qe8HskVStBqMzIy/2s5CsfeGIwHlHFATgj0jyHNNeFZhcPx9tGAFQ8VG22
APMwAfNcP7+sw5iv8h0+Y6OlgYEcMdGx6vYcAHQTIVCBORMFWrmwx744JySIHilhNssXp0veXnuN
6ENwxjt6VIOr/Dvg0FrJQ579Hx4qGTDSKcMcLZubXLsd5boi+KrXIBm5n5jDlLSAnGl3+W4OHyHf
c9ZpjjuUPH5fdyLr5kATYRyV1lgn401DQoj6hcP9Z2KjVOn/tIwIms9EdhXzvDwaETEQAHtfUqJM
SP/4YCQaDJRpAJH1Hd1DnQoH/PygsVBghHGEBHROX+JyOvOBvuoTo8mjXyNQlXTo1IBPGY2BagTt
38MPEk7ASCYT/MtnDkfCqJrmoKQqaJl0NIJIfy/q+dq6/N555lZeyMd38od1gfXvoVhDvavl2jVT
reWxszRHxQhSej/NpFfWDB5+i7PZRzdeKCXCzJd16nuOCMoUKRhBfdXMYAFBGUp932qD38DMgky6
ip1W4DuHFxr9WMe2MjtZJ7yZwzE+1kdA+4wWYeyJE7gfFhAjKCRFNaL68g4G+FZR81NB64has0gJ
x6v7ym7aoidJ6HbvBO4Oh2hDtQTu1j6qoEopORVYnddtu3YeYRZh/suZu0Hy6VpI780rrkHQvb5j
Vlsh4gKY8NkRyPSRIBA0s+Msma/Km/jUI2g2CwqGb6/xYdfcMm+DPRIAdMWjj+8gxPke5/pMHmxj
YbgQm4Fto095WW60jjpF+zvea1+CmkJKbLIcP36DTTpslZiqykh0WRkW+1NUn3WUMB1/3tibq8i1
TsmgBu2a8P7SlzB0d9kVn9OevdA9xxWqZ7dV00O0mbVkUBOhiy/Pw6jGKRItyz/fG9zdnYvgB/l2
ZpvHNamVEEbPLCA9KJkF1upKuydK7NiRecP4SureLJVjzy9VzigoAQ/0rcj1jySOMy1Si/nfwCbO
RRkZlYl8QywWVxFWYRT+U/BwpPAdCCUZonFDcUBm0tUPr4OYlxb4HL7/ZgWq78grZRfDendlKEV/
d66dW/K9qUUVlqUhHtMDmer/Pi4xAWa+39Rbh5lkPF3+1UQXSAO80gqeuAb1h2Plz+YFqgzhVL1+
rstxqFMJcKrwgdYXOxoa6uMbk1LFBfIXr/hz4aqKEOUS5h2dRMhv/k2F/LssdiMDcLAUATCmTpmC
+OZkmaVzMFMwAYu71Dka8B7WlO86QjOKGgdl0xp5lVFXh0Jza0zbhmoAXfB0TEMmN8hEkeWoo+bz
WsSjQ+FV4UFaJlijdvkz5+PWLXxHNcYLXLZBj3cNE+/JK7qiVLn2gkt2UjXvl/1RfC6/8V/VPeJU
o0rB/DbtyDB3sAyZGjF/PAsAhiMbWK4WVdeUdnr6H+ESZ2sQtKsor5WtAahMQRXbRN+dDGfR5PIF
RM1Y7O4vKNAoq6nZmv3eThult62bkgTk9ghn4vSgyxZnhgRvYbmnOmS4YjmC2rypTGBRZkus16CS
DspMMdEqWMgaLH/DGfAuXHJjrtJ6xevM/Ijo+XG0yPpfkGFUGZGB+zFfeKnW7JtYMtwrXP5Om6LO
XXHT/N9Xva/QF1PDQTAZt7tS7CwNO+7s98ZwlKrd2z3BQAtBq2K7DbRXTdUy1CEegJ7T3c8ft3lp
F8q5Jaiwk/j5MGOrxfNvk3+Wi6rxSzx7KTRwlW8KGaZXBnxRoF9j5ZyCq+GaBHtjShKx2kGY0Cvl
niTUtIDMxDpBaR73YJQOqjxDpW3NT9ujHvdcTqaOCqrdH0Y/Y/FtpAIdMwnWiX3HxwkQPxbLHfaq
bxXQTYPul9KYnkc1av0z3CDoy80xUS9c6wDGHMIeMLag+Zf5S+cM0ESxIULMHcGAq0kLNPZs/2Vf
WuIseqpsAJgJI8TsZi/tB/5gZkHASC9oJUCBnjSAKGYcHFXn3Q/GN9r6BIhEJNaumbdas+ITx/g6
pbL1CxOuXkQsAgYByvzM+jjNFBO3fnTi8Hzdyf+t45UdCaOJZtXJykh1DtkAC4IQLX+7ozt9iueB
3T5S8RyBJjlDdUsNJy/yETM5bl4jrMWPb3DUrlxmKMfUPRwL10Tasz+//2BVtQmGGxvag32SamoM
AlzPum6Sf5owd/anvj0dBec/XXLTeBVatEDEkb924tn1k/IINI7j5tHJacTdRx/zx19uJ+65KpT6
kObPezAwHNm3xwI9wT559hO+ymUEo34Ep5ln4GTTEq8ZNP7RBSEPkYDl1cT6W7GyB/W3jzybNaSw
v6WUtofd7NfjIn7pDST7QXMZ3P+JXHRr81VzMkRS9Dce3mUikidJQpm4GzTMIw9G+1lAPTOv1Eai
8ElOdzzbwwNyrqFbZ5MayWpZHQf3AuTAj59iEa6+Ud6EVd4QLo81LqRyezdhSxx82AeL4IgFBdva
iAnfcJ4V0Ita6VJd/B8g5q252VCLCrCj74OxsLQLC6PJa+t/Crh9TOq2IP5muIWdyPB1V09acDec
Oi+DMYzM43UWQjyzfVEUBse+Nhoa9gK1wOLjTKybOlo77PUlJiovxcINx5e5bkEXnvQ0PX1PkzGA
/MVv8EZCCCKBsQ/43V0TdvZUMEzf6i4cqBT0sqZd+uMv+mKzLsVJe3h0/BBdLfTwHF7etF4tSAYi
JQQ2jw3k4UNFHrkKF/pyGUwzqZaYJHNqpQ2lgiIqATP16yZ7tsEjuB/yGtvBeDROR/AYLkW5CjT4
ekHoyEjzrARVWaFLms3TzgAxndQqBPJN2KebvOPK9SVM5o1Jn7RdyJrn+96H9Pj8TigqBEERbvMB
y9tz/E2yMQCDgo/+kW8kqleW4cbGs9isgG+l1cpGqwarS1jRyLdSsXsW+jFGcdfIeFyi+cFdCVjn
oUduf27/WjE6N/xEXBuWEvF63NXrcm9ZbetWtGzsvtUK5mwfu01i2LvNPKejyX0xa17bGmBCJ/h7
LGVtDvAsTZPXyTomNoatJD2H0eMoa8hCBdUQZEWeQAW2AZJ1IYQIXiqRRAyZMj3zwVoaXc+x5rWx
8hEHr1Q0m50uKsW5ZB4ASD1RXkE6acHEb7Ri/4TkfQeyGbtIIXiZnV1pfufjBwq7KUtfWhK5rspt
QsxH/P2yEyv4tlF3/NGKZBh2Sa1d2SI6zL42CPXbF4aMlsHKCUqbugV7ImqCUaoBAuxNAg7drz3p
BcidiTSiBLvm/tH/bBECcRzy8D/CBLXp7BCE65LTVzK8Gy5eM0J+Qny0fPG9rZzk83vokHyIbY23
hVu7PrS8ABHN/QMfW3bU61aIsnEdVceCyBNo/x88XdId/1/CdiBzXhJ2m+fraDZ0Ptdal1k21++s
+3bOViHn3dgB8ZP4JUUyQM5jZA7Lh/PnlMe+fci0AINyKR4etDsgDB311PDk2k2B7/l6V7nefqwR
FMVUMxDYqbrkC6X3t+NY97CP44b7NMgVRBkjKeiiQ9lPn6bJr+2mVNI4bNqqzUsElCc9Uaxn/KJ8
rVnDRnWMD5bwZDJnvXG8cnm3yBXRffdNfcZUqocEMK7puCWqrJ2SQRghbjIGjn22dw7iWY9PfkMY
RLmU2Mdgy+LPU4i+SdQg62VHTC/2U9VHDG5YUf7FA3QJh2sq9vG++JU3n9F6oGE/FNnsuCE9RMke
aP32PHFT7bk4VieIejf6SnRSjaxC11WQwGJ8xfKnUZtowqoSxiG8rUUS61ld/jQIhEOo8FHz/Bcp
Rlbi5hznp/rcCnB1RCF6jWkQdpFmGqFDiN3+xffsXEa+L/VuOkEXQDiiknL8Rm7L8tO8W3w0P4SO
cIziaVCYxWOtbp8g1UfRy+u4WP1lSuVIz1v8zIQuNhH5gpDy22cyv5KvNEP8DxyxT+E6lNFLJtOz
2xor8jeInYVYCFZULUNgQI5o0HImWE6NC8hzP9viacjTv2FkV4qFwmMfm0lgE2jYxX8tDPg20Qu1
lKyQI7z2lC/T2YzUoBsqEad9aUJjVCsVItcrF8fTqU1PcnifXWDiY/3KVKYW08qhsKGk9iln5Bko
TWEuDoPpUiIbq2FHh7V3d3a9TZZcN2CRC31anPtFXrM9gH1awzKabOHgiDgCBBMH2pUyL5pPcl3u
zHV0tqoKXSM5WAy9Oa+Zn1c2LRs3MgAgwxIFoebloxzHdRlKpWfXbEKLL6Pv42bmzTlAOb+LXJya
6IcEtrCzZuhGrw+CaXQ72u0Tl/MFvAL9V5wTfop2YQ2uVQd9wnOsWIoAchPPi0DVJuMehluei/a4
GTxiWjt55TCDWGArBhRBZr5ErckySgvDXdGZOXPJdueJh/24LsJnW76qc2LhHEojqxDFlABS0VXE
lJfP010bA+NDbzHCL4vGzblxYsLM8TqeQXIVx6BU/AbRaKmSsrDxPgxcItdLEzTxhs8sCoj4dGq/
zAlf7hgoMM8M4B0BVQoSDetzXD0wFBbyFi4kz0hfkiu2fyP7SPgpn+gM8+d3Zsrul15SoSZkbMGJ
G/sPxPLu0JPT4/SbYATzvLOa82CzOREAvrYesFyxK1IPnbnbbcy37u49avUfdo73XIeIeA+N+dQ2
hytsFhSoKOsWewHFcpKPlU3h5Jd4xlxjhoB7+4GjsPD4pOF2uGvJSgCRPBsZ3qd1cjmc/mcXE9gv
S94e25enCVZ4eVGceWPdQ1N3ha0RJLWrl1jmDp6GkYYZtr9v+jA4XcjHnVAASaeJlAswwjUmtHap
93gu3vRLPIUZjrxte+QYtfw3R+qaDH7YsrwenIL7+GrL9kuzzVwrIJfAzhRzY3UdEgXsGAY8sabq
w/0bdx6yallMrBiI3Ho6m+KlMwkVz1rUjElw9OyIRzhgoSEXHBKEPCNTudx9ojlKiEPZjKlSs0CX
688ArPQrYaXq5F7GJ3qJ3uVDMNgUsCzEeQAybrXpsiy/jL4tqRouX+N5zcJNzNHjIZcRHD7bVIru
qBCGbtcOgnwXL4TZ0xx8Qj9unUIfJC8vNkDHkfxN3gxnYwHfty8JfeCpWnbgqS3BZbnrwUQzTRiQ
1NvsYzEc34skMWztvDZbS2X2e1sd7YDrDWB3t1etTcawbLk4L/FNosliGsvF/Q2QEhTNlF4AyShD
5cNudRCBRtDQ/7oScf+EfBGUMxwRSt7dh2pqnvLi+3mKSbSEIW+NSsSBVgIyOGthmKf8vU1dw2yh
g3fnHmRNLwv2bmJmlgw/pCKxnb9EIz8msvbpD1LX7uHxvicM7IVa2OU/MUjlDbEwAQE43q4jZINT
dxGqUK1jwRtOMQA1IsGONHQ0eoPYsx85xEmmJpPR3rBWdeoNYyIMeBv9A5HjBRFzITg74/Vru/35
9+TLHVq7mer3SQNkc2MWHhadDGsqankQtPUHqg4aX8C2tWhOvHlCp3Xp617GdsgfBeLWIrEonxcF
4chtleUzQuI9QePsls+/d5jH3fsSpupBAexCcP6pil51j16phPqEe9bFnMUbe1jgSVuZQvXvMcrN
12/eSA7P5CcVjRMc05dE1Y/yB1AfZtl2op0a5S9ZvduJE6Vo+8eyvnwOS7K4CgSgVbwwEVZMZayl
ju4snOHux9SawAAT653z36b9WuKJsuHzz+2mxVhTxE/ANSi9a997flsFtTNJ4XlTSQ4kG254BdHU
q8w383UwTbFre1c2ZQ0Ivw8FjPIdwOtNQF1G/vFh22zUMUantsnN9/181Bg9BG+2dq7CgjJ4GBlx
ApGMG0NVoYHeoM37BZgQF/eHsoZuphBaTnCuvC7rhzrY6ahdWD59M9TaHTYkyNqQhEyVEhzhpbQ7
AIAg2tluRdo23cdtlDC0LgFBni5JFv8jxzxO+OY/9F1VyTn/M2Wd+Z5mPAV0t6SN4SEjSxcrkIh6
4jeeFUcBwH8O5hb8FDgciJimBXWlvRjhBfTcP0cAnRT+XlaqrdP9J3A5yDW/38D+RQhTH3S/IsSw
fnhceTcj50pVN+20KqhPvTY39eTudyIES66Sfrf8ytrnzJzmVbvUTEXiV01SacNazUdhQfDidklI
UdQ/VSN8xIRH6RXqq113eNL2BP84ag8J8mJ/onqVqm1nqXm7LomWUnnEkqLyV+qx+Vxy6zaMe2Sy
s/UkuyzE5FuDE9Q8fe1Y8boAxSOnsO88wRCHFQfuQVoUMmMPQln89anE7S8Ujyli7SLUG3OxTuRb
xVtdbwULIMMl3BeuhNA/a395cTEohJLBONXdFS0g7KnPOZk8TNPHhNV96t5OxXC7dSx9CY50Ad7t
C38NvEiE0xZHu2Qv4puBr4wfonVew6sPwcEzRGYq13KSfRBIujRP8JOOtjnbmSnfYbIffEJiGiG8
k9rA117VOTKgRZhrTtElp4wFNwPMmQIp4eQ9jjFA8FgvJDcP/x9CdIrKFdS15raAqtm/vCfIxU/s
4BXPLAnwoVXtkZdTBmzi7kIImcmNKqJS2aAXfLu5IKxZVTXWFqMwFE53uaQM9vTAmaYBK+UCyhLd
uAx4ESPOcWgEB33vioMBKrsWRH+HKH8MiLQKAFuTGEA2odRb1VZKi9lvu5nFppYIlcFXclRZ54qk
Q3cJddRVg5Yes7zsovWXOrwaQlV8WqS8/6NbV66wG+2viQc51SxMNo6gEGXZKceW7nvcUSMXv55y
tK+i1Amtfdy/rR0k0prIoeSRVLp0UeGAY8fiMV2MpRDk5XjPOXWjBKmQwEBvggf2ey5i1BbdJFPP
m7NTzBfQmaPujM8UOCplqI8/GVVZRF+bFuV4UPrwtOLV43TbxhtsKvDwfpYtXx+dkii7XoszY2RQ
48+ganNMcNIudmE308YC6uT9aMSG+qpXRr1+qise9n04zrdK1De+JjfHmfeKHSpFTs7iNls9Json
RtBzciNGNPz8oVCgdDWb41IVnbykXD7UAmcrtaZi1j0f6u/FsdCYGBYBOiks1skHyDTxM3fAuAvc
Bomod+JDlaYY/d6+P9jd/jNEJJVwIP9Ca04gN5VAIfpxSacrx8DenRiFdbRn22DtfYH7diOgeanv
vRmwCN6k6zPeYkUBaoXUhSIGnPS2BCtogejhvBH1AfJykxgR/09RTZqwZSJbuIxyPqUipnM8l+1q
Sifbdit7F+6PZc68STsGE8oLp7Em+AlQ2Y542r1pIQZSTLHu+j9xrCpNf1/xE6wsiDTHRM8ARdJr
zz0bxh2W5kwXsjSjPn8uMMNWVktEV4sVMGX7y0LsjsdO134fpEx6/tYzF6z5awCbNloiRUbzSaKw
tOpEFKbHFOvLsCrmwRs6/ghuKf76jaQp4TVNDHPlH8wG4M8m+247MCF3F4dFE2k9+cgAufDG2lKj
AJ/ae2gaV+Bq9HLp8Ijbf5FhhJ731sISpwLAj8tyBiK3Q1Sz7Gsc9MUGbIzt0Y49isYD115B9jcl
qQpNh30NfzMD0Jyp7sjTMtyryZjTaQR9IBVSvOlJ57e0KHD//AMgkhta4Yvnjf/vX2xnj6YUedV+
0PTwG1DYc7mONFc7iMB5YpsBsu/H0dvpsGOboNkGH/hRsYRpktwYEDJ4ObLnoPETqB0MYzMToW/o
L0mqb5f4P6nuSYCOWGgYw7p5+EbgrWHTElOklGrGw3es26wN0Z6X8Wht4Vl8T8ObQ0g60Cadr4xH
SarfVAhIRtVrPd/5ygQv/OILmkodjOiA9RIhMWuJXG5bckZyuf5bQOtexgUSKq/7jjPtOsdQtU8l
/ZFwAMlk1WdZm31W2iO3PkLQn72xhDp9wxkpQGzME2oE6UFttFDCkbPoGwc1EUt/TKgXaDbrvtJ0
Ue0c/54kUYoIwAO41qNKoXY3hsmP/T0H4XYRDmNU/A6Aq9fWUsIlIdFQt2mMckbxrNeoPcTsZtEi
asvjul//Ll9W0aoGRgrmXWlVD+AVNS/slqSYDvZqzM2XeYnpVL9pv9ZJOIf7kN3A+deMBTqkHD6I
vIWG5Ub4C0ZTe3ftBRYFigGBohAmDQTF8h9Zxa+n20eBbA4R4pq8Pa6gKNqQCvuzs7BWaUSkwBbQ
2Sx6HjnoA1r152hFEEt566fNQaY/Cx2rPSvTqNZrqgW+rMqiE0RAH1RP2uVHigo5Zq/swWFYnEEs
gwgXTQ+3G/XEb9E5M1Sf7CnV5TZSb80/JNWzHhqXQIcoNLicc4/6Nawhudw890yVkrF0mdWC8K/b
fscaJOL77WlzFkVIp6TKvw2L5O5iu7L+nrDUvEkeGngVizvKDmYXokYJx4lv0sm4nwfrfhVQPzUb
LNp/TU7Jyx9ew7KvnScf/4Wu85OkW4k8H05bgRL7stoFVY+V+nI8vaz1qaQMyTm/3K/Ni42mTiyf
k39asmFcTUvDbdbDPozGFU/WHnW1DqJYeQKIoh7Yi6Smuc/+tmvjyXmOItATL6HFNcqbSdRDjjMl
wNqXgTDVy7xcZd86xsnNTR7VlFYQmNqISRaLXUTqQ6udpVMfBKRcc2gI0nEgLCzRFnS/XRP7Nr7+
wTySlKTY+A6n2r9Xrpd3H4AJBiySSZ4B7dpHp1gVsAzr5sZsdx3oBhTdlmlc82n3FqPKeHjBE7Wr
XNUnKvyaUcvd1CoHNV2q4NiZ8KfuXtjPf1if2VB6wBN7ImrRmXcIZI7m/TiOTcki8p70lcL7bqt0
Lx7E/be73lvdS5u7Q67YptBRIE+HaLe3fiH5iKKm7MYeOziFQhhDuhw5I3xi8K+Mvz9BhOfj6H/C
zjaFGPyQnmj1vKLQTwfkgLYZsfg+7zubU+2eRnlmUmRtVPKBcaSxl+0FU1U1qVL1Laj/6HcGpmLO
gR8n/PWblJYR3q/1u3k6Px0w0c9LpPMSy7EOHYUtOHoiIQ/Z40kvHx34Z7sHAuchopMurob9sTSe
PcH2KXqTinBOH0Mr7YHre6UCwJ9Xie2jUxpJJ4ZXVzgzoNGRIebb8hZ21w93A4Qk6crP1E60AtFR
XFlAkzvmR5sW439TdwPkpDHh8hLqCvEZRSOwZelzWZuXER8/7NyASCL7btagy1+UgAnQ9C8u12Ns
1kA8UJ+QNeyqLYZkLm62ZNJiap51EGlH3WKLmJoSjDMD0zXhNG9kvY+haHBKcu/nE7bAa5hLA1S0
7Tvu8Y7T9U6RcklckjRAXjyNPUGEgogAIM59EmUDmCtupsdxNcPZ9t92SZ6snW5CrsuDF/mEM9Ym
522nDspUUJjZLSI2WqN35ciZTlwaO7i3o8frwk49FRtlDT41Y8VBdb5k2MXwrRNj8HtyPlLjxrvE
wOyR3uAzK4tvfr2LLCaddfUIS4ySZfPjBGMhDoF2bYZsJpd1a1JqDmn3DU6D7wdyTcl7//gn0ary
HkK85Hh3454Bjovjvj0+Y08pkzX2YIjWzlRmLjbzjnrIuEFypKF856IZWU4owXZEBkwiioNtqgNw
6raJqQ3FdbPupVBbRUJ9G/4zpG8vIizt2Zb6JekEdGOCOEFJeyythpwbitWqaMvEexGEZ8teQwJm
Zc1/bDwh7dhEbz2RGucwZl02J7ftlRWVZHGgVyTs6aqRiid8BUJSTrnlbumM/vYEp1yVmzYrcAGL
Sx6oKaXQhGZlUzg/mlPJD8Lun0RpZEE+MlgSxQottIZl82XCwbnSbOUXm4oVQxJppJBImCejzWm6
QnIwuVIVC5HMvselcTIirmxNrFf196Zqv0qUh/Q1D6ZLpfFkMR/dAzvoEV+XE7f/PeW52T8YscTS
4uHHx2iLDOlErAPD+uR2xgwXMoZ3NdBptJMsaYHvbZn8wuYqTj0qVScjTVHKiyhWnsN0D/sEZhGz
4vGdCFQxp1/c+QpQZQ+OIbvY/2tO/MEoznIHZYnIO9OrIR2I3hJVE2oaoGOih2M0Sed1R1iJdkNQ
tXQAqONnB+/OIIPaho5f1UA3BPVN0goGcNevgcpSNKNwuXcvldabpTDEzygGaLu8Mv83Ichbyuu6
Rxa3KNInnSz0jBdL5ZGqpQjrAKgTlJghWcLIQEqrXIO6btdrh6FrKinEZvixmtgVgTe8AtEzXfh1
4Lzymq9L4GUF2JxA7sIrGBvDCj88F/bh6BIhI08HdAfkErK4idF5dr3inGT+2sPnaC1JmnD4UZuJ
GbEZ1uAzkORrRIVZQZlCrjUkKCYg+C0PTeFlYe/0CXYcjUsv+dpgX/iVsPm7ZMUuXAdGFipA5Q/A
ZGmYWLVcMMJn/4vTotH2yllQAkRrCm2/UpfqZmU23M5WJtXhF1DsaSXSYgBCd67gT35JAUfcEbA3
YlUCIgV5iuh9GgpEG8q7VwfvVV2gzv88kXFqEc3UDGVD4kLnRZSXhp1iU9CXvBbDFXT94UswObQ9
bEnmMzyCg+vNazm7vHgig8G0aXSP1i7X4/tRrPx1y+OzXvt9zeceOr1TYT0t/Si1xQf8HI7KkEWz
vv3qtlTz4DXu5IXgrO6mzXZdywd56f+NyS4EOBmKRk19ISBxpEHjf70sxWt572u6pSb7LVwc3/5J
KCFFr88/6Q5LzZpDcfWu5QEGmswGfMwrb7SFmNOaCpqxfenMrZ+3AXqKw98O0+3DApo7m25j6tHQ
E/wWfw2CqEHD9oUfEZxlAlhKpp+qdzCkFyAlm7ac+Y1CCi5ayH9vXfwIj/c2H/SLeq3LjaWuaJY1
pZj3xU9Iq35pGHj7M5UbZ6k838p/ZcjfBSMQLnM5+CP+rUXc/gQR7g+q/e5dWc3KEEaI9tdpLoLQ
sx2GX5d/5gE7WdsNPqf/Z7Jay82WqQ9nJUoNJMwJytXVeZOsErJAWHydHqbmLnpGQLkcMeWpMplH
VwZynb8cE9PBKG/CT5egWoiDyp0Ub1d+6WAw1ekjxXqjnGyYEZPCgyGqbppdh/33z28rQqssU4P+
g2ghEpdd/fVNdn/M28yH0w2yq2C3+NBGeyJFTC6fHibvijcFydEEJ5HvGm6APmzL+sVlampVU6oO
8dM8vjoK4QH1YNsRmT2V7HWXGxf+P6Ll+E/wWBbvjrCxtBYNhTK0KcAcXeOmVMBVn7SCbOh7CuMm
JMZrgHBmeRJvAN7xrQctMdRNhCJrr4EP/1AboMQE9N/+M9LvG5vCAjqfyZd6I5WBfTfaAyotP4UE
u7rOwG4dfLwJC7tdBK+eheuioALiOP/k+QYa3b9yvxR9h0pk5mjXe8e3KLl8p2BXVf7/mBBj49MN
zOON5jzay0ftUerzlw2xu3N7nQH8KXevNP36+RBpk3jXfKA/Dfhiym9JnM95Rd2H16EkBVPfT1DC
Jh/AcYhW2TQXgXfo4iW6gShpJIp46mDHJRE0xW5C6jFmfwc0ZHhRsPEzwEYrmWyKSeyitn9LIXgN
nGcBxFbLKFGyG2JtMQ4kF4pMtg0PrGFBtbz8PBJYujAbFwI/JSs1HXtp4LcMeyOOSVoTLam1Z5aB
VgC+g+jUJI98Pt6mR1KqYIYSUWzJ2ugD/7kY+BZqDbxZpL35RvqRHFCl2+fqe16x55puN9HF0r1f
srXsGGVQRBUBhGli7B0i6SMI38+GMD2E311fVntmz19+1dajdigE/gM+VPLDRjD5qY8LZ1v+iETH
KC3D0yJVkHDGr3/L3c2HGdrziD1fce+c0b0muo7RbvrlR2mAfnBACTGLdfkrRZmXgDLjw55Zh4DM
OsRlQ7cjNKEMnHu60+Jy0CQjjbGCmWX+K3fJHYA77BdlxXFACxL5HlHtpVRZhV4yeGf4FtP+4LBw
FYxGCs7oh1rGaz+hWYjdaRuEMEhx7GoF7IaCQm0/ZRy9eVsbYjGqwjvbYMI3mAbZPkoD6M1tEM8A
sg7g3DOyQzSCAqnyzngXL3zp0pPPPcUBhSI/yuLq8xNJC6oKIEWvTg/WKa7avYkqpbqh5hkgNxLQ
D03vNCFQTdWLyTCXcmqRBeg61JEn1oXcuR/GBa7m+rUL53FEp/5Be+JXJ2mCWCluMxqciTDQt5cv
hYX9aNuu8mJLRVXvu53fJ3rXpDQay//vaXUuB+o44pG+Q9YKP5n5IyT7j5NHrK0WhO/m6gpInG8r
FvibH23kOmhAd7HomJ2ny82YShnw6SIDjd43G+l7Zsk39Ep/TIlzmY2o3pHk4dwsq7RNlKNM3LqT
NaV9EdV/FePP1uzvDKPO9l6rFA4HPO2ADSMGfmC9zJlOnEmsZlHX0B38vb03AiLjZOZ7nHcaSa9U
Oj8Pe7kUPT26t5z5dOr/30vIvAVXBd80lwweYQKuJtZ9Qy6nA4HEODKIeqlR0LgDpUzx3euCOdqQ
/KxdKtHhEbuyF98Yi6p7Dl+wDilsmhKnp3Dyqrvq8iurCwlZFE6b0S8rj+8ZdKP9y0GWKKn4HhDh
tmiue00v/3qwN/vpmg7qDezZ+D+wwqjIwVr+AJnEQRwCLr2wt4r1Gm3XWqSMAQOJQ/DCGXMvXQbm
hLFravJ4k7QByM2mrfJ0gzbN1DU+nl0EKb2LCVJL31z/6QU4486KTZCRp7/dyVObOCrQ1oXugGYc
+ByFtnDGJCbVoK00hBU6+oukFoX4JFeax3igUhJ+uS36abRgclJ+D8fCun9pFQvhx5RM287BPB8+
nifWElCZJyC039pLzqgChW5PZTvYRYQkfgPPC2XTSVCbU+E+YSNkRhlRVvdUdcvu5ihdIgJoBF3K
J0XHhhIPYURjWQHhKmKwVqOlJ0OWYYxKrOzszXYolzipdov9KRhNDnq1tLVbuPXTZk2+F+Z/tj7G
cQZlZWbG++jLfz3d+mJv4Xw+I1tVrQqCz82Js45w+xHDW8kIaoRD3Kwxl6o0XPMcPXkN5yzwC+mj
xgDTzF85f4ik/BdZH3GmCSleQsce54oi6sA3ZkYI3F8dAEMuZtgpJQM9x8fzjyS+ATn9U//aLFNq
QJh5nOU71ZE6eL9BsXkim5JKSpG4fJcne23m5KkRDzvGYLWQ07IYeH8ELJ7ik4JBDtzSHPNNgRlM
zzKcWQ/nmpCWkPG6kzA4+ARssw7ffIEy6KsLGlydjTo6hUPafjJBqyJaKyzs8QpFvKfriU6lycKt
iXlx0yK0IJHWwCvm2HKW2WnG/XhNdRoRGa9wRXl6sYPcySRvrDP+os2/JJh/0r/cHT9F+1613sSf
N/yzEqRPZGDgONoHbpOOPzk0cwO6+M2gc3F4cotDC7HLgzUHz/KAqORf6iRMMUnzUvPJ6Tcfj/ah
ybB+8h3D4SBGrYXVnZDkNXHX6ey8lG4hWg+OinAKd+heJJ3oqo4HbRQdHv5D/ElfoE0kps8v7Gza
XtxHBNAM4rUuAosnYUlBH3gkP36A95cdXPHVLE+N6G/nyFLLIWNYKzIPCdeAXmSBcXAx+zBBnjE1
TPNcf5Xi/HOrUmxjcabB48L4TWs3sB3fUkb71bVq4KRO79jM9PcUv32DAl+iPS3XaWzBpJBidFa7
wD9q4M8nct8bwvwHe5+Fi9NUwjfamfKYe7oQ90i7wSfkW5GOjVys9a+JiN3FHmMUmTjQkEZG71uV
J1O9sq9BpayOzygoMY6d+wkeAcGa+6OPFLx+y4zKXfd/liEHDBW7tHKT2Ae4N2bga8Ie7eZGMzOB
qxs4k+ui8s/a+AHKjtpxMrZC8FkeNM9xN+dO6l/+PmjZO+t6s8gFFFYPM6zW9GklQUigMzZvfkIX
So4QlupVFaDUhBSZih4ctZgPPfe8g3guCCMRbe9AJauGeavJ5AyUuaqaohH4VlAPIT1Bhpf/80Fi
fFluY78wH+OD8+xqKCzdA5F4NFF/N7usd65PLGsKJ4oCoLYSRO2FvKloCnPRf3zRlW8uoy4QfoRw
sPnIKRcpv/kfgbH3m950LAc6+x60XVzlsEX6xoaCAww0ci2vZKGte9NgnwyqjYLfJ8qVrG1Aeepx
wimfMjyxbONuxEyxpvPqH11Rc4CzJv8gJ7sSO9FZLXGxzUY4SstxJWUEI1Qzsxrm1TpuGzEpz6bz
iwmdB9C4IGe2BsKeZICa5oy9fvmRGUa3RUrgK+vRzCKbUGm9IpHgqaZheIw6/QWGzVETNkRVPQL5
y5eNTj3ANtR+hzsTcQPNzntkMSaufz+dGQ6DlpJIh/Yfy95Q02af0jNuvGm1IrXfqfzjWf2EE7iI
sbZ/5OXs6Wvd97HjXrV5E9PZ+1Wbb/UyFcIBFO6ih1l2OYZoLWPbuNiUL8ER053xSZ+2HKiQLPiO
cXuiPEn0CkLrQ0MZ7J5aTN7sDGkAL15MEKY4MIFiTOmlFnzfuI8lzhjv/5a93zETpsfsfIt3au45
YBHfXuHfYsy6wSThVKpiLlfYT37CfzSjs3yEclPDq8ycfs/mZ+NEEtBdrz9jWNLNiN3LV5eq1bF/
iFuAQnzHs0WKy+emJNjMEncvdKYSMO0b+hnYQIDVY/Vx3qnwvdP2QKQU+J66VIJ7Hx8kLNKXm3er
wyUURCpDZDBwCLM3FCX+L7rSM15C0ubcN3AU/80kIjAo6uh2XcVzK95nGLZ5DoxVjawzVPt6MrD3
0LalMEKcWOs5R5r3ZKCQQlPKkMfbD3OiuBlcMOeOVdUEe41os1BWjYiQtGmrT9RBPNgQkNe5ZsY6
Wn1bUwmzM4+bfUqeVVPtRM/clPuydnMUNqWZ0uQpt3JYUkheB4/DXyomV1h83NgLj0x6+Gpa+wrH
ToUPkykeytDKqk7fZu58MuolMAWPFmElFsi+P9JTietrRQ4ZwkDM73sGnGrXGCSI/lbWAXFhSxXS
zCLPtIJD0NnQuFuAYI4/+N48h6gaC+A8Wrey2DskseFcLwLjlJrp/DKgFnRp1Aw2iysjLHS7aSGx
e2yiVFh4HTbVDs9SzEU5HJkQGGlUv7TFQ6vaVroZE2B79okMxiL5NktrJCyDv7DomKwPgm1VGIVI
PQ0LkO4H2X4MCqcuwFPZmov8jVPKHELm3kblCWk4JszO/J04kkYgoZgJOjoICuCuydCVm4s6BSk5
R7uk7bjRFHsf9E/uKuS7RwqQCU97/E/4uJGsLygYCdDyNu2SWHWfMnwuApAEeSb2FaeOc9YaM8Oa
UKMr7INT+Xt2LcT4Wv/LUVIR/VsFq8D3bM5WAoRY+oxSOvGL0Q3749ypQyL6s3LcQajPu69XiAsA
T8WiJENc8y6BzCoIVnxF3U9I+Mqeo/TkUVxdEEuG9sgImFOiQm/8nupTYqsdXiESW6UWBUSpdjOQ
gGsxTGNSWMG+CHsgF9RbOYLRDSSM78OKy5rmw6j7Jk/foOAjOQZghV5ZEMUQLJNOAGQBeDPaQF3m
4ExP5WAGX6xOXwQgvaz3wW9xMAyCViXcLcMtlLpxUk1AY1iqDoGWoK9yNixtvz0DfE5HnelMBLnE
XniUUTSDYENvZtVDf2cvHbVMyzDzew7F1YyEB+XOIp5z2e4kd/9qjJvDkoILxql6NgMcUgGbImD0
GUzSzTRkxKCJV/33X2PiNp5v1oUWSbxag0xGJZRan6Sy2FgtQ8s3Wg3pyQS65cNNElqIbjvMu9D3
7zuhbSo0P7FCZORQ3nm1WGWbKpQnvKUmSPHYR4gKWeBnqQYbVufjR1kMvtzyIuqpJlmUXjxP2ZMu
CYuwKOvvCiyrkphXORUXmSZElpXOWQpO98sl+8uSpQtU1xJGO1eEzFlSmK0PTKJuMhoeiFuG/ds8
Gz4I3oQ+OkkSgwF9skM/vp2dczBpWyZkYCoZsZlbp+Ai/Mnd90Ue6gZjxFVsWGhzbl62PBhVTbtU
YE5pBVmScuCzLuPCOoSCGVAST6bTXm6IQ1K1fOOG9p587zXekO5r8eie+PYFqDDHiGK50wgHDc/z
sBmocbvgtO2vnbce0n92RWeqtN5pSmiASwMZWzpPpAzCHCk+oJTKPP+e4aIXe8a8kA/qBTARWD5T
X2H9SE/2ryrdCOGsq+/gdQ2KHIUK5rBtZILxpabz2CkP315mWDuHmkW5K4ZiBsKmIwOAp9yjCOIk
0h9HOvYgyH30iBnYP1PQ2sguz9U1/NE6H3CC0oGWRVTUHIdofgZo1MCRZll3qjNa8IsAhAiEcMR1
HKA5iwJQW0VBcndpsLcIfpYd2xr1pLodR3Pj377WOCBmS1DrOcbWy2FZiRqEPwY37kdir2KMGUF0
SfSHRj5PFd8dAENY3Zx38WOp/0NP3WiHJWNO8csGpwqCSxpjQBE/i5NYM0cfhajOq8jgkcgWK9mp
Gn/ZdDgxuXkfBTNZDOqMvM0DYDu138HOvDd0mjGLCvFcnV+qn2r7nD5GF59iNwrxbxfgpnVnXb0c
lRY9IXcXMNQDrR810QDlmV63Sh9HMfyrxzktUSWRW3oMke4T7PerVRYwko2TDM3nDbSm1BbdwmlB
can3hu7hBXN/vw0th1TS7RMsrC8BaySTp5YyxGlirr8vi/Gt1uz6L4ieZG4o00qTPN8fzTugp75w
EkezNK76Oyzl8A5lJ6Cd7HphllAtS9LictLU2E9QduUm53wgelumgZgDMOnsLS/I/StQw70ovawR
cL4+HiXiFn+j6ZIY7KYjjxDfmpBjOwPmmSR9WL1aW2aWenogSaIl1LyKlcfTQ75+AnBNJjDYXUyo
4G5QjQy/bZTn7MpzBjenRBkWedeodY6Rp1P4exV672/puf6GnVlaEzmARWuovhGILbRCOvGbx8ri
BGkWUVnY9WsjUowad21l5Dex7ELVAR6o4JVsomyb13QclES48VofjlUoRBqs1U3ZHF63q/feCauJ
4UfadZ1h7z6+pGH6goW6gC8AwZU46mb5WiQO92Fh2/WbLt6W9/4joio6MeqoKc0QEmgffwrgkKgN
Y95oTeFsbVJixTRY9+7tlvv1QwJKWUiMTsAwP6c2mMLqjs3SuC+ALH9I6X0ynXGzJ5Dp/DHlDEFU
IH315Lque6PNTeJNrsaaE9xfugJdour5OUj1LXDMay4q9Clqx3qDPRuHdvcDRnkgmNAxuwef9d30
upA41VzaWaMvLyeHOgvP2eBTiKbnVoVSsTkH4OEKE4uvSxFM7N0tNypeiKLyaXrmL4XgMXdID6Xp
s0xvHRpmKGwtttX3lcDZ7zUTja8ZeCWXiSiwRX9aJcYE6SZFlWJnWgI02oz/eeMjBJCsRR2M2iC8
/StrYhYvzuD4qbLTirjL3regs+wPsda5BC5usxMgKHHyv8s55DbniuDNjTxd9iEm+dqv6/+DMUAr
v0YFAVUuDFLwmjcmSKbkLOZJRgel95TLiaJ1ZZPPPZSLXjGmMUgsr2Bk4jgYJSdGBq1pmoRf8JZ1
j7K6yiigj33LC8JE4FgVAqVXqzNFwDgvPD8TvNn/EanW6jS3kx+orJJnqjZE6KX5ZnicFxfl7rtk
aCSVgUo43d1Pb+c6ZdbFuChzZTZfh6vOuLFwtSH/RdZZ3RFyNbfVYzhqDGKifExN24wt3uNYrTrE
bflCW+KCTezmKkeiXtIobJP4hwgH6DYHYTrAGDATQWSEVJC+j45JjauXOCY0iYSM1Ulf2VvzCkAg
P43jikWwhCjDtzz3tVZ3/xjlaHzT008WaV+AVQ53dNsZMuyX2uBQi2qXSm+6JONJsPFVbeCI+B3g
l1Ehi5NGNG10pFV43LOZhinxXtPpk1Znm97hlV0eChhSy9505U+Cb9ZNri8T804hIUqx+U6tw1Pp
nmiLuc5Dgv0ED+rakviTPa3XqUQOpACUEM6Kao7tQ3BpUbkhLW9JWhIh9/34mf01qTulYIimIPkh
xZz2GTSepM2VKl1SFCNNjxEFrax+lH7T6tTh6VPExi/jGX+gs3ajDaEdh4UXgfbFKKNnFV4xGE2+
wTMhhw238ZyRf1fvh96EbaNfmVMTS6ZeJQfRAQFTCwfLpIpFtULjWmwM5UJq36yKzzJ2F+WZMre+
QQCbK3Ho2VXRno+ezuGSwLQpycbqSqdEwiB1IX8QONIzOSldCN09x9NOJELYEJf0NaUtRXCiv4L4
LoMJjYOdC/M4Mu+eNhDsUjigXIlNFTVF0KAYCncrLpWyR4V8PLxguZ6uvtAbLOOSo1T8OEMcOozL
oF0OuLdhYeZhzH6Fb9MH72NseXxGaH+xyMi9PWRevvG9fbg6+i4EGVQx1cD0nUCPe+4wjrF8pp6m
bMlVRVB+oqWxXE7YM7JbDiyLDLnHhLz6XTSg+qFWksprHjkb8JMJiV5drZ+8drp5alc+STzKxAWv
Gy4jb5jgbazP1QNjKE9dxLK2amR9N+J9FMAERk4knx/vBe18WTLlUlCQpDngajzVXlmaJMVPDQZ8
1aHeFaiTvaROVpn32zOI/yFkDTgJmDnDH59E19I9TNOqfJOCxqsRldLVwRB1Ef9wzW42aNj84mmv
dobzCu9MzObRjt7c5F+5R4dJp+ONtUFdzBLtmo88ft+nSk2zVpV/qYypUF52Xi5qqaQEtwDQTDOX
IUNt2WASUYdke8R/O1yylpR+ShYknsy3FW0sRmvzCRmxhLx9TIe24TsNbVsaDTEG3SZqQo5Bj7cs
ThZD/7ZNqgnY9malWiVKS0Qx2Y0xpvjrfz5MTdCbnTSOWGNu9B1g2O27SE5nSN3mvAjPxnJ5+IQg
1sm/qAMFo5B78a6NrBxAz5Xi3bs90ovrpZIcPx0PKDktmRZOm7GSN2DiAWcx4RgnTW/6MRVZV/EM
xDhsGeV6GbahWkye18LwJmwtfY+DwbLHfT+ptvq2V9TQQBn5eEKxhqjFGZXr2ix4DtqsU7nbeIFf
gZ/CSRQCDR/Q016PmLlsKRlYGL72UyGM+aSPS9fXBUh2fAnw9Ek37xjDSUywc6eB77xeGeT7fvjL
cm8FidnlB1dOylbLmgZd7riI3lBQT7yxuPs4fuCKq66UAitsi1TRVxX/uZSIJoRS21w9Bbo7yV6Z
lz29PjNc+09zWiWKQktkZ4pf4XIi5sgI7wbAbtcjB+SmC1VTeCsOzFLxhWTifGPFpDceYc7fMy71
3N/mguPiK/xmrtTELImxMhedcnhqEdT/Z8PqJHgFqDLq0lPPBuK9BN5YQ65gaCgdUQ53GiHMKcjr
HHbKjD9MGvgSFIXT3JzLBxX1E5XIUszGKmRmPYtl9/dEJMlYr6mUOoCUslhinNWfuPmLWnNb1Q7Y
nQgtv/2MqslGePsWMEruhsmjziVu5lJUj6hd7RFYuY4u2bgmEySQbT3eZNLU4PTD1jh1c2xmdD8k
aB9eCwA9svsxrS858xupdU6uH2MwrfY7/szPrnnqYptaepr1f46/ERgjAWNKdnXms/T82F0UiZJn
wsvInKZUXwxjhNZlCW4kedj/BzCWSo+KTUj/JKgcrhqri/4JJi1K5OgNusJfUBqJN7HA443e6JPx
/Bpi7kjnm0UU/ThJcnHvgLcvb+tsymrj+AN8oRmf/c7E8JS2ruzSLJwaJiLLWLaDt3a/8OQLa3p4
V7F+B5O0XHrEtdqJ4BEv830hiDELVN60a5XPs96R9/MjMZlp+ju5NRnUFgXKaT7yP6epWCL9c6Wf
le1v6QskLYmeNd0DyYd5CHl/ipEo86cLO10kJB00CQ8eWhTVg8+dezV/r4JgvAVQGbwGO4Q9/COj
rLDnzxf+dCClGN2SLgV4oqwJYfsHYPEv+ivZ9d0k3g+Ll8QUFXoVLsUYAc7p8kxWyQ6iTX3k3lzg
xZPAuEwjC8VuUGWmdIupeizsUwvfAAfWXXxEAa4xTfXTFYHi5C2eTh8LUfZABxPehewWDChEq8wt
jUi4sLCoZtYFGwDWJgnqbbr5wmL1ttY/nuym0BpTJ2J7t4uFLOoTftGh6Ft5XYJMs7dBwk2Sjhqn
wyTK6Y+0FIadjOq3duMeTIWI7Vc6hQ5x4a8BUU/WJTKEjO2TVtoFOHFGQ9XkSJRVvcXRewQ86iwr
UEpwRunJTcWVFsjPQ38zwhc/+TqT/SGt7pR9PRKcuglZMOGStaHMgK89ZK6/fy7tAjNW4wq++H9f
WoiSOSzbyhG2rBruatomeOMEi580D6q5704czSOnhcgMPN+pVq6ToqQQKSRlmiFegrHrICdWG1cf
j/dnsULkN1F2NIBd86lV3UmXz+0FcXf8LGLmU86ca7OptTRwlZZyfc6KhVZI1tdnhxPr2DMX8Qh+
PLUSDS8WxC1PFLJMflmciy01b6MkP0zRPBv2kZbf+Bhf/onIcZak6tuy/9XXq3o7ZMe/MGuTwvyO
+b6zVpDBKJNrO/a5TyCEmx0Yf6gNqLRKIJalA/TPHo/GmJSEXE/sO+HQixAgbf0cFGdPLcX7zjfY
VrJOlvIEFcxc+fG/8KNgNYGvRtCMvbX7y+wtLYw19d+io+nnjupL+nlK528bw299EpFLVmZQ3/gE
B1Dg7fw6N14oRXjYWp6gA8w/MYcCktA+g1LTh0yGg/5X36UtuFKdFHBUbEt2GHcApiXzjOPa+frW
jQcuKuWeru2hzrIsZPlwTH4oz0MgzWOxBEQzp9pj+yBM7kGAqTahwgO1NTAENmlQXuTws/XPskkY
kilv2UC0UASM/epZhlAmwsk4Q9WP22XsVwah2sydqR+cA9jguLITvO9o4ixBGm25uQ4oEo6wE8Qk
MoVyti9ek/rDN8VysHPHDWx+ZDBALwUhue5CRhcbPrQziqF5HQXmu4/MwnppYVCn/ZjDPuwrxq8B
ixdKVmcu9svmO7rRfXB7Szp79X6FtHVmnd1AEEy1xA4c1vFIGayu5sm5WghocEqJ9NIhHol4B07A
Du+USU0AHEXo7AKXfmSrJDXZbIkuXSHd7yf8SVttiz1N4XJGbIgVeOjLdqe6QOeNYH5CiA/FyL5I
urOukpwtapyIYv+UWcZ/CeOT+qwcijr2jPRIWWZP2iaXQhZayl1hnfa/NVeb3NPaslZBtRLFIhUA
MmRtA/G6uV49R206DgFfuVPbWLDG4w31vVL2wz/karhNEVFy/1EIOmSqIa8Zfkc8NcimSlydkLA5
WiV2HBaow18/4UOhVC9HybWKD5v2MIagkGqrIPapl6CafYiLCrsohX7HUyn6xzmgEqPS38jtWyM5
nR2QVP3k4eDS8Ngg5KxUnwRG2yDaGLzyWRCAIXiPx/1CrtUq/1NnN0F8A/P89gs0cfRniBN6JTFC
MAwdZtrumPT1RDCvpFnCtuJ7g2dcPjwFmofLXcgmcdaX+0QKY4btE1eBoV/DJfBQRlU2tnRxwfc/
L83s1TnB4iqwOEZSZZ/uTU9X4S+1ovwQr1+Kk57TveBOawcIBiA2PTDp87vKDVrw55xdDuXLbYvl
YhumCh5C255sxyw7I0b72oZqNU6UOfs5jYcnkRGcQ7GZp6135ZhJtNOZ79Klk/LB9gmo3OUqdd4r
yD59bp0D1iZYVTc5xCNTl3t7gXVGMx0PWJvKXHFfuXCclHXCxDipVYLXnSI3B8Ps0Z7nRcGlImBJ
IetWq7rEw3hmZDtPaXXHuMztXIogifT69VRIcpPBwFubugzD921zWXL6oJc53OzUwqQZ98+E2ccl
gYs+QF9FhPqIzxB8+F35jszCKGAjJlVpB1cJXpb5Tdkb9XyhFzpXfNRdMLWAIYC1ue58vsn0knjN
31dMzQAtZjSY2AFR8FuhRd5gLDX/Ft01TLWBqKUSbwA91ueCr5BWCnHZVtaStDbq7etlnYnGop+s
9f59gvx3c9BgWl75/JvvByuXcMzwHfidvuULXvjyzJlCL4FqqkSoghiku0VTB4DFvKyEgglyn+p9
zI71CQNEu6t+5Fu/rFMWaiUYhcUDSdHmW3RHPWXYVVjiu3AZc4JEze9tTvuEAzmcsvpufy90xgRB
Nk4m36dCG9DOfEwHpHByM//Q7DSDNnBijotGF9ss1Om2XNY61+8wMEbaajtz13S3CHlBYTOdxFZy
YLEYoaWiVaS6ECb/3CrHEovi6WgpmUQt6G2gpVhzY8T80sS49iY20ChL5CBbSc2q6EKQ0jKBvAr+
Uce45Fmb670lnKS4fxcFVPXBE9Rt4v0hAucmeDzMUfGtvdbWZavTwjmJs+SlJMsyPa0r0S8xDGYU
/F06deHkT4q2lMOgZJ4zOfG7ZgMWqK3Y0gPlwbdVlDS3CUAKI53434ofuFmqG21LGYL7KLb5UJV8
lxhRZEQA7sZdT+/nxtie8iB90xA2PPLnmXM23mjakj+JX/Wv67ScnahGtFYMqrE6FktvmmnUOpRK
tv/jdW0rspxQzi/+R29LXCmHsv8sjvZp46xzcVzOnmwu8e8AoFrThjZyUTEP4B5+6ouW0+Ooijul
7XtfdSDGSCEmOSNKzxlwT6YFZHBVsNrE5qI4idnU4GKAkTNIQIzbWt6zEIgRZ1NBPROt1Juxusid
zutDc0nOKw7tLLIOjWyocG0TNcqcR+OU8jHFvV4AVnOhiRT2pHW44dgCgAOhHK7bUBHqcv+ZFudw
BbwTJqUbZbRafxRFTc6DhB5OVOoTdwTlGbJ5cwISD3R/JjQKqsLVDv1qJYS2xGfqxis0d512pDuN
YKjrSc/Z6yEp6PaQ9K3fTzPoY6ePgPQt8U6Eg24Gm+5cBGC6tBZbsH09CmBVxBOdmIfjecxi6sDf
d7wHyM9huLhuzsISRciPZQm3xanf1BLatU7XSv18NYd5P8dmzdeoQCCk+dIRLGFQWqMNbpzjdBy+
SrZLlnjhp/8OaCXUadkrrXiDMKdcUqI6h1Cj5NMS0eXoE3Q5LWyusDZ5QXKboUzci3l8W82XhWZ9
zg2DrcysQBfim4bWr/uKS3ZwWk8HEKfo00Xgegjw9751FxeaGhXpr8QimCQQhT0rMMt92PZjWN+G
AC88KtINm2Bufe/LsNJIkj37idG7fw1Cv0hQiMST2CuYW/g/kuv1NzmAF4r2kmUoK9ttouZ32F7U
gaDUgyVf9onPyoOdYmQ/HJ8HuJ7FB0b/424iA2XWxe/laqMRbzJh8YBpTPoRHkymsx3+lJ2FGFSS
U37+gJjnW7jzH/d++N34Mgtpn9WoWFLitgIMM+tracUwqAZIDM7JhZBFc02tlE0K7rzATwBHVlXm
As3d/6L2Q4ndyEhq2OVSg84EioW8NMAaC8onFWpLEReTbZX+rta2qRN6neC0D+2RO/bN9OVNhuB+
p6U7hLLAJ+QmCk/iVLPMp3BA+pfYGGbw0yv5JD1kvxkVLawBwAaacfy8SQ1EWQfTxEoMtBIH3sWp
6Cv1SoqMDQvn9NvN5cT6kPVfY5sHdiHZlwGEupiWZV4iljVzSewihlKXkY1wgsF88AcIfGRlGtV+
fZTRsp9SImicOtC+zWhOSfXMyk1aEDQtcTV6cYM5QPIWdhna1jilepiSDH7rRx7pkRaBUISUdO7A
wmLvl+axKXjDxLNWGqRtJThDWZgg9tarz/NYDGqUnLipVByVVfRl+6NV4zwo8btE29CpXEbqFXcy
l7BrR2d8kxT4Mx9qP8o5rxZvsOQZftzX/yxIx1FsRKMsL6DlFTNJ9vicMKmfg06zOOA0//yvnrhU
gIy1vCpKeAF1qU2jyzR2bD4Yo6u5zrIiYYa3g0RpyK8TD+1+LyborX0epC1pHePm+L1a6wusg3z7
pK94wb6JfmgqNojrkBPiuGlYOSvf4zYjDOfx8wdXfzC/VSWnMOFkLpiS9PSWkwLDeWRy6bR5pxoy
q+BPnksLgJ5UwdWDo7afR3LajQdVm9QbmyMfcO4UGWSzbSApHKZbicrGUXrE3Aqut4loqO/0TmPL
kj1GuL9VIfEPG1forWQGHPuy6EDyB8ExYxN6XukhVfyofambxVsHxre1smUCwlE9sor0cAF7l3Oq
dikYJbAi1Lu4+qN0FqUSCNmspI4KKhHOHbTtH3OMk4Lmpuolbps4CQllIrvFiTVbNkbYzp4YCZNI
Ln++9Hq9nvv7ItQGOBZgsCIGInbaWlRSPLFXDKI4zlqNJ2oVGfGMTmD06zKZmV35bD5pJS4n7JbO
+yezBe3eNF3txgc2SfrxYPVMh9IgK3JsAxNN2nHxlyKZxR8goeBds0Y9jffA5r+xTbjpR84n1SEh
bKUU/EUsTEsQZh5mfE70sqB2j7yoI0FpfR4MpiERYh62l9m3ynrS25vbMSe0J78zfcYsScN3xgpU
kfowBfiiEuAWQmoepFDHMVyGU8oj0X7zZVBFF/0dxmjrKHjbPLZaoQF1EyxcCCMKQg7hK3LU0krS
bP1rJjV5C0mJ/Ar2nJ8KAMhpwNNE6NOuC86tVnTz/uN4h5SVe7vltwiSAVYOnUJpjQths7Gvnx95
eBhCZPOYE90OcR+XZvb5v3VCqzpQfHVOL94DRjkk84enUWst49mc1GdM146yWoNp5yVHUJy/Sm+8
2sijaT8J0cfK2Av5Jp+vXLByYc/pbInDkvif8//ItT1Ge9sQylnc1rp42RHpNVaQ3EHexfkh7qxg
BsqR0BFmymxLiJhBRYc9acyZx/V8DEv4A/1z7/h3KVvfP4+2BiJmE65qm/JxLXJqf0U9eQW0N9Bo
MPcTCH5ARNCdRVvHgdIWgZIYQtw2bEYl7ceoTidYVZqyQ+hXYVGl8DwIdsMQ/7BerDH3C1B/5X1g
gsfHG+ZT3hEEmE0mTiJ16A4OCIdIDfzJToIzDD0/8XyFaB8cI39fXKOEFO5kf3PwkbNFeFI2OMnZ
jNOrr242cvWfCh5StG8F7xYF0wi+5M3ZpBXX88KLrU1xbjgwLiJsCZgEN0LWPx0acF9mqMNt7gNc
vUbIhi3WV5RMOjW44imD0OdyXODsZAlYTvh1tLqtFwbiOJGk5IUeeqjKF/IAGdEW5Io78nYwaXl8
ozFTn73b7zXu0HUK6dnD9MDI8OzCUtIPIScdNOPiL28aj1S5hIrjlaQcuiZOqIIEnlD/ow4AkEAB
EsB6MrOf6WQGj2sVm4gvxXViD0IerHLcW9UNhsT+zdbn1xPtW8P740hYgiNx4c80MsuaMToYJZCk
SSSfs+s30bmhYmaGujkjOp/9zkH19TOXnb2fhkodQ+AgdP4WQwf52KH9pGSYJaKY0CavSr2qAxt+
vNoR5DcPeo/YBhezrOaeaKRE3Dxx2F/JR58WUrvhZnopmDSHC/ui7Bq0V6jJ/8UPyd0iyDhOzXT0
i4BFdJXsQMQ+B/cTtLci/+ByIxzC1uCH7tr73MgzZAArRrTeM0FqmEg1l56mi/dPE16xgR7jS6MB
CEc80QkfQa8rFOIWM7/09loYuopz6kznMEWNatVEVf8vOqT/CWY+t9dL6/LaecLBNSbnNfvLgPwO
VkkBcgUCC3yjWq4f8R9Ef+suHVAh5vrgaD7O6uJRX85WxvvK+TJ9mcDubLSBQhDxBKXrlQW0bxWB
ldXCp4nPnpyetMS3hY6GxfofayJuF2Z7dyMW4iMLYJQ6DFo4Od+5oVaK0yfUPsGMP/JwheiA7s/e
XZYh3P52c5TVpAmIffmsSyUUjMGMmiliRJWOdqOAilvfvTAVIaIFQvRT7oMRTW1J7H5Xwtsp83Xl
jFBD4GUr6JwNBaUFygrW/l/psBg6dr7XhYXVTBTn8EK5iVSZW57tKrww/vB/Kg20JaxDZWqiO0Vt
UXfB0WU1qDSbUzQzluyNFt0UJwWCtPs26c/3T9Q6YzRdcU9Pa1SdsFD9WQpFk5zlzz+1vl4cD/st
hafIr4ab4OLv313J45kVR05+xHVCQhf5yMK97dSeXztqnRsKt/bgwEtZFICQdMlZcVGs6YlThsVs
jhg/WKlfR0kHpkJ4JdqRgGZDeUM87zRGBLp+iZ342sytIuWVb+HfKcCoN6yzL+Y0QObUMmfGkLuP
2Rx8jq3soZV2z2u9gWfRbJsMg4w3OIoUpY87/Xa6xLbHQE8D/gSD2oqqP5L6GV/Wk0N72EfYvFad
4vyce0W0w0nyDOAMHZUGH/wBUQ+yDCCWl0koqSWdiwVQXJMY3rk0rOFKSv2d5fAMGP4Ayc9J0wWo
0QlETrIAU1Ca65/+8f5xQJtWNjkp2tm97ezWC767rSB4AciHFedeKcfysrRPj3vZpUkhDdCuejKY
3Xb8ABGbamUx0phTcxwWV9MxNT01Phg6t1l23i1He+NPkhjS+3d3M9hLFtcYUF02grWlzZM6CwOj
EQIk+AAf01b0+qIAoHRHQp1wyct8Y5MJRiEJhaNbdgwg/0TPSehl5moJcXqCjqlKaWtgYiX/lLwY
Y11enB5n3GY0C67ajbunnqtaJoVEJdL6h+cOmJQNwkxKi++9orzxZoW7pzKC6WLN0wXL/NarK9ax
VIwGSv51pWO+Vzis7ptIbPlVARZ04Bkq2AOo06dB8BqYeTubE1JYtRtFzurthxG3H2lOJPwyoxEe
Ogv5+LdOGARzxOYhxvbrAbaAKwpmnL6zUE3fXf10MC6MLdRxTR3WtiYRrINTg8h93SsDTGXDJa2P
ygwahFMx92AOY/6GecrGAUjcGMJb8+RcTxcBTvnDgOPakxc9U3rYoVCxEYi+jbS2hsgqcooJK5FW
RYeFeRdSC0QcDBVAQPrKJfg36thXUma1pDQxBp7KFVlrO7LzB1GazLK6gjKkw3UoK59qbjwhB9CF
eTBA1lP6ssRUjidmMov6sRLlIrmt973Foz9Ophrs/hhbMBg1HMmEFkkwao62YX+KSSAGXzWSjeuE
vnGKUg2KUyYwdUEnABSMdtQl2qVbF/0MgqvvpySRvOL7itbQdTbfYcAOKNGekc/lYR1H98jxTvOp
CAWvcB3ZXAnPPt3moxdF/AJHiW0VFVsM+uS5U2yncktZ9YQmGMq0rKhi487KH5ZxrWpXfTlFm/i8
20lqWrhCU8hn63RApIn0yrv0N0qP5k4240J6fXXtVuA9XdJU1YlYtCnydyaEIc9i+P7YclHR1QS5
4zyeT5kkrN0OqesiH/gPwQM32LlPVzCt3gNqCE5S9Og6SPYvAJ6pOxPpx2/MjUDyLFIZfdv0FXIi
YAN8oCNqapLTWeqAVWTVK/+5E7kT6U8bafy1NIRQ6uS895WvYASR437al1PhcbQ9y9+5ugtswP9i
iIaZnuromB9e/Bsu+G0csSVWTJNVlnhspYnQ2rRGQ9lzAa209iZDCGfJr6QwGcbxC5iattaYAYQG
BMHxoLq0/KUcHL7nB84vkx+nQ+qk/jPyETuScVoYcTJz44dxH3zpNwwvaxU2CeUXuQDJrBlV+ACc
WLyIkilASGTYmdO9QHGCB1quvPFz/s5rPHFWAXp+3Ye+SvwB1x+xAiYAV/a1xT87kl1e72cPklOz
OTNZOJKbVoXi7/wiMoEoMWMC6emo0cbikH98vg9sChZipYPNXhXMN6kV6MF6LU0CFMStzNOBsyYZ
5d9TGdx64AofZcMJZyQt8GznO2yOs/fuVJf2qY8H66b2vWYPBVvU37GakwMag1oEYqjfmdL/7xEA
nddnNNPlBeG3yt8uQysut7ryFV9NhlT60HlIM4OwRErowrj2Uw6okkwF6SXrHIUeVtgdXYQO0pZs
GSYlLO87cSHhCEmqZC/frzQ5g5BmlWoyfNbfZ4kPu+2/BgTLuULJJCGXbNT4R6CU1zHQLghJy/jl
nyt8pPZgzNtpMjp9kxyGH1qM701zJB6c+hN15B4jDsoaRS6yv7g6D0iu5E61kskRyl+juCkufMj0
7mIz5ZGDax6vsBwwoQTtsHrvLnnJ6zAD24RWIYVvnGTMQoqEarPYloCe0IomweQCCGbC+AmkDm2v
t9W5Fi7CW2T3Ay/a6PB2xNWWZLvAhy26zoFve+usOCXbxU2YKEedJ963226YnMs8yQk+dwRWWt9u
Cl5ATapMt4kToLS7bdBwYDiC2DmRq21gnQSyL6sF++goTaEdh96xBfgoWHMLelrIHCJzM8OrKCjZ
hQ8wt7HwD0Hth63gmnhG4nUgePK1V1FOuq4Bzc56MzScTmYPuOFNZ8SUTCsf0OkL7Q/a9Oj4kLac
A1sNZ+dCyI6VZVha9YSAWLgSr/Y8csm+LUytif3Xd30GbApvNLzSqMUddNM2DA6qFZ6W572El6xB
12w6Q9Ll7xj+sCugb4bOjdxPM2TRzyfOEHIJ0r+YNxbAmNls/1cP3+QsvB1t5ufNUotZHfzAO82n
0vQA1KAS9k1AKtC/nEyp/zwwe3xhWKmBIYMB0QScx+TxgZIMSFmiN56uWi64xLKCwfu3FfoAtQMP
7xYLROdV2Vjzp5h5WUTsVyfRehv4yTkTycoy80rDX2Sj2/xP+Fondeyl3YpVUukjgye463GsdD25
JNmnUVcsGmw/Hr7B0kjcns6PpbJDoAenydh7xzI9wZIROxDD9LZ7a/TF6K2dFpTUddPBaFGCgZDn
j3239KCsncP7JDmdZgFQvNePW3y4q+021bkFY98+gZqzhrx8iiiqpFs9VER9QT1CVao3SfNjhLHz
B6ZpyQ/RdPAR8cZmOOXsCuvxK3G5fPwoERqDwNGb3RALPjHoS+sGckWbw/688rt+HVrpNmN3VJsB
B3zNZJrrK0GD6xAYaAR59wswufLS+TAHNbJeeUfB3XNYrC8Co3YIs3lvkAJuywFDX8qQ07M5jsRA
OwaIksc0xUezzQEWym3ww4lPaQnYMgn953FE+Xm729nifrlFvuXiDMEBXTdfLh5aBDAaEYgc1wm4
WwAQNCoTrL4hq+ImEBXaKTZKXhx3venIOMrc5cExOPPkKUARaO1fMw9hksR2dOSmA8+H/j61fZL6
5mVFre84g0W7drihq85gSYTJWsuAErWg3e9XTBJ8YuFlmCJrRrgX3rVj/AJr0yWtzvp/CJwERvC+
qKkyxmdBX8qcNEl8cTDRXgppYTy52aZ13kGbsZl+fxUp0ECxUkZZ0e1enU25pAh9iG8GXbu2PA3w
w+7WJZGXHBBfnPBoYuvOl12Su+Q+lyINP8ivLWRi0cmiw78UDwIiAic0CyglXzX6lyX7jKOFk9mx
Lq2MvsF+2JRIFG33BxwyVMDCn0oq6JKxp/huwu9LlOrlM+9E8qGaQ7Fe/FcfBPTM09ei4vz/IBIM
/SyHqwTuKmXGNoemZExq12Yg3+m2J+Axog8/ZNIf7H614d0mplLNIACqYFA1LPh6I5+qVvLJUogg
m5Ar3AS7NImKHc+mEC4DuWIJrq3g7mT7wV0quHxWZLjRyLPM+unleD6h6gWa54ntmrcvaWutdii4
v+TtMXrFv9ZQRM6y06f0pNsUuuNZVf82DRBVe5Waczb79Zq55wBVJKMxyd2QZnXLBmRnSdhwsW3n
SbgJu3brlSwhQre0F8rDz3245jCAFwqh1IAiDYgb2EUh2Pb/9hvWZF+uqFlgcuQzUw1mxjIn8dld
OSf20+7BC8SeS6Rl7ELa9Qk7NKbzJ4H2Y1036QmARXHZRTG735AR1i7fhw9gpwuPgUqFm5GxxMFV
QUkWnQbWriZty8n1MLa2WK+tjVSvmrUAZ/znqNdBufeGhVCZjMsVvvMCWoP9EU6ZOdrZP9gYNrOq
ZVYv8rpkol43i1iVJLLaW62Sx+O3IPdCJsOJa83OLldHMZxpCnZAo52nbRPFvP1NWVKq4siUScEA
52gdfs/0vyWfKaaQsZHOHPPvAH4fQgVuZs3a/0YwkKyPNnhl4KnGqFgZcjfILKhqPJIn1QedGGZL
zZqjHfdKo9RXHEdwfEeN6lg0NzEqYOvc2FmKBsKa/ssPRywlJ3HIJombbOUSCFWiw+GkLSU1C+aR
dtYwk97kCpuUE4HPqQ8Mzf7hfIt2qF9PxZUFOHLsILuwe2T4JepNGebjDHu5eHPHyuzDGPJltgZI
TyPYKcy2msro5Wi+ejCMskCZ/Ml1nfQYRrab6ddNoIsIHijAdg9HcPYGUQrFtTdmOOTtZ+Nmlgx+
CEtNHLTJBRpoJbTwbDzJwUpTqhSrs3IF31PyHBqsl0UdBECIy4Ss4rSUdm9Utz44zyOYcjkUBJNm
bf437lugrPN2y+nSvOGiYVf6fOYd2akeVLkxh5HzQVZRqcT7xIiN/S0ffoJd0h4hWitAbNMfPEmL
OtqqGBbGC2w1OioFdEwdoLVvUvewPxTFlQ0y6B49p3g9zjNxdMBa5dXJAZjOpsUM2QKNsVl/qDik
02cQVOmpTsvHFrpbMkILQ+KHFzwHOD9VzKCF+YGSk/0Yf0SHrOB+RU0vpNGJ4qxSa6O9D+gVp9Rd
05PcGrfsgwfi7l9etMkgqqaGFuV6npi4jgSJH4pvM7No4H0/Wxfg3LjJr3o4L20gK/4BFZqvYMA8
1udiyYOmypOdfavkw4VMFcjAJcWr8dR9anhnjKMLokuf9kG67My89TaUh6v1JIXzvUYKNNgD85Sd
7D9bIRuV4sJO5NpUF8WKkeEyJtoBynkwE9zj18QgwpWxNKhRGvy8zyRNEydmJ6Fy/IAUHX9Vx7VQ
m3RjS2eOIoYrbyDPTfDcN1+kHzNkWu+8wz1kHGEAUeNoXksjniyM1piqAoPkmWlZUZ74q31nJd/e
rjd9JxdwHK1bZaxTLQiUSdblLtp9M9+CNHQUtM6yquLc4UpJli20mcavJtsUrWoaTUr+nb8mdk/0
tC1/B/2skqaQH6e94B/eYhjIrEKvfbCAhDojX+2iGFD4f4afz/gW+92tUZwYKIxCGdHgr7XVbqgk
N+6yCOP+plpMDDw9sQ0zPkYZYLcKwl8q9kq92ALW9M+vS5kH/qy4gvVHc8CZA2M5BlJBfIRYe0hG
+2dQKfO/lOyfAV9raro0TValruHRnbeWgIfWSR3J4ZlSqE/ZFW0bAdduGc08cwIOhB+f7T4b2Bf5
hBwxfMZLfoUl3Wgc1VPC21YF2Dr/X8MnzK0RBuhtAGiVMwtDGUDRdt3q+Tclp7ijvmLmypMkJ/xX
xvbX4OLyBLmlExLARFQeq339M9o0CElNna1zBiTh4EkvhJhW8Y6QdjUk7Fq0W/tE+62y5ChS53XL
An3NDVOUsfJ6z/LqS2V9totxXQG6F5HuOk8yLvKIqax1CYvbZaVbDp6EVTdLu3sZu/kJaRHbVPyb
Iqn2vsLQc7avswIgr3R0X5HPmmESJ5ZP6pZhzLEFQSPecDSeZmFJNSWgVQbaymwEa6S/Cb05cg4I
xgEFxdhYzcZJDD7hy5p6h2uJ0Aghzft5W/3w7effzqp8eVXAF3Jaw6PHUPg0PuAyxfNVHFhvTr52
nTZx7QPb4N/wT51LfLEepoIR/ihvc9HslsrwijFxDe768Tap29xFd558fs/8Uag33Ifr1PVnq2oU
BN4jjey3yj7vBCiYw9llYO/NktdzigKQVnn1/Czhj4VxnsdjfR/ikZ3t32pBBjC/af1po+z001EU
kzARravTxCAayRWX3J5k3WMqIpa6y12THUV1mH5aqZC1OBnBBdCu18bt7qNUBMOshyY4oSaA6yqm
IcAI/OlfT/5JfgDzv1ip+G5tIokPdD72Fr4OeJGn0Z8R30WlA1a/g6V7FeqARD93gi0+ep9zdNEi
3BCs0QE8eE+4EZKzlXFbbMlhlBx/A9WNOWoT7VTtVg9TP/OVrV/weUZ6wIo6Z5X1funpgccsosjM
cbrgWFUoOk5EdG91YkFNS1pSQi+n5GLqBJZqfw6Tttzp3siJYUWIe/rKsUEtXFu+d73Ug5HpgdRQ
BfWeZ19oLRPRADQPlcztw1B9+AkJEyQfFg7i8V7sGgWsT1naekPD6TxkYiwqBzgJFACKRrLAXCAJ
kWdLAwqAHuBZFYtTyG9sqKsCYkFX4On3LOrd6i5b+EH31dJWfwhW+YhuIiVaPELlYqGkJQSwAkpY
ZIT44WcIQdCLvVzrwsCx6rpKSYXfLHIpAVGJRayEn1nbc3G5NZ2RN1xYUD8lgDiZZiOB8WPwAfaf
5GNuNg5NADdLXl979xX3q6YHxYBl0NJC1gtMGIYhEZRpyHAK3+SQVGBAYAa0IIYW+1OwPph0vpAd
Kjf6RapWvzlb+VUKCkTzdkZNy+BD5ks58NDoWLpz7Mv1yqsPtI5Mz99G7lh9ozdNXJfKkncWq19b
igSeKODKAOxR8Lj1ZlSUehj1bHGDYYfNzNLBO87PljTsnpIuzTWf2+wCtKse+BSGcV40FNNGCk1D
OcYDOEN/a5pvbysB63q1/CuJcALi4Cwlshte5JX+4150N8L3vSuAp0qIkfjNFDuSQK5UtfnrTifW
t/vAXTmmJiivQicV6ubMfMSR4NJHPuVj05xNB4HMxIZHx4+SQRrFu3VR/SqrdRrxtADJ1PibiPKt
Z0jiVlHM6oUOwrUMVWEKvdge/SIZltulWA3PeYa0vei0LSa5zfYxKaovcsXWwNEBMn1eNI56a/Em
Sev+OKwxQAiwvAk2iN5fW2yYD706VaT6v4ekl2puhJlc+MHGDmX0EqBtKvkGTHGe4rC23y76lKu4
sTKbf3/DKCdZezD8Ipf3bOFDSxeEeiMH0k4L96fYrkMwGhNIoBLK3ERdwmzMii9IZp30cdhUsZKV
lNjD3c4XnynGJjC53pNooqE+0TYaV1SEDWK6MqTIhwp/Y6W+bHMOKLZdhbzLbkQtPgiKhva04R8J
6RHlISvyeGRtQWk76hKbyliBsGYMctz2ZwOtS9XATNSpTThPZKU03HB/gnlX+JWrkGphU4PYVuwl
OEwHno7vqWlrL9VDGDvsBFzlhaZcIqgPcwaHn/HTJS3tmJiwXsJtfMEHW7DnP5NBXMkp8uFqmhJW
Ppspyi1YGv4Dt0gbi0n8qAPAXvNPyUPmMgfO/eBl3vP9gS4lb0e3r3MHNGfuOvcw6T5NH72rozaf
0V+b1YCvlRA/NlUEQAOADlIPD3SbGBI5q4K4wCE7koelrtwCKDYIMeUqv8i2LYqdhytVx8nQ6wAv
CLudk9ALY+8f3vO2vWNPbobLAmYaj+MCVQAflwmizSmy5tcM4LM3pJ0Bmc2FxTjzRnwZqNht7LPx
28d16xmWCaMyN7Uwlg7GbDIf0Nrzq2ucy0DH24zWSIq7dMJW8M5i9DSSNhBwsdq42iD95n9XDOus
BUvvkeyPKBMZT+FzUyouuYx+GBN2viDxdiszrTK093akky+yes0nppMh8nNnqxY/XPXgbcg02CJu
xiic2rwM+/TEGhwuluIusL0uFv+KeTGo+9rgXlPKk+f9Rzw9Iny+9L1gSnHU3UvX89p16t1z/pki
epl6zl1KB/0DQsa3nvNst9u4wyWPUYVnvTfBnSCsbBQJhwUTnahkN7V7SEh3/biuBjh1qF7fmC97
JdQIOJNSiRpCzBooXSCMYqWL/7MXO394XxNX6l3O2p6seSAM+bw8FaGPNYzvuS17M79xFKdwSMpt
r1A/1AsC1/R6JMOWm3TqVbDXOYld6dLW5KUrFCF/2AHL2ERYIBk1XwWEBqgvbmujKn7RLtk/MZro
CSwVgUbeHKtezqhsqEen3TIM1s4mxNrAEC1xtpYQcwQhW/ioIfgjB80R5AvAI0bdoL+hVQsQ1khS
4VPIHEXUFQpfQgGPBbTovWoYozUroh/8d+sQAzUAmlhXW2Pw72Xb+tqpADubS50lEeCfSqjA5+vW
GJQlfg02E0aUnqL+P0Q+nrSVUO3+IvqZTBEstVh+mZyEQsTkgG7toY5OaUqUWcSa4A0d1hdCU0Ez
fm4S61O22zSmFhkgYQfOl/X3RTulLfZHEV+07D56SWBoyJSeCGdrkvkFzCNCDxHXze06XhuW7tY0
84zwXl7J4lFPhJQ5fTKSG6sTFEAucZ6dQQTfwZeIiPsS80oAqIdBRleoL6YJdst0v6Ml2Y5VJyH+
3KYLe64mJF9zq6FsUDRENRIsY7VGn+lmy2xe8vuir+BdzdP8va+Nq4dZ6uBIk4O5z+YHVDg9Eup4
a7HIm7hWdWFvev3p7iq+JqpzyDUrRx8rL6LHkbJfSsFywkKT1hAXB4NVRKYMXb2CU6BH00BZPuD/
15JJoz0/lQZKE8K3U+bNNgA7sRb2zhA12vc6GS/q27XJH5IrF2AE9ZgoFP1+b4HYqEyykV9s2PG6
6jtOnKrzi8byZ0WDl8EQkDz4RKLS0b/LFnP5fMnbaFflKAM3N1oIpk1+O6QtJHF3xaFLGLh6UBMU
6Yul7kKFYGzFUhiCbGzYS9WEcQVqRhEHu0hCGqZYtCkcQ5yNHUqmBCTu1M7JHA7joGQPr3IY4PBK
80KeQbsT9esSmwCudZViGTj/yW6IcprpF0BnX5zIyCc9AzsW/eoyWiUzNJ5Tf0NJFmTboGGhkM4K
27pFLmEYAIbSTJL9KVteCA99/lnH5wWZ1oTmAFxCd3FcKblSmNfgRWeRh6yOuG8QpZ/x18n5bX/4
oYxLDz2+Dm9C+nuNO40KkxbCdBOlVzjsdM1vRrnYbWP7zUNbiJX++bOgi6oCh/uBo1+qLkCRP6Q2
orFQqLuA0m1dV+l/GPHgcv1cZN3wyLnfYF8piYg5/H0zl/ZNKnyRo0DPQ6l4kltrMv/VcMXQqQY/
kPKRZhP6Sa/IPMkpa+itE+Kn+g4Y1Pxm40LOwI7QHyb7slkymtch325M8TxM12ynP9KIupFtqfJc
wESZX032paR2nJMLJrf9Oef+F7pp3U92uZJCEhzLlEb3XTLsir0exUHOehfy4I3Narb57p8mYyE/
kPaDV1WweOvofW6qLU1Z9SAdVDeVq9bfsy1QHeqB1KOFFvanrhMsOHCID1S3eZ3y6M1MUeIdJZOW
n2eh9h0w3nIa3iBE/ZLR2Ew1/8g9xKT0Mn0vTy/0OmEg0ZLB0ydbakFeIWmSZlz7Lenxlqs7Xkq8
jcghAEyNunCG5Hr90lZtRGlxw7t8475zGDX9L3RY78xNhA7Sed+x8mwC5Hbq15PRWMPWxuM6O2y0
BUw2j/PW6aEEHsVP16TxS5/I/b9OTJAwI2g6cY2SEqtme46ricZoRIHYV2h39BMBLANPGjRM1N/n
qRT+BVDfoPWXcUXRZGbOFzqiRz09BQqw3lqWJXHbnglz6WxsW1iu/bh9GBxebyVgwHg0XmkH8vIG
q4NoG6ZGPqL7ls+zPAeRIyRS59vcof30aTA1zZhd1XSYHUr+/KTDYDAHJZydXGic8OqIuRhxm7IX
Qji5HlAh7CWuH0/gXB4EGvjmgNtWAVP3q3GObiDM90ESyh52WLmZCp9oXivSBM0untXkKLdoQ7T4
bEXEzHVibX/eqGiP3e+KWV6BTQVPRC8MPAPLIKmYOFPn5Sxev6lWtcDg5EzMhFkOnXA1ub35Mdct
BmBMf2c8w4lthLsHM84+q5OmSpZvM13csuSJDQ30IhJYidshr+vcDj/2TJzvzcD5Fgn6xRqILYeC
oRB1juFHDctWuZd5BgoPSPC1LdD89H+gl2Q/4MEfFGx1b1Nhyvxw8rJbVzkadMfxMS0Zt4wAmN9X
qauM6yVv0oBwuTr/BaeShgqRqlvktYUAwaaAin+MpcYmWzCeDhfTd7hLkKJR/Cgdv5aoTmidO8Ep
QhGxjsui+/l2dElcwKUKZZRPMqafDyO4c8M9OVDDdgsaNl3KBJ7eylhg10Cm5Tx6C9k8Cw+IY0I1
mBcbVxCWx4JZ0zRJoHdyLhKY2xn/Rj/t+//08r2FUe21fEf3sTU7LAwmd+HoiOPsWAX9+WuIItxC
rOUdu1z+m4RwEKBjWjbKfTIXEp1IQokuVC6e/F6dn5wxRxpb0BmOtVva0qliGz7fPDD5+afxM0fj
lqfkZdPAHoCgvzlohs2SVHrThXs4FKWJmtFSBlwREXd9fsOWPeAWSfNSpmQ5i5hzVsGchB8m1Sn7
CWGtUFx18eI9I1aj+o8ilaQxcEU7aGP4j/71IvFf2Yu6H2W57PG9GVTZJY0YOPumZkWsgkOOM59K
kKRcYOakpHyZbB1a+p/Ok6eHOqSBSnyxWvNSSbEEVsoLmgqhNRiEZhL92+efJEgKLToReiM+jeuT
MmC5tGScXMSVn34BK2msylPyMCtTloiDpMVpzpZ9UAWoT23ykvO+MikbvKhImcLuFumDYZ2/u+GU
cnrelEWeIjO4vhTsn/NtZ8SrgXSqsPG+UTzDwzaA95JjuVSvUuCJzP4FrbouoT1MTV1ho7YPGbsb
HFS9tE5upoFxHytOlPjlLwziyI4QoiKiH8PlkeYNrRDqHtFknE3U9NCldw5PRPjoFknoAl0y8ilc
m27Shp0MNRUod5wvQAA9SBqcTIJY/VXOxfOBaNo2XLLmLtJFCUY2MtIdqdniDJ7Gx5DLvx/j2sTW
QpbNdPxkdHM5DBKEuxgKqoFJUVbvP+Z2Z3A5pZcQmhBwkmN76MNxPYqF2s4Oc9+PBqdUk+0r1yZO
rbHQj6fIYETz0bAeYpQy1sqhUCIph/QrlGpz/JMS1GsFPZGuPXA4IO61SameYeTH0r7+qQ4LpnjL
nVHDL5Gb4CrcSsorQ4HBNiIm3J/Xit7RogCpWpue4ujBzeOODhwG2zXON7veuUpejgiu/mQAqvpR
7dwIm0HG6Tsc4iLemwftqbfY0e65vasrNfCRQiNzUdOVMdjdb22k0OIxU/WM03xXvB48UXDVmOI9
4wpEj4a3Tq+0urlpgMM95gSr7u9L8WQPkAvch+yvflASGMFXSw9K+MmDv5FPfOQCNCcKj8LJ0r4c
nHr/OO0Xp5pqEATIlKenb08h7RpzWXzJIhvL/Q85k3t51NLYONNie9WnutKTcN+YtfZmHNqUUX54
jYQ98/R5lLnNNYSGMhmm3A/AiBxz3vKDPdWuixNVAY/TQ0GENiMglt3N4v8qeTG5xF7QG0ci0SaJ
JhoplHzzPxwjuEu9H2G8s8GluW2EiEiM7ilscDfiAMs7yySoW1HR1pVFw64xaE1i0bH/LWMXdFwS
kGuOqVg6GYugmqkC6K75urJwuR8HxbC4mkXnpodpdk+dOg8rnioARrSoUjjg2B3hO8dqoeNeaf4p
/L1JlmHGX0LPHrQiOaY0zx8Tnj7QB26D3GuOPCZOrzz6Jx9siaPtENhx8AArCepKkyQNYwCMNSPq
LuV3POguiX80w8VeTlMsDk1xJqhbLEfDZt/J0psvpoxSeLHyDVO28C2vucXVoH/7qS/xH/v/u1EE
eJ4/gdeqS+sAI1GRKQH5sfwANRFWdYzcs7sIs1AihiIK5bq0RKVCx8YovNHn8QnEwl913D3z1WcM
XqZNxfgdHwY/7paqJFNiyAB7/XoAe5/fFEv6w2SyfdQDDGR6yIxmdNNfdJ2l3TNxhNkOtD8PPo8L
wBiXMPM3IBQalCjuH69TadPdTd8NPqTIkxBoNGyoseA0wVOcF3ZTqPlPtDEFHQ3zMbfGAMuMsWzM
BTOhcLq0BbSirwOy92Py807queK3WoH9LFaXJKzDtMI5MiF06ztALuVdKU+lnn3AUjIyX+42rZZN
jghyu0f/7vHN41Uo2hOSdqXRWHDxx+s3HuRokoy5rAlIQYotqQyBZ3laSfKEO8wvdO5aRijGS0zg
UvrB9E0WV29mHnqy/MtkYoOvR7GozAIdYs7EdwsxJCbszq8IJJOPPOH1zECQoNBkH3p3pTR60QyO
eBTe/mERO6dSQW/lJsQAVO/dftJha6PzlV0A2ESceAI4Ut0lh8G4kIsP28v034n02xfRrG1gktY0
ss7LkM0CJfsRrmA3W/urarrW6ZnScy/XNY/rqFyvn+zN2mgtjvVIGKJBO6R9Xfaj/c37+FxdDnh5
+BmXh9deSv3vnBrF6WQLCBSFtSVccWCn8hwdz0/Dxn5c6azwxt4jeNM5TPf5Si18zpVfGEcx7nz+
KXgQ6dN7BMpTyR0Lhz3RE61qPfTEZzbXq1P2Bd10iR0wriXVdH4qc3lc/BtBb7+ecK6apxdfvz+L
WI3Fn7A/QeT+3PAjgQZJCNU3NHZYUDyRKeb2912snvQYsi1aHFfnTrDtuJMZLvCyuI7vSgTicFA9
O2Xq6GpURuPhwd8PIVes6yyrVTiziavjGVio2QkDS0XK8pzS/FQ0tIHq7ioXWQadSMsBNKtB2JxU
cXLE4Y4JcRoCw4In5lTyiedZ8mPKI1QliKMyAAn/NrCST9n3Jun8ASOtrShbYHxoQRwdEIUHDSE9
W4gRt6XSdrNWOhz87JrHoCQAx0H0v8es3d1XL2H2XWMA5p1aEWYX/y1ORp+VLgKi6CvbwKCXAUl8
eu7G/nfRW57eV03OAFhi8bgfx6j8tt000kf5jkpwesBqiZomNJz2uSKCXeeJtrTVUGHYLyDTByr7
RoZ/eBfkEA3c0zUHHfzU+B2iaXjd6sohobJ9MNqz4oGrQuS4mQfHwuW+uE1sFKTe5+T8mvPuH+HJ
fEgRp0RF5jpiNLVksK+qbiZF2zMPjANucYAqvDS2zQOdTNefrmODs5RwtS6VjLcEsA0N379cKuIk
N+LX4tS8B/+stGT6E7EpzIcIKkq8y5irTnezJXma/kwCBgDHnEqhM5oMyjvg/80NTUn6xQsOxe0W
QUpzXrxAdGY21CWKnapxIuHBfJnNsBxgVVWQAVixFHF6zcfgp+KYgx256cUwBJ9JLR402BxRoKo5
l3TK25XaNsDWnrXSj0sixgPAREovFJYuygk21+LxAQgQ6rxo6dh7d6yQTRDEsVMO/OQqaW8zdCYo
afYvDRgPpodDmFM1aouQ2JSd63Bp1e1Pv/PoBt/oWwkAhSPqEw0BorFUNWvZl2J1KKoOqxTh8RLv
D91G0UAiGp5l3QYKvMV+82S+j+3/k2suZ5pL3d27Cseq3IHfaSekl5mw+DYS3+N+Sm2mcX2jVy5M
FmHNYqEelwN7QeXjXtdvLEgdQDoxtdNrN3FjBshTMQn6N3o1xEU5gpcRg+PlfKiV95LAB3Inf1xU
j/XvOgjC3vNJs3kP984GR7zGgN/TFIc8ORET1CJ6vztv/0tpTavq39r+eLzmCWFwON5dvQS4qmHb
g7T3sYJMVHmfsu/C+J2LB8726F1lYwtNRTtXxKIFXUoPiwXkcU85EqEXl4MQb9rBpj+9KjIJVqlT
N8aDPmHOMRX0N+LqlpXsz9Pk9DrnW2BanQv+lPvNXUcds08+/2wadT3DrG0suqReXZxWju96WzWV
7nLJfocrEmVWHDzRaXiYrH41dNR5nXSmCaoO+IGKSiGAPF3cewCP54D977YY6hYnxkc7X/Ki5dlQ
O7Et1Oq5wf0d4vq2MneYBSi9aWAFOXN8eQtY3Z35mx7K/Di1RxLKbXv45L4i4OiewJA8O5apxzAq
szQLETx8h4Egna8zovxd+BibSW5jQqnbWddt3RyShKJs0OYych3rr2oL9wBmwLaBzUYHnxNDjiKX
9plUYipPSFFnVlChe22FbCiF3fvyNWSy/8Bp14mbRlSEds0lIEikbAMAE1X15BhTeJM4bpAofjga
qoZZ/m+Ui+jsddTlzbBm9NfZugjfY4eQULvkxTAMeNlZ2EMt8zUVDMpX9uUTnfmPQnMPyMIGbgRo
QKuLPIV27fOvhhLXZw2XIGyBxtHYRYZGhthjDexL8ucC14de/0p9voLKhOdxPR3caM2+f3IEycXx
oZQQ0tzgcgpNNvaUjp2rz7nqI+7gcko1J+XWX0mTm54k22bVU2mGnoEU/xu0kzw0ZPAmBdcrCKFe
qTGw6w2cAUr3i1319Ig8/XKlx+cDg7QNQvsZZ2mZvq+a8dTe9DLZuWjWiuxgFWGQq1RtLM3yK2/h
bZCOr8hpMkFyb+c4f0A6AsS1vRxeMwxkIA+wginEa/1OmvZddY4y/Z288Rndyxq5/vWH3gif5GJd
8bjoWkIWadTc5KFY7Me9vzWumxDTfbvQVi51fpjM/wBKurA+Q6Vp1ZhqactlTyub/n7Gu+hsdZl+
gh3IhpBbN1E/ZupHLsRMfWwk8HjAzsTDa3qQYOngx4jenyLzV5nT9u1QtBTi4GnUbYHm/3TeKtz1
6nCcTC5uX25RjgNluUfYvlLef+LnM367iK88PWc69vRtbr46P0nPHptd7bMyV3sY3WCtU403ZMab
k+9/DrsisVZ3ndciQAhX8Fo5XZzhIaDqGeqpfzzynme3olJuH/GScEGkZ8gwUnwaeQiDHBVd9VMV
qfxufyHeihJm403fjN8bwOpAaw36okCFhS6l8jswh4tSLm+h688ZMMElFhUhEyLKULPiuVj8Ud4Z
+RInWQBx/gy0YkBTfcm0tplxHleXIVs9M+QmrOGoi2zGPpL2Y+A6zY7iDjCvq/d56+RkCnRH1OHr
15gMlKuQn8DozRM/khufdEe3mo3nebnJELs/JepDBpotvLs+66McXpcGxvUO6hrEGhBYYm3IC2e9
RNNVH5kZVdTJIf6RPHh4TigDlOL7BU1AKRhQUNm4AA7cr3gz/XtPv2YCwVq0RiZGh/0MaWfQpvmr
cB2fAWE5fIsSVxVrmv82tw50LdzRLiz6XLCj9GiDBUmcgZGFNvqzGeRFgfb1WkVuQxOoFPhmcqcM
XhP++d4fOUiGrDpVCL5uETerfrU5slhv8K3aSw+3pWBA9AsLXz5osjuoaXavOPUxn4FoBhyZRh4i
4UkrWA3kbXln9O680ddS9f4eewIV7MJOFn+IMXab/MCgJbezxz16OrvlEMdORdPf7xOkbzG/V423
lE9b2d8yF7E9JnMcfHVUEmGR46AB30fS8IN5uxZzQoABme/fNiiuGNUz2wT5roetyx0I0vjtoE7V
Y5atZDnYFWlXlwcxBVHTXhmL8vlR4HI/1a6azmd0c4tNdegMYpzK1WmAV50HhcKXp0HgXBWwYvGb
qI0khCCd2WXpt61QEDUiFa5SvEWeS6NpcXLcq+APNGWLS4x0hVItiVqSs4wZqWl4/iCmNRgJnj0R
T2XDwsktWn66IJs5Dw8ONMeYzYU6Fj7N7LJuWrgBaYziN8F1dxILraLEzjq/FS3QWlRwSgOI//Ha
NgOSaMmAZrKUecqL+UgL6HWMwMz5d8FEvyy+kgbI2sAA2onHue3Dy6OG5wB/FUmkSPg6xpP/dJ4h
v0slA4L+gC9LX/m+kb7QhVAZNRpYN5EomfIfzYlX/pQMqCODqhyDFDxi2x9LdQcIGSyidfrek8Ez
4UM8BRWRvhq9R9Yu9eRw8wIH1cO2u+bUCK9nzObw9bvOagDsmxcrhqV2rih6j25T8VcdhrgWJcc3
YMjFJEHy2h7ovpqHqOuPBGHlErEYli+HQLgql8W1KxAMqJDiRbF+FpVNXvJTh7G8J7Qk5NZ0VPCJ
wkcmSKh+R+CKRtskfRGMkWVH3XCFw/ujfWaxu8AnWK6sWDXNbNmTERnN2NKaLOlPZkg+KBztT3BB
6TwSXgje/CFn1NF6zEAYtmH4qVvhcm4iNAMYlJlHYQC/Jp89Iguiaw3atQMHWTwe2Y3FRpRp46Hf
BKq+FUKXMYHpHLwpWlig2KLFysVXOU6ryFmVtuMRKod7rfjrB6M1HC9U8i+XOKWEV7xaw5PAPwXB
Thtq6qLjbjnnXKnN1gKtv8vtDciakZEekKPA270wKtpTZxNETu+L63mSIt3KOto9hojs8IFQzESE
XxHO48z+jqXIfIes4V39xWV0dOea3EDTUf6ZPufw0CcwrBZIkCK6pxIN+j0SMbHK3pUxMkWDC/d4
qPvKLCeuSoMMTGEpNb5R7yZO7Q1sQAVxMRZGN+ZWD3Ku5Ze1N3jOa38YBTreWwfoTDW0i42f1xXf
iN/2Y/LyIQeXCmWcwZF4IYZ6Css2vCz2QzLEyj39FxMmlxd/iPtp8AIhmPY+iNurpoY8bm4Pn7S/
gtGown6bcsoeyVzVBa0j0PczLZxpM/ESVxrJkM5r7bW7YXiTPh1CnRIUL4EVEMv2EdWRtVjMlD+m
B1hOKvCPsHKEp3D3nuZLGsaBGNRwjKnKsQiyT2Mt9L/b3UPOMUAhYxImKOqs9IM1N3KBojobl/z8
6zuLFxXjuaFLi5cv8H5q+nrb3p9GmUoJyjgAiEQ/QI8+JAh/18PTWlmD9QQPvF5xGvSxkP0d+R22
W2FYzJCFGKebDWq6Zqf01Z5mdB1gItWRg3cx+Nfo6a48+GRt7mjsoXlFBdtDw0f6ZkkSBUx+cWfQ
+OPLmt2QoM6A5g87R/pG0M9dWvEzWB27ptjbQRbxOkiA6P9vamyuVCAq4MP1El7e7mK8t7zvm0uU
5w1nQ4hKOCUt4zCdrijP4KueQ/HNrPvgi8PiD5D5t7zS5wdF9ran2JEgqyOVv69gPHwFgsHEktd2
zCjiFQuLFGMOPoKwpF9BKYDuexLSBqA2WhNm8SbQ2zFFDsmKdvEpVZ2KF/mtXr5oxb4bsp/+Ajb/
D1KrJqZgeg2K2qAIKIoaCQlzbGSLfAPTFhcDaS6TTCq50jxFQ4EDdkYj99tpm4Nd71WAK8r4Yt20
SwuPRcp+9icJOsqssYSvRQQ0DckOX/D0mE6h9oUPfczSq/FPh+oVyQ6D9dLUMqDFE+oG2AGpVx0K
SwRr+Dku3hiu0PlsTS08KSq3t9Gcn21D15aq1kt31/YCWE3BQ+1wCNzWIGXp/cvDVT2EQJ050dQg
hCNk3taaXZyNpqHVQk0lSEZVAvvjtZA/5fV5FpO4ZkQYID0161ptAk76dQOLezU+Gyew5eFqBepg
ZRv4Hm+xslCZ3e3RnmRuDDj2dyVcjNMRIRQjpHG/NXP9jC1OGCaRNiXb11H75zCauDhbCYcDqlTI
4zDSN7RJFAMBXG8H6+DMyl+HghaOjV1wyP6YdcRk/Tv/eZPfwO2uiSzNtPbSM5wHY9her0hyDRb+
nfhrxC7i8+u3Xz0uayTIHHV1gsogCiNQqZeyXc7/neX67/VzKpeJuPzabqzKhFHlfu90JcfowNuZ
d/r0nlkuJKagWjD2tCRIKubqYQjnOJE+Osmsph6tqDbmiVaOv2flvTRE9ti6uQQHMq+zuhuK70Ab
5QzVe7DxqV7KAvPpJtxd5AxNivpHa6MJRJYRSm62uiyxT/N80C6SGzpLKEa7Aeq0ufRyuNGLTFPy
/R3uiXPtxP8SU+yg95FBuUeq6tZHfSiDamDO2YmO7rvqGiKVFl9PLRdkaL89DFXuox/lpYGXXsVF
PM81q9LqO0g8IkbF6Dld6GbvXmKEsZEnZMIlSqXKZ+VnwNE48Fnv+orut19GokYkqseOdAyULTC0
hns4Of/W9SEIfpkZTzQDo+OkOzhdEqgdsGY+S2gfig9r8mqS+Cm6tiyRrd6Hea5398xurNKxQIq2
eFfAYnjWDIKG95e6iUo2F/mp8zlqVEDnvJoPNX1Dc1829/gFRX5e7b/srjEmwdDlzflAaZTD88Ah
FAruHgcbT9Bv/rE8s9zUGJFv/kUf+bH88BfcnbbBO2broI5CHzwizAtK04kPgFwZlw6dTC8nKv/F
iwBz5j9jpeqmkg60iztXVm/TjRFMU92rjKWLcuaQIjSoVuTqpAOAX1z/cPLftthqgv93V5HpFwgR
YSfFHHiPY7Vrgev/UE75iq6biAyQAgd8VqjsANPsqZ7XZ6NpHQqCCg4doQochCA3bSm3GXar6xQ0
PgG/+ptqxPDjWyeOR6LdGnQPO7iub8UT3AwdXhMYldh4VAf7Z9QDWAnkLmTOgXqcn7VBsMWndr7O
g+0op20FOyooVQfg+vVVFePOhDI00UunUApaCfZXa/leOpy+lKsbIGdOUtrB50Pzhd0Ym4baubYk
QZWFhGzU1loJCgB5W72QiomrOHX+6GiyzLEOdRx6BmPTgpc86Jrji52XmFEONirWpmI5bGp78jDu
2hic6dV93zPGUbXiCD2MfGTj7kH/NHKhTNUMViQUjhhV8FbzQhQjJY2DQci7b083VUN4XWyzWObe
kc1STo3w4aIlMe/uEzKxZWIUYF00C/EMIRp87Q4S+ZW3s7Tra7isAqBdfQEW7BS5NwCeHUqWEdUY
+XWL0zekbAO8SUaoe8Kwi2S+LesifIut3Fb+y7DdKUeAWrbRQu+IK5v3AFr2zXLLRUCkgPzeGtGB
l7n4ppavd9vhZliWSAFVuEzDwfGVAzybfqe047ZVyeR0bKFT0rh/M+LtsW8Ft7sU6Cj6z+8u8605
3T4jEo5vHY81kq6cCPC7agwenYyuR1TTFzRuvvuqdNKIgrGLouMJljMXLE+FkssVFuuIvPQ+l8sW
4rghKFd0QW1A37NGZfWq16yEkTFNSWZ5+3+jbl6fQj/aBFpoomB2hLb68WEHyehimrxdUEIrEsxf
nx7rsosqCkTvmY6QI6TpdCvHSXb0aPkzxCVojdJLaHAqsSknjLy2azCg+Gm+WXJYQP7V1e2B7UUX
oJZ51XsQbRuqXbF0y2umqAOPcgq19pmEN9Qmgb6dUtp0WoiwyZAZDWLSQh1mj/4E677McriD9+3w
J5UDs2B6wlvpl14+3Xu3jV+2BwmZz/fEKhlz07y5bPpH1AbbvoKHBWF1N6aa7lf3g5qFPkvX7fq/
xyStcfHsHNzxQHydp3t5cKouaNKNn6mI9L4LlWXNdu4hpHF/SHfK8lWnX9OLxjlft3n34noo4EVV
Y0Xi3fIf6zOWr9uxGVbCPLRvtQ0n61qHQibZbuMpym/Nc3NfKIgUMPc5wCTgQ/GZir+lYxQwSXVG
als4ZGo3d6AUXxdbQn3PlZGzGrAfzjpEhYXNnPaDMWTTTaSdgUleJw/fo6bLfQlDGaa564ZGmURG
dFOPlVU3rCQS87ygmpoPkMZsiDsu2iRTq9GcxDRiDsCNaYUuN6PP5UwVyZOIsqLd3whP6Hh1r5fP
r6WzrU0kaIqNpEtct0Dlh5ChQL7BmEQGBhqTbvGCR3sIzHQ9yeW91P2PH8wad470/wfWMWeP9u/1
7fD0XFFpZQ1pnk5zUB/2mLqjoj3zZcBk5+7MDMamji0hvgwW8TYYc5D/3gWhhOzR/vGF2LbzObQh
9OseuKOXmKgdE7xw5kN1dXuucUDBnThyTwmMreKq7RmrTikbHh1gU23X+xquswpPU2WzIljAN8Io
l+IJ37YskUXtb6ESNCL4CmOgkrk4uOtc0LTATGNAlMCAHv/eV/J1uCUy8yCZScGqaFondBL1axup
c1CfIyajLz/1EuKJprIHrEvzFLpq7WGpC12rQSzmtYcSkISa1/EptegAREDQkCMKEBmuV9ote2el
5t8SmUWNbdBdJdSSgnPNfHc811nGGVnFZLsBWpgU/P9UlHkIe2wUGzXDkYduATGZRTK77Dj0IsXI
XKcC1HV7x/tSHKEzE1Fpl8UX3ga64ithF5mQtmvOED1uzzIZlSmoEc6S2WRKH+sAOuNISmP2vLbk
6rWrADsl1SuDOqCK5xDFm2r4kNC4tTZ1W8DDMHKE1yQU5KgL5qknGVQ+f7kHKa1JjJ1GSZR9Cz83
MPrqNPiaA6wB0+pXQik/QtYzZPBpnZZH5rOrO12yT5JvSR2YAeYKs8S4KxFISHCfGRTJsJRze+0L
i+7VP8ogWKLP0pawqcBdoqP/iuFqkxLe3Z3lafKA5kEmxNGOAP6a06GnCsQ4CpeeJCefNNaTjs7e
5Mt0tghf10ichlPL8YwX2e+yC10g8atpHYbItICXZ/2jRWW6LM2VUA0HfAHhnXYj43ftw6B3iwTr
evu4KjBvY7PIVey9RhLLy7dI+29bRVcHT4ucON0T+HLCnm+IoJLxslH+hPX5iiFoyNPU2Vnk84bo
1/NOAtxJKsIKvq0soQJ4qqWFb1zaeLvo3fp2b/ktyY/iJWIKzdcJ7d/5ebfs4zJmrpoUmes8dJbw
LCJ3en1I0d3X8vZtiIvzrfksgU2BYBZAaQbErtRCir/kszACPt7HMzpo70kr9MEhUOkTkIaW1H6l
CboHl5w8hWJZ1MW8nIsrYxVERxjIz6iQWGsxMYgMEj8uhRzfvJ7ImTZrvUxcl+pWUnh8xjraoWFI
Jox5m73LQLP8dePioM/SN+mTMGgPVh47wMiXQcJtDaP8z/eQuw8yoO5Gc4XrUt2reLUR/1bcv1Fd
shI3XouCowJpfFuZ7PFm9tA5uHPUSc2et9PobNZiDqFfDW+2ourS1Mly+Asy+0Kkeq79pgk2D5sZ
sCF3d6t+ViN2652dTD2TL8hc+qpuv9+x9Lxh2oNSxLwKlxlS1+8xXq8H6PyfB0hICxebUmx63bgh
vNt752JIXk1wSIJdyRADfsA4TInJSGGufCYppRVhXZgeIAY/vtp8RDIuj3jfZwmflCP08kCV4yey
AP/tKZK9GBp+cVG2T1k733S5g0RxeLFLMAN/gkxxwP6r/ir2mxQljAzx74cMOVpIpvyolSaHPE5I
P6c5FTDuIu/M4OMwwa7IcKMeJxMAOSTvyWQ1+cmrlHEDbsTQ14Om88pWFgpXQUwSiBaTXf4TRFDy
cpIbQdZE72ohCQcm7kmlLdHFS3CMnxaxADKBQuJPE3XX9x2bMoGVwfoxVSMyOPFd3ozoGYSh5rTp
1TEmpEusg2GyLjlqzCkhPgFX8FZKq6QeOgOPWMrGi2WW2g+0yj5r+vF5A1myIY7yjiGaYi/dFlPK
p3dGoCq4lRwiuqqOUsTv3V4QSLvTrUPR0QfA2sQXOHuAFDpiODJabGDqzztFdAkU4hR5BZWs299D
2NFBbMtYEzolQBlTrgxlm6kUN5vnzseXdr0DKp3YOPZTnBZKm9xqy4XUDKQC37L9tNJewX+iPppV
Mkd94DxefB/hNvdr8gbSkO9uKZK17cBYab9HdBbhi/gti8Evwhi+VqlQbmrb56jAkGwxzngiB6EA
HktuzBCcQQ1MpM2WIRZJGj6kE7v1TFeQsbuuUry5JvJdxbHDPS8jEmvfZRFnXdMMSEXzL/J6ecpC
SyiKbuNTEh4vBUcf/efdLuProFOVnCqyXsuzpbMgaf9g2o4T+c/yyZvy9HOvLhK0y+zmVifjecfj
ATFlBILiyZI7oCDHJfdbROQqZhjK93bx09JUHfpZaea/O3GiJjAKgzcSm3SzSLZdjQlfDpUL5y5X
ceKqqT0G2lw3G2V+hOiL/uXaVMTFM5QxARcpUTClYfgaMDHWL75AoIUUM0HZEN1j8qDhrsrGl8QF
0miVjkY2yG/JvyM+ES3eyrSGwpKRqaQEuK2FsEVZz8Ug/n5NWEJl/oq5B+rfd6vIs6y3A0ZxFkJK
t1AQ3WarkGZgpTi16r5S4udXlaabhgetHK1USHD/tQuYopQXLSa9p45+Xu+cvVjr+GDpAdhnKkAU
MBvT4+F+n3fOxmi3Hb6NeodfcVI35D16LEiHa+1isfeux6gAiHQB4M3HrQd5SvOTdKi27jmtw8ZU
eKy+8n0YRKd6jR6MGNTglKGW+Nt9QE2uEBR30vVpKXz4alIFjJJM8p7W7nZ4qx+OomWan8ZHLf76
XTfz1z9ntsAaT5vQp1zcjGXfWWYNubWQUhAf5VpltryWRwPd0YgpOSugmYG+MazAnIyrgm1fK24v
CPEx7oPkd4IYz6NTI/E/Wu5BrpfMv2EvtFOi7PVQyh8xhYIGNBsQ+k3CnHAqeP+daRSm9k9unuIe
e8mCKzSudiJ3lK5Nx+Pd1dP4Bhzvag0foUueZOALNijsXU/2/kXavnGhgfVWdS6Smt36ButfQnx2
/Dk+1loxpTM/wmRCJ9j+G8Ke85bb7lvVCu7cA+zVkl8LLsjfK4CC8NbJO1m9Fw6EqkR/gKZh8GwV
kztTYLHmgIMnmibWp6EprCBMexNFimrxYtXshPpCis/VzFgU1VxxtlONGxklarFGGeXFia+LU9Eb
1r7lUlFCS7AVQ4m3dq/MhoG0Ci1yK5LMBuxQGxlNhe8Uvhohkp8Qt0sa5ZLUM8x5/oJopONL2mrp
LL/INpBqmK1Y7le0qMg0rJi4IWcDuVXQeuH1PHTWaugmdNCiMmpRU8t543HYDUFCHlDly1lo+laP
1gqOBRthvgjVIR+I6R06hZ5QtOMeA51WoXDK74GKUVPeqTfwLRAGyuWrL2wC8gesZNdNVOPlNIXP
2AHl5seygUp4exTciensklmiW7Yw51AmNhgZaEVjZz1Byc0IUR7VXzgvAm5EMXfZhn6d5FRKvoxK
d4I/vNJvZhsgeXVPQkTlQuVbfH/fO2ufbs1WYW64n2M38WycxykmlCN9dwpNYLxBIWp18T3VH+nQ
v4BlmeEWFKQMzteT+PvqHrwwaUYWv034mHdx+V5E6wV/TgcaIb5RY7TM9jUf49UwfgFeKT08ZDVj
fdZGdP1srqFJt3HUBFdA7CFmEze+A8vhAM3EGu7HjYVIuwXVV4Y9cRP1lW+qH3XYdJiAdAUZuQpu
ByA1zqZBNwaC2xP9YMIyOumL8F7Z7KCFpTjYz/xEHbn9/0nKpHuZtslXCFtOsOloWo5FC33Rt3zF
Hy6mj2kOmi4lbACAUPcAUn82qB77ZAsIiy8PsnBccXIjBSWcSJkOd1JzkMQC+nivZjscfMu61kEL
+BWi+N21R9gzf5s+nLWZXBSawP2n8UEtUPWfvpUPm/tCxYpAjf9Geb9jj7d8Mj29sX8J7SYcjq8Q
KVjBzA4XOMoyBhRxDxidIKCTcyUqbMh6vcPr8W1jSsQopvkzL9yfioXuphdfH5slF7XXoQ3s1MFG
D+n2MJynuvrVw1ZJ1VArDteKleCitka8Ny2mK0QlEmbTWxBTNDrvG+qz1KHODJPk7z5gry2LhkCT
jPWEqtVbBzQzzME4Gd9c8FIFQQxaeqUkVjw4rJtvqRXhE23gnZ4kq9umudKwCiNcnhh1uvEeokub
N6wVX8fPMsIkL2ThNvaX1faloy6oBHFUFlEra4UPXNDr8M/TRWOOhpaERjsDh19Cd1eehSe6zzY6
cEw0hq740gQ98PsIW2LC98IaLiHbZnbRc7QHXvCebyjRt98kmLyWbmQV787nbBSvKqAiCaVZFVEO
l+it6gNO132/7LY+zuZ7PeQxmw6/CsVFoPb/423nuxf+4JEv2pVSNzwx1iNq/pZougIAKHmfpjDO
jLRZ7SxFzWwe/R8G6JD9gofOklEIfb2CP0KCVK3YGk8xt5YIx73dGrVW0d9t2Pol0tVBwVk6vjsi
ZCv57w4hiDgz2jVVZuavdvP9AghKy1og86kgGOd1Rwr7O5UrQ7V6GVwghILXUhj2XIr7ZM6vPapm
ocbw8FfChZ/dWUkNNn2Uncn0fnliedCHGLr2ZZ7AXTvu7xvV5HJmQXp8EKA3FqnAXOgn8ChLyUQh
PcHO2hrA5c0o+HY7ZXXEw1/k4QJ7enc61QdJc0RmU0suPUWeTLt8O59ZBOEazdVPqdgP1EIMdBDe
Yvhn2IsMnxUwONtCfZv41RPd0rim2E4o8Bf6N9Sxs20N3T/0qb0rL9uYqhoo9lfTvKjOmW3dIJaW
3t9rfCKOhC8WKu+EiqYsz1/Jz3v5m2VHBpV7lNamaBNZbZyWtv6cjj6mcJnDhkXzEqTIFmSycj7q
1ScODfbw3sc3vjW7e5fBIJMQyn8hLuxy52oHqk606hiHy203iZch7Fn6F6Z9PejCfPywoMdfOFcx
1Eg2+JbkBbvwVpLbNxPFlWh2QRJ3oP0bMgpPNejRlLlkNaq0C0EYUgbhQxeciwcqoIbBJ5H2Y5T/
zf4e8Gxv/2ASSxTzXd7bz3nZk8rrnBFybUX/6X4jXqf/HoEmIdGTP8rmH7IN4NCE1Kr/NBTIxCwq
Gk7BmnHcNKplXobN4Z61ov0OqbT1nThhM00Uza7DZFhJuVdK9Ie5ffmRqJIZUcRTXUxZnm44PLzx
eEVc4iQUzqGS23qO/ZIHsyB8MQTGX8sEDK8UBr4Kfkp5McgpuyUFyeGL7kFicZLINS1s0JDPb2VH
W1DFjFfyYI5L0OHLmET4dV8ONVwouPQnkJMbYR+NQy8O3zl+mWte6intqoftMR2CmRdHLX1trK4l
n56vlS0lB4aBpx8/omJM0R1aNDtE1kRFEgZAJwAb8cx5c2QhzJe0MHLnY5GZH1ft8wolCu1TzckZ
cxBbGg2dQFKVC1Q0ZHEUo5gpLucwII+CEu041F3+cfANA26XpUsdyqIAVdq5PaFHUYspqnmXQmqY
A+go4PON1Z/wmXor/n6Nk2l+QBfmcn60pAVSOUtFrQYRwEK+ZI8PQdEOrGN67/TvkA9XFq+DPnWl
hXu9flBvi6e0bMK4LOKg+2fZK7KGiRiCLpbhCz5HQFOI9B1ZNE3Ow/faG+5BrNm7cGGqwZOeq8CC
b2J4Td7Fe6SmITjEKKLw/BNn6hhwZhNaN3rwbQPLKljbMQeAkrz8yguOfVHapXfQjWM0hv60jj/4
jrSkyU1lTgk8KDQYSUUJ/Oh+lo3To44nHOrP4Sa4qNOOa2bE3zfvqP10r4akUYB/HxcJ5CW0Wzuu
Qn5OqT8KBBWVRG0U5J+XK23whqh/vvecfL1I0fncuh968euCQiv3mi7FAGZZe5HLRCR1cBItNPRQ
eO2qPbRSsqVjjmdHMPLNQLFy3cIHt6mzFDggGfKd5ITGIP0a/8m6+M59dt0rOJWj1pu5+2YmLlDK
qMpDD71hc4SaQLmE0+xDmf9/6QXpjJAzNTrIl0vseb1BMQ1tJD3xueAWDMYD/menTJS7455Pq1cE
Az7a51z24yRbcut7X7pIK+BseNqzBRhiXXDBqRYS4iM+BbVnb0+y+vnGvpMQaZePSSQQq+wUMtS9
F/1CrG0500jUmBRtniKeCt6GzUDJPfeqFlMVYepoONp3Jr3cMOanPIQU9I2dxddVMoNXCxNvww1S
leuBY+9byS5nYTCqPPv0gcOcwIl7H2P+K0LoTuPD6O1lmt7Z9LOgiznM57J/Cl7TTGPyAp3lrRDI
GoLdNzdTbHhtL7Tof90Yni7Lj0KUY9lXsCFp28tVcCn20l0cRLp0DT10Ier9yFJJEbidU6iQnT1J
zsedIE+NZoqdxOk6XG/u4H2L7025hZNrle9m/TPCeQPnofusifzjtXQ0ZCvJNHiV/s+bqMwBNNrH
ELTlXXSiHnCXrLqhtAUomCXOv70mNy2ZM5AujzJ+E5xrw6SJZnNQkMv387oWbWozyjLqdAWmLE7g
Yg+oeNzJUcogHH11LmtqNaSrNjSfARCNYHoZREukH5gwL6zVV48GTOKz2HWMcFQ1jVT9tTCsAzPq
eJgPv/E2/excEry/6meZWydcz/6gfP8NEiB1o+nAr/4GGrRMLXPPAa3gFqUg+JVCNyDYLIAft6WF
qSV1090ekF51Nq/7LHGy4X1pu97bxdITj0QZmSTWc5P0Mwl4H9CrS7YDbzevWmEo5TLe2uFZptPe
4cXTnScuePfYhNtVykVwRAdcKkNzfiWl504c1IunI6HbB++z0Lo56Tu9u/ZNV7CCHDiLFkHJfloJ
Ho4z5euBefGx3V5OqprReRJY1ZiqIOZJQcvpIrnr+1TKFuv3d0ZKPY8SDwR1ITd+Z+wv5lg56Y7k
BHuUjqXNNupbj3QpPP74n9WLbMa1VGer1Jx4K2IAwyY0rc7gG3a/Ip36DW9lxkRdZJrzrVqUCG/v
DSjv0Z+/vy04l0VA+oG2S5Zf+rDBdYxn+soKtQJ+5m+d4PpaRcBGNfe02bVpOHthMlbm6ZV1ZoT6
s/+AyZ3erN79e+cgFvkIT/Sx/QZho+YNe/CZOxEkOfxr3JZnfXQBWZ0Ju7ECjbRlWND2iGHELoqM
0yifeFgjYIRIVk0aFr4KmEiOobCsbYyavxtL+M1LpasugcjCUkymVp2IbSZfRLp0k1jzO5xJRgZ+
5i5IVK64D7GOoaeRFurNdD93uHEGydCf2u5MxcW00FKzDQHc4YoyWoefqjZpOCvK7nDe95W+9g1c
cCuAjyrKIg3/5vUvIAJf13QcSBd15HDJyGmp/BsMFhcasD8Xizo+1qievT0V7oiXlNuufnUOO6SJ
l5XWL+W5DIsUSZ9uBquJEw2MFAwhfeBHpf5W482+sMG6PMX+bPE4r/UiABHP78VBhO0I2Ap11G50
8jGmmU1IzQ5ReW2fV29V2nLO+nXgc4GBZT9Q9O3CQ0BxDx/3VtrmKp/lVTtGWbhr/GbfNMvTe6Fs
wQXoHP7UPcoscgFCn43i5jJ4As44L+I56BV8SnHnij7XuL5laxcc1YVyPP+oU/l6QyoUdqAqbzj2
ENPLJhTMUeTQnNcFkL0EgjyXd4ldnYIIyvJMYq2tQmefcXU7URqzHCZCXfPRZ19ilC3e+zrMpZiq
Um82rQW16ag9hHzz8pUdhdLCnqzmjvUimSvDkMinnDqpy9kp6RLAxYdl+fhEW4Z7Xyc6hKQIPrxG
PhNTk9Ly0p+8mRv40VB1L891UvOh290jCfgSJGhnZnaBnjXhGtglPCEzH1rI7lPFuHVyU/Y71/Yi
K/nXMwf2eZY9LDkvLgrYUuVBD9neveMnvoTGbcM3mjy1eaBMj19Kf4F/kg+YbaeDwuNlTOoSAOj9
MdP1JkjzVJPu1KrD8C5/VvKXXCMM3UL2hLn7cG0Hru8Pp8JiaAtl72hJLu4RCCof+dBf9SyY81Ml
Eg33WLWRQN1rwC4l9wwloDiCUfDEZYeMaZEtqpOJuZD5UdRK/Rfl9tlLemgx25Hh72xsKRBfFy6q
aWCM5ZcTNU0GF4G++iQNsliF675tRWAgamlRYdkYmBiYZ9B6p1iO1iagXqJWKQ+RukJ12QZkmb5I
stBI41oqI1DsKMvym3LvZMxrgV2/3tPIgkMjm9iobCEBSZNmDW96gLccHwPCL1w5X3p+IyGxf+MC
5UJO5QmCFDAL4v8qe+hJxeWKN/LPqA/xEBBrtiPbOKJt/Xv3kvHlR0A0gRKpkDDel8+uMXdtnW7e
7/2JoXmQmMpTAZYkYI9S4e5mV3jtFyDqs5APyjoYQj3iusEv0InWSILptbCf5ZgyOaGHkD9KSdFq
ZGA813C7qtXPfR7DcmgksYaLpHpx1bhexerpwNIeJ5Zi3zoAG9adFmrPDeo3lwLwPbba5gJvKop+
/yEUWwsHZlPLkRiF4QKqJg26rqlQkHJcNwftw9Fy4npbbhTDAcKNekuY+beFpMOhlH9VJBdX30LU
BhuvdCNoYaQrpca/D/WlZIE6bRrLGY9uI2bX7O4syW9Daee4xV3SgSXyIpAdzBF1uVJGKsRiPEWE
ZGZptXXeqtQAi0CaAGoCIG9BDw6QD7gR1HppdBhdfXWKK5qGc+IGx5d3Eio/qXhmEsrZd2Zzllbn
PLtuJSi7JX9Lx6mrwKgNODdFewLmyc71IpoFnHMK7ELpJdbMFOaCijlYnMoQ5m7soE11J/dAHZYh
lAyk4VjOgjYj7jY6rxTJqQoym3yaY7grhwnWW6RoYCtl6X62CyXzQxny5c3G+8X8Gk+flXkuZLOG
DglvaCNWnuHpI5F6oVA/WyjQWMsYWHTsZMFxvxAQUr6dkOguevJIxhpXDEyW3RyMchFAvZqmyXLL
s2uPOmTylKLWad6YkYrNgxQtpUVTK7cgHYbrJ2K9QMish8HArf1pS06wxfohU8O9c0/iSB5SpQqs
GFT7X0mxX8t3FPjT0pTLENmmTkLAdIFc08lSsxFiqOHUXI+PzpThK4Yev/1rDtg40lG01Ji8s+Tt
crDrVgHpvcL2pq5ESfTa2kMeZLOTq5e7E86mXK9nb10Ks000GSsyYNbcd6dWKg03b017id88c59v
ApOLMlp8ooMDx/1mbRYYtCLOyeXQ7yEXD1FSsQqQkPUKTym6BYuEvLtdIxgpgIbwURCPQhEK2PPn
1PDBTT0griv2CWNEKiJ7EcarcR4xJy7SxL0TLdI/ysPhYEzIINv7hNHqOFa8mKqCI9YI6LEYvmtR
jgwXH8dAXY+1xEtdotQo8AmGyT8etE5PTghgpN37iEGCuA0XY3XRaPQX4d4KGOkOk3DsFnelv2EP
d3qRB1Gsgbdq7VkckTUmTw0oZ1xTUInhWZtj0zy+0JdafWju6rolqMA/Z2MD+dJDl0TFgBHpfuWl
cXbmR04FGktASz1iLKFZwCqNeEa8shOH9V7WVMm975ji7U015yLz+RGRGHAVA36R+T1ycZXO0tLo
sfPkE3O3xGWKZUu07eh/YF8fVCfXY7vs3CY5B0U329MMzUayT4cnv9k/bkcN9gwLOdtStKk2cMzH
mWNKP1PQ0fs3iPVPd/J6OnrV4gPc23ixBvpNTVGxK6YuMLQ1kCefQWT7AP4N4dnttDmkX7iVSbqn
laM7fzNVa1YF8zSm+8PFJyQev93nj85vHCo9hH3I/IISwunE8jeiyMmDXW7XpGUlUFzBKhL+3Ne3
6NGTSXiF2zmTgq1imdMluScdwrm05D/m7yNjSLKmhSc+F2r8JTks8S/nOUCwiwZvzVeLRmM7Lt1s
wM8T71wy9yKADmaE/WpPc+LYzICFxZfMzfkoklA/7C+Q3PFcPi5ZlrvePFyN2qt+givT+lDYIvhZ
IVGyZoN/4qu0QLIebS6JS2YI2mJ8k35D+M7+6+B50PFfF5xw6nz2QGWKyqUi/EZ7FZKA3aVqO2W4
P14TTPQR1Hy2QWCIMxpeJMUco5mXMvbAVQ125jYInJwAU5j6ybzlVWH3v74dnV2C7GfGVDqK5K/g
F1/g/Fz/zEQ5SoUvVcTLTkGDxEOzY2/KBD/UNAO0NbOu80kTJMPqHdXHMtBc5FN4UIV+hqTazT/f
NvFsTqiPudqmUDGdSOB3PIce0/bNn9my7YOHplC1owcVBbwLgK+3CrhIEZtSkFbnRpaDZVWNKEcD
gFmPQ09Xs7BNdzHblXAwIi1zaYW6yGc4Sir/FoDb/XZvYsK/Niy491ecPbk3Z7vV22mb/dCpuFdL
M5SBic2vY1IWONDG/KlU/TCaDP/7cDghyfiPfOfYKQgEUUPO6lUZYhhSEQ80fe7i/apl82ltUuOK
13U8yt2RdSqBD4ywVJgwv49TFDVC5BsFw20XLjRWpbhG+J0hcheHE/eelkndT8Vv3btcInhpwCsd
fKuN1WlDotkug+0M3sNXShi5fX8gVFutYDoQRikwgCGhbW/VHX+EuTGgGjzR3oyJ32/QPrQn6wLK
dgW9H7Wwfr8DRbNGfvQ1FfmF7HWR6iW+OWTIqZHjqMN4ByQk/eYes/O2/O21Habzf4gdClaMIxyC
lEY6wVEBqGZVQgLOBCPsijZEm8Ye1EQLyk0gdEOJh9e4mX+AcEjbO7TRkRHWUPnmIQ0S/3iHh7oj
SNAb87+9yhKlTFtirfk/ZW9Q31V6kbIZ4XmoVWGVzy3LEJXsObhWo7LFAtscBnusMU9YyUdvXeTw
oQ0dBkbe51QCj/bD4eubL6rdoFT9rxraIx2uv7dGpJQz0VHxaQjpb/M7EPd2C91NVzJ5SL0JIpyu
MpBNRa5JlUW8rUasel88w0wnkzywde8tSaP1cGBfffkWIlkYBco54tBsukg1ZctcVT/TsuM55mXF
4Qt6Kj/W71TPYnymg/T/Bs/IppeBwTYDXzCPDSv9jay9tmoiYKuvWyrR/KjjOzyUvXBoBa8h9eq1
SZ7yaYo2YZG5k95ZsguTBQ2iq1fyEOj0FgNdeXGI0cJxSsy3w7RECuFoEb8CKBthwG3Vb7jAfvS/
YLew+cKF/yj2rSj9EDBjVQ01KQ1ZiMVydmOi/3RGqdVI2m3xBD1rDl4DeJeIbH9W9czgQT3SVnMi
QRRTtZn4Ipxt39R0IDE04f3DY8wzpxqAfRVA5KpvIUt9gwUaI43ZxwxCIO7ZhcOAVq+IcqAIo/yo
5qMJ9w22Jp5opsbbL5hrf7xtbtyOCGN0CBDeubzEQFa0Tyl27+B+sx5SuSBqgo7XEACqncEfCKgr
y7nj2bquqAaSTwg7yularlYRvXeYVRhLNnmD68OLiyialC6e4KBL3zDZL9+ei9f53jf17IV5HiQJ
24Hu5MkMek0sEpsOtUaW0+ERGSUhj0PrHuRzVy7HQQz7ENWxca8mD1ZWSI0YmAkOrWOlxQ4Sbrnp
SKvnZEdc1HUDPq4rtOFYT9LOKKAuGTpn8X9Ra73ZrQxAYMcBdn7A9b8ojQYGfko0kyqQ66kPOWqd
5899EstXjYBAGZwx13Jkq3h0LZyEvc0MV3vVttTnUwqzUGXqlDf93BmgK4UiMBnRjCDT5wuxSRJn
oWHNFg4o+9+i3g1ZWtO8PuoNnNFOaS6JBr6qFvuVlU+qqKhY/OlS5hhSDwCbUPVmKZp56Xo81AWm
8M58wyrUAZS/c751gqUGcK5TS2vT6LvOhU+75b8O9gYoy1g6vBhR/hGPSikuFRhdgNKplALXkiFK
spupzc2FjJodUlEFz+RCISfs2AJ0uxXuBb4ByvrqiimgZ5FaflsuPCWThwRMCYGSwl87I4VOW/EQ
eHK9yHW4EB5tYgB5p8X4f+Zfi6DvX7asd2MIUu10BiMZq2rWP/U5Y3WLmpZK8j412VLu1NlpRcUp
3UjMTe0uUnKAMWVoSImAsSCe12xMaXr6wx3H/QIJmpqbwSJLicmWCcCSjoj6KqHmohNTGkmBfNO1
/5AzDSQzoNjzR8Dn5eqXRLR22Ehq8jUO0iCd9oVweDnghHcsS+d/VnN1CHVGhP4cV1a4lCQ8tHct
5yXKy94zzSrH7bqQbIFqiPODtCD1SKOJUTRNV5eOQTJCcOMxwo9Vfk0oTTXGxIeXDgvZNaw5GKJR
PSpUn1F6QhD+CMoWZ5TMCl+6uv+FH1RxnvfsWkJjIngniydZSZ+5UxM007/GsxQcSbqLZZg5LgkM
JV/5c/BTXjx6G+KLDz6yNSGEc6ayu7eSbFbEkUeJhMuapSs7rGf5VyypiNonx1THj5w0Uh3wA9HR
cEKNE/+UJ/AdklHjSbzzo/lawf4WB9G+TuamMp/ANBHX+5q3a9CJ7F+/7dG0X1rCwFvxNuTdTmZi
TpY2Zez/K7/ax0j2bsHsl7Tj/5x6VDG2CC3r0V1tOkjQ7ANu/5sn7tQfHTnfaRU9g+GRZRyoK2Ei
fNGO1Iz+hIKI3Cj3bVk6xqYruWjziRq01i+CJ6j1k6Rwe97sDA3PFIlHiufbOoJqAfLD6w8b76iT
o/aHs1WdFUjCj2DR5+ykTqI3gfZwIwQyxvYki65nePiX8/FBhec/nQpquY5Expb2vzSXjzB0LtWv
LO9B21W2itnabLwOrBsBLCNVMNXhiPugi6zmjlBtssDUBO+mFd6piu/jQAeCVzYpcNn2dK8l4CAn
Zf4xZOR/kiYLgH9bdNl8r/r/BaMOXnEcJEmiktH2mzkkhL8Gez+kpTZkAug2zhgOyNR2S89U5fOy
aazul3ibQnBc+7snIoVnqEcnfg4NulvBTby9bIi8SbN2rE6l9nF2KMS8DZFl/tWRBNCV/0+n0UfF
CJd25fNGL+5C1oiDMDWIydsydFsdh/o1LfR3W7cTjG7HBlqaRTEPfmfZYdrzio6EgzzjcpK4+YGS
9GyOXoG/Tn0qlVda2qxKNrp3RtY79TNi3h3YL5fscWO2MEsaO7lX6TKT8MtK69KlgwwaLhQjG224
b654vrq15iKXLwMLAQRjE4FDx8xqxxreH7s67R30sen8mS/yX66rZ/EQfCVBsbMgzvtkujTQYlHM
rOsIJSBPJ8NYOR/WWWvCyDYWcDX2FnbtexSEAYcNMRgkZ5KmjavurtoGo3+rwnAFLTfav36YsmZv
7e7e7lNDqvR63peK+mfpLwSgpuk095gfd3llIqiGRuAKONOFOFLOHU8QzSHUDNmNA3XlI++jDisI
9IWiiXjfYceMz0FoUZP6qXT234n0dw+zBeUFb7vaFQtfc8TldakznnRMyy9inLYI5AoCLPNmrq6T
wNIV0wvyMdDUedpAxJ4fQHjsCeBzRnp3MnndPviiWw4b+r6g0hvvRarbbsmgfJphXC9g/v1LnJBT
oJ0wP//Om9fdGfNnR76oTqyhO0ObeRQSuki3ZkwdhQ9LBGKRdyzbybaHjwjjlPRuU5VpwryWeIXT
X2zYZFjdo5lPWtSsp6PmM+aHml3fpvmwHEwwvE8E/CSoMPUcgXAci8HVYsXMIkJdBt84vFek99go
47Y4qpsG6TAJJq34Jwbwqk5KofshsJZ3v7TsyuOIryubDkn9CyoBogu7R005D1LDveQDy1hcK+tk
IUTUhViYXTCEK03WQaI1ps/z+tj1NJbijuqfeudu42Glq18owamTlXOs2A0uxw+iSpCuZvUdNndb
MtNHKEVPreHwhf0xZnxwxqqnoxT0RF7uYqpeWMAdBaF1CTkufcRon5CCIQ6mT/6pAKgm+BNncSDp
bMcTQIgC89pmMTvm+QV/Ba/uG+MChRXFZ4LtdEQDgSGNZaheAGmcQ5nLbFr4ZhKHVHMYiw+LANyN
DGuoG/w7t1AcIa4+WiFv4FcTHa/8X6JFfBWUKxeXZSf9IRrajLsqN84PWVUM0h/D9bzyo9VMAZ0f
mONR1alSa9DPKte+UIa+rNVAMpnp4biSkelyDODn7H6lwcw/rTA91nVpFQh2hD+Jh8O7OBdTZAHB
mHEzGJSABeiD1BOWXRfg+izEVXdxFDk0bW6WC6HAbnRmY30ZrgFuJYSkIzFTB6vzhYf9o/6vDbIp
LX7SGHVI25IvV5W0zftRaN3/XFEDyMZQJJ3HagCFRd5jgj8OzQ3iUHqLa3KibgjAUZp2lmy9NlUN
mixX59BNrQlNqYcjmbswlgxhdGe+cJS1SvbjdzRrFB8EC+rpl/m1lEfCCc7p1r43qcTCUF4upGt4
b1YYAZ2e/llKdkzKzpS3a3sF76Kp29eMEp9J0m/3EDmieOxGc118ZUvEcsQHogZVZMojwy3Y2MO0
Z6HQq8OqcIQBFXyjZPbLZRYi56bROYW2qJlD1xC4ufPQcE1zlnBjXQ3ApwudK/UgnvLKFlwPsaBa
8pKHKif1y87CHu5sC29Tz4Ed2t+i26A19vUg09W/YSOWkLd0fjn1rluzMWhF3QO7XQ80KfQrC19m
7+MPj4tyJqBEyG4rnqBUHzXKRD11IeUEJDi071+exEa7Um1Ko/KASo0RiwVtyHT3qSzhs/tgzaMt
Ii3FQE+SnXxVpzhZCXRAd90ZsZv64c6ehf31pXTiyUEBzWkfqiir/QuoKED1TIkD6qKEQN2MTg3G
P5/qqhoagQM8HTl+ZoqcF7xIy5i0xKv1bIc3Pxs+gCq+14rI3UzsUqnHiQUeZmuxBcs94Rfzh/sx
D/0lxOWj9Sy++hUEtJTokq4W1yyMzTO3Y0qmJtYRQaOg9L8/ftS7X/TgPZv4i4oDVNy/m3xGoMri
rVBxuP/2MqzRLlIQuMRZbOsqdCUfw29iAYl2IVNVFGUHsTqBAYLB1iY7oL53Cd0tVmQIC5/BUqoF
ms2gQhO0xshGQNQMCCA6SVi386ggAWeIb9IQkJvX+P8lcRhWevlSjVkL1Um+W9ubzjtHF+fkUHtb
pP1Wbst66q8kbrsTk1d916t8PArImVxNwdVxVycKboh+nw3cJSHFq3iK2+IlT8fhWZxg4Yu9oAgq
zWrOuoWik1GJJ+j2i6we2SbNWgVyNXpsySLqdi06Y76rbp8L5POFDOhgfd1MzoxQd99342Xrq9jv
Ft1OGtrNCAjEa2V8KMJSPY4IZyWSlqBrRrgar7XDu7C16K7NaIXVaxZJrGq6f144mVJBQYIw9fbc
Vt245YRSy98rAhcoUJQ+CduktkWZ5JmdCChR5xNdsf6A6hCsxGexRUM5voVYEft4TYsQCXfWjXRL
cmHH4Bq1lseSoVq7kJkgSqETWfVnhMbIJ4rCgDQn84hect/0weSOU8AmGzduPcY6PgtQd9bWdw7b
FmNOWjupr1LCerP3gPOQfbqnbMQ0YlFBfZUWp/R8Yehfuu8sdl+WXC5llI2gB+O7jql4Q3t1R+as
37TKHJVkclYCk0RfmdwfjuRmJbNUV3YS8yJb4pidopaK6FLv6ztEFPO/moVqkMEO0aeur8aTb5n2
8fRuYfgstLPe4i86PbswzMSIRGAaDnHnmEmoGR4pZWlM06vqI55YpixcusvkRey4UFBmVOlPLJr+
uJp6vTuBMTF91V7lztXQrbdGeYyx1O9dqGrcIVq9dn3wj6xgQDRPmjGUYQQk2pYAXV+1Heba/+4I
jMiKDoz2Up53bX/vuwOuW4C/W7cbroCwDw5ZSYEsdlPizm27MyyKDES2NSXHRm6jFwSU3sK8GOqo
APP5BjZ6yRgBPfK9tIU+wKgPWCMFl6/KaMxqJjwUgRIeOzszvL7gA45YNiL5+becr/pMkuOcBt7j
DgeTgTEoiuwB8suPLxFJ3PFWDQ2xeOhdHWn/Wnhwkr0T0ksI/XPtwZlUN2g39w5r0zPtXv84qafV
LSGWrReZzyR58D6zmUoqSXPSVqieXkTLB27HqjeQTn8zQcLmzizkFJz0NQlZLSZShyRhClmhWsz7
JtPPaCvEqpI1LYi7O+PBqAIf+OcfyYedhdGB7o2+OWZV2+kXal9u1xod1H1muVaaTFtKbsDjwqn3
EdxdQt0XaLmSxoc4R9HX1EyvjO5Bi/AaWZQQs94gEVH7ZoNKHL+3leBKG28bYUC7bVjvuO1NR13O
J24r9f2kMR+tMZ9L3t+3w4P0kgb84hYXMBRfM3QLCLZuFkN+gZm8zynImdyaFr6b6CINXceEboVW
CovRyFDMxVU9cbNJWCFKsxKCbOph7vrZPkjazXR33DsBxXKSnxobCScTViTFQUx8Wahddx6NJ/28
Ttr/m76oI/C5LA0mxytvH/f3wVg7Vi8NcdVym/3mkfi1eFRtBDgIwyFn19dvot4aFMicZF+E7QR6
ur97x5KtnfQN7Mx2Cp6eq3xX0p2YMjQAPyY7zgh0IZ3o2PRA9hw4K2p4wXM378dqwRUxqTgA1W4e
KmqPbuY5X4ljna1nQbgztdCGwC9gjeavqsUnSlqWuivTLmb0XxmiN0fEPfTNydJNAUG8BoqWAeXu
P7wRyr9WpnRPYhumJItd7AXqCFNx3SKr0n1BpbF8JNcmprnejnOvUHvlqs3LB/v51RpsMQVLehPo
Cbyk9nqLCX+/rmDfwQlyHAqMgl+yiTVeUpffTY5mk0j9wUFx1wrzoVAQx0MvNBOoW43fPvU9IS75
BIa1tSdJQ4CAxgYHfSAl/qRSNLgMo0FLeEQ3VzIM81litr4c8ZY90N3WPgecwoiR2Qn928TC+aLc
rY47vBOZonlHRHkK8AhaQxn8ZuajBKSp6uZtCOSHXukV/y/UgfjG7lHfxPevzqh5Bdd1vgMMM/S/
4iSaykpDx6/oAf1gGpBJB38mXtzsumpWw84WEG6EHY6gPwy/aNjTx5jEFwqRgFZ9xRuYPbgtPkFx
HOZM6+zj1J81sjlRx1w6ofc0D4j6xnPOiUkV+R2KPq3vmhCVj1znCQWwymVbghmhVs/M+L2L+R72
zp+RXU4oF+dAi5EYDecmR6PRj7iMxXMU7tgUQBQsp08mPRxbPNdLHsvf6Hrm/lVuNDagqsp9/B93
7P5wvLuXU7R0uv38jcQBG0XC15rDRSegngLB8mo7FPcAbzgB/uoel+joicmXDoRPeaBcYyqNxmjl
U8rFsgYr+mT6QTIVzlwVUIL2Z2S4336kbncYXKVBUkRvMCFN2A0A+/86k8SXDLb/1olR7PyikezM
kgyV6tNj4CrNanAYZrQBFD2vR+EaAwAQVJPKAhq1SuQX4Dn3kGonIcd/y4omHbAuVJjpgLKwFUnu
orpMq18NZavCnf4am6y6lYxl9e66dcni0cgK7n/V6hJSAweibc1kC/fRt+w5jcdMjtrXLmV/Jn2e
6QIRhdtAm/hNYB1mMb3gRERWE7kMDL19Xo+z2XtgFddxwnPf4F3IkkVS/lHOnX/5illLyDfVY8eA
/nw3MycoXqJO3Hw2m72krEaNvgM3XBkujOc0OJ7RU75gbrun9eu60yUFHgEhQT+FmZ7vUSyNtgKF
Seu2mHXLHvNqG6qPipXstDAfOVGYsGugTiczQKd0S6furIpc5RDkFn8aQXgsGuO0YN+KrRXq5OYt
rmnO5v7p6cLpe2poc8M4/uqFu2QZb11mGJmgXkTxHZ6xsMm81xJ5rBcFOVNu2lqAKZM05Gb5H9GX
qKJ8MWxDwjT28EeMrgN1BipiTZpMcDIHdjolY3bE+Y0+gpDLkBhi0q5br6tsSuoplZ8JLaCEqaMD
ewy2unpniMCfllWXQNCgJ0+Os++EJwIcqGVR5uHbBlclV5G+BmRG3UyqK5qJlTOickEUl8VzMDnC
68CEnosGMBQSwsqJqrKYvzZQ7P0FXhRujxfZDyO/ABBm2WldW3ZU4BKqIugHIrJbLNXM0hIsdZjM
ciVKC6zxSJY5zuvHBJlj3QNxx0fDu/dSh/WcbAGDupZoxtWB4jks+hkrC8cKf1kqY4cdTW6GE4+L
to8ZUwV6DhQjbVMxSU5Ng7EjRW0j9iIaPXPNBkh3KIxmEme8E+CL+AUiC+OvGf/Z2LWz8xU/BvDA
HPRVvOi+goy7oa3uloOS3LYMhLcrF803ytmlTLpn0HDgiVZxhxgbraLWD0gpDxjC8XrDQTaUNKE9
spC9qe2LT/Plh8sg+Rq8g2Cmnzw8Wk6x87Bvq0MXspgrz7lM0AMilsKBWE7biy4QBQ60W+DF5GmI
8Yoepa3iFCsYwxj8NN0ZGdf48ZicZ0jM2YwKAWvzQn3MVo0JM65flt2J2EcK7w8+is5BpKRui+qS
v0pOLtN/yhbEB3DI7jMWy1eIh78wEwWrIAB5hRFeMyxqA8m+U2IaaiV0pcHSmTBLnM3Pcx+yW1JQ
WPWl7z2xOcpkTrKhO7HkW4/hdTWViRp2nhZOgvfD1a3eY7E+zwhTGvgr2fj7NigW3wf2jwNP6UKH
d+e75adx5vTBDmfcM54tDyoAKRPDU6TBhrIoqD7FDgCPsQFOQscxg5whhn2EvI93X+RMZxK75fCc
BQfH0p8Nvik0drIame0IOQ7BhSZHhuU2u75q4d3jWqedALegdljjvmuy0KAd0fz2+X/E87rX5plG
wZYCKE6xGv6S9zseTwkpFjC8o8YfwLmg29qkq/XhXmYGSkJxqBeI+MdOfHYl6pPoyVfBKIFmzSBT
r++ctys8tklT8yp/7+PqUK1NasAh7Z5qAof8WCnKgCZ1tI7h+uU3worRWP2BuoTtYzHOGbipTmPV
gA/Pv8e3oRYrqKBDqxwVoP9KniU4UBjpyrPyIhIrkHHz09SqHpMYuMmFSnEtU9kpnEoR8qEqv4f2
E/1zT3hdclc62IIzToRb3VtQynpy06VxThSDaOIXuwnRDeczfNUFZWkgNuxbiNBxtfGzJpJ2KSv2
vxB3s/ZrF+riutOo+O/nCUm7U8N4qDckhDjMDdbdkbg33kKCqBQB3kD/85i2AbPtNBPu2eLKK9Y8
JTcJNBfsK5RozzsCxnMrkmPi7pf4i8XvmFyzbk0qx7hBMO2CSR6ebFMpOyY6EW2Jo4k3yZIXgwvd
k/brG27/cSJheXTHQlLR80eKaOIPYAsR9M26d3CfKGWtywLXDBcYP+WYOTLoJfGJX/2kcritETJe
lC4hhEELZ0UsVi2NunMBjP/SWuRRnU8On7X+71Saf30LSBLev4TkJM0wJ6rHoEIQ0UEk6XAP2ViC
q+fTt/apQBlNlXIZ89a51ixc+jjG6jRlcdvSn8sMvY4Qjs9yh1QgtP2uMPsNe+KfxboLqCzOA418
48liLRKpqCVwnf3KeRcq4LGyDs8Ovgt18ZLl40a25yrsHK7+9rAKtTiC/PApZm1+SYIO05S5z4lm
9QUUzYoywp7PdrYkb1BCBv79vT+Lt4xjqBzk32TYmYd3atf9chUtQauATAf/nAW/HWS7BAsfRFiT
qBTTxjMgDnyAx0UsfkFcGY8bOeunyJslux5d6mM7Q9RQI1N3JR2iN2xReaA+hJjYLhchEbyzcnIN
QABsSvpbVHTYoKkFT70G9rrcX2Wd1g7QRhVBcSnwcReS3Qz9k+n4LnlxRFpLLZjLnlQnTzAgdsMx
XdxDu/k0xfZCCK3xWkJy2fsNvHNbUGHVu8rtHj/0iyYI6Avsw7OJ1b2MA7GeKVS4qdPb2jRF838H
B8ySsu/JNMqS3iDplbxZZnDQR77ohjOpqWv/oR3k92tTORR5/nWPecOKWiZ+b8ez7bOohQ/KDbTf
Pky4ZKIkvRyOVhP7y3L97pE5vZuJR5KWdvRZr9gg/p/og5Ev2iPTr5EaXU0Gcb52E3/VhWNXnArQ
6TpO7O/WeUmGq6iKu9iBFHb/zLLSr2QNiTl1xL9yvrplgzY6dEOXn0Amy1fVXycM2wqQIdGqD8ri
5RmyKiEjPdyzGCarPO23IloVDebqVJqy1F4htJLfKh1jZJPa5AWmaYkNXmiywe+RYrHvxe5cFuvN
5vw2AQLejnDTFhaJsd9Jd9Ajaml3qlKt25luww2O44gbrYHuBCxJiJExzFzUgG/hyAtpKZsLv+hW
V4Ze+nEDKOTQ1my5sDimHEr17SztKm+YhdKbzU+0zbLKZXadpQymTs7x84vAVZQl1WByar1DD21Y
l6lS1VC6l1jjVpzE2WR7V8zvy03XPI2BMIC474DgULPRcz1h43ITGj37YbAi3inaUa3NahgQ4Om2
E/O9lZyOqv/Bb/1znKI6g/+E7RdwAAZmvsC2e5yx94a1zGbz88Z3lHhbi93KGmZSSFV9FHjpOup7
q//FRgx0wvWotdqvOLVEBRtT153aoRa+MopcxpP1KCCVQaKpT3esjFH/v8OOtrxcLRP7R+d+NWwa
lzBc9m+XC9/1JEO8zm4cnK8BU/ymoNw77LkoBhcujxXp8U2LdcIJTbdDUWS49jEx/2URpzlGAfc1
jueP20ANLZsUf1NguvxiimvrwgFHMTb1Y0FphVQVW/nEScMELKFaHY4nieo629qpU4PNplTSp4Z+
YuLQUGBFHdAgu3vKc5rYQdGHdBjIxXdHDKS/QQcS1NddP5mOz6Bi/nvpZf6VN8mgvbAb0TNvBQVv
PHl1FnuNjaqbcP8ZoWJmK85D29PsjrUJcJ0qPfvjwh2Pw+0f/i5k4vO5din7JmbJxYeWietKOh18
msCkLPt0vbFLN7ymqfsOD5gLemvvU6TiXxg1Yl2qQl3UAdZ2lqpp4hdDQAg9l6IuFF4Ou/Ql6yaC
3JunoezEv5o7B4gwgRHoqQbKWxQInOTkR0jfDMbV2AarBIelp3aY4NB8itL54OIB/mGHjxzaVMI5
mPdju8bAfKylFFR1LPNDwrOGoP/HGFRG/JmmxX+EKXjO1ajHics8hk/jgGp2KZIV9b/Evje5F53Z
S0s3VBq9Fjf+tEMCmq49S1vy9O4EMXehTUhWkkFYkL7rmdSL3mnZ66NMQynYt5gSpD3MbDf36RyH
fmjrxbAm5SbYl5D86PXuqs31WBQpVK5uXOWG+3IMuNP5yLvuuy4rw/HEM6r/NK1H6jDzq1N00IMf
0u04w4U2kDDp9BHjkog4w65YZpQGMthB7z9iMyVsHPOM1apjY2ZSkpgAx5jyGuv3oQ3wzVG/LiSI
qyYfazQMAEYI8UYuw9NurnXdlS97xZaZzD2STFhlN2aoNfUdogQkY0r9+2AbpYiBozRNHJKFBEVl
ssC+vRIM3eqQH/IE6KbNis3HmerxgUpQgKXMQnwnclG0UxNmbPrx/Dcd/pxA89YVSuGFGmIkAEOs
uGc4/u8NQoKTKiP94/3asoaXMODYq6gTNfCz+EznDkKEy83xxSDgP/rwaJGcUPBNCCpy6nmjhYcv
rjB62Z3Q9EQA19qFB4RBiJUp9S41uFG5wRfHW+9NzvBzUATTSqTMOjCOuOff1sp/xryM2OSxzSeZ
8dHMg3SaELrxz5aAYz98DprgiuRV2/IQGk13Wb4JopghNSIUaAguoa1ZRfFuuc1fg8cHnVLvMh8H
gMqgWm7iq9j6/5vr3Cy5rLQ/95aOUNa+MvdNXDzJfWwj8L6atfYEGY6wzA0D34pvdtyJ7FcmlIcr
tChjzJ23NQ8EzTwgQdou7my/JOLxKgFl42kCHk8fftqFXTjgDKB1PCii4GbEGeHSmd0QElQu025Z
/Rhve7F6JoquhAAlimQxalbbVqOx9v9whGN2OcHlqqS9dklOAcD0QexuB0jSmnyC0/AN5mqejHkc
4Y9hfKbSVegi9YHj+2VRw4hf/d0TiHSg6V+nRFUPTo5atRlxsXag1Qw2GWm3UToNY9GDBWF1CVaa
O+CCYBkNtqzMRCREJmm1SdIwmJe53wJ/5DCrslpjKNWeMIqHz74eTiRndN6DrqMhapEQtYgVTPiP
LMkChgRywMhzLatnqiKlBGUZ8+N9u8rrSJbrEtFslefHdsFPxL/z8IxYkMbX9++K+gMXuPX4InjY
9IB+CAguqawdbKJXscYb1LWgUTLmWygJvYJFR264BMhdKcvG+b746WeOjcrKYRefzD5vmDGwP3Ju
uFwhPEPL2v+VW400Bof7zuhLnDjNbnT37jcQXiGwttfvpWupFLcs9Jm3qqAdokcL/uCPsyjCWf4R
yCniYpJJv7tFBYLy5/QwTwtO1mGzCN96WeIVkmYZpdIjXNpgyDIKKGeBucKvUMUxT35efxCDUsuK
jK8uewsaGR54QqySxSLn1AWQVCw5gf2O9K477G7KW1kX/QrsFbrvV+NueHVoEYVJZaj6VSpVvvhP
4SoTVFPArb3QLnBPBsPaz7AkLZwbx4/rwMQGWkP6YDbuQ36CLVRpF5PwNOZ4XjwITERaBxmkNFQf
/x1kKAteh6aO7woXUboCHtw6K+9SF/C0RDOmmrTFsoR+Ux/pTr7OgZZQ2hajSqtLyx6Z9xMc1MNM
Bf1UL+SlXOG+Xoo9Kth7UDzxMTQp8SmkTJ0iKh786K5h9C7fgZozfVoF7//0lfIUzfCobfjMstre
7rwbUulX6SBk9oe7SfzwA07C7ftckdzaLeBUqvIYsKDPCx31/T6GZ0jjC69i49PBzO8jw++Fi1uC
dTf5Zsj/TfvtnB/5MqYgYClNntzWT1H69ft/KRfjFmSH1iJF5QI+myz6LSPj0TdawlrxWqD33/J4
AB0LFhaxdvffRvC856SI3j9XlQhF7NJX+G3tcTKOyfR0WlTZiI44ikcxtiCzOQuyoByMjwDhVMBi
s3mCy8ehiLMm3BNhnGc0MYJm125K/ucMYk2SkQFlzlpgtZeDtFRl3hu7w63J1xYVHXBSh6Rj2HWE
+CWbwiISnlSS1jFnC/aNkpJ6bFl3RX4dYPuxOm0Pp8tfIX7+lAZGLmZWypFlmHrQ0GRIJhz8OIXx
y7xyXQzllAqOJy4XBE376eQOZ25M9d1GodYshTAePxeWIbNCRZ5qxPv0UGGKY1HKndqvNKBXk9wq
X6Cn3ocZI2+aqBi4eud+WcLEJ/vy+esCZp241qCMUabIicnOaHHmovy6UWGCmYZqq1ufSLrg2IhU
m2DWo/Fy52SWe6O3fxWgD9EJpY6XLVrHW6gQeoqjQPfyCgp+J3sEviYPzL4atx0J/JafRdmW0Mdh
PE9J7UYHxFNr/nDYCqYM5MH/+mXuPj2hxCGBl3HKrQS1PvdTP1zxrummyB4rNI60sN5LIYWX6WC/
Z4+KF4Y0fdJdSD7yIH0BzpXStgbY9biSpOyDXkPGKHfRxP8sC6G3w/RUHaOE8j+46quuc+BTk86n
GsQtdGNVr+ct3CVnm+1Uds3OsQFpytBQPlkRW0gkIKkYO3XZU8AtORdJwJ/bFFFm3WDHXPUWlxS4
cREPRb0E8KFnE5Pfn8M6oErpsMbak7aokzWp/x2nrUh3CXi9cTzLX6fKyY73IBz3dPvyCxQNRtRe
hPUVt6nuQVDZvYhZI942iqGXrK39bETzpMyDFoGVdcWs4B6Qo855X89M1fsn85ZwvACH0pDUlMQu
FI5aLnwlTLms272MVzwTLIC6QjJKPpBqEcVvF7Xj1Za5/1Y2OH0GtYBOHDAq1wnGpU84QrgOrg+o
8gJvIPly5Hsr6JV2tNA4v/lN9f0E1tIQX58TyNm3ouwoCbBoBL4PyJa2VCCa66MUV8vX3fxRshaH
ocEtUrwdc8dtD+IVfLicaGfwUxFvHKnBZsE/1KiFHkz6yymXiIBwYlMr65VAYlRv9vJgVJmiDyph
gmjqUtU5ID251LRpukKr3lCUQvFZ4rIbsYJLC9OMcMc+TH7lfHGa18WtQrxM2iYhfqNt6J5/JHt6
whxjOTF32xmLWqHQcvn0Q63B0r7BojXNtBQqrQ29y0rgfhymCEMkLf0iTsnB69VMcZRQ5TLo73JY
xr806fS+ZsUs43xKjW8zhBFQU99+Ld2Kb8ZaZjNOINRK6TFMsU9ZHpOBsmVtLiYRufT9mslQcxxv
iVKrzDVI9CyuUAVFaHkXZIgLqYByifnbf4Ivg8CEjklh4SEkIOhgMvgOoswMf8dqHfU2TzTdlClj
i8D9ELrMTGGZK33f347gx3NY5uY5F0uX1Tj9fWQbAK0mCU0IxB4VeTsNrm7vV8QpT7lIpeyprs1P
S+clrC6OlPfCl59tIJP69WlsjY4mXDi6CU3a31pxU97FVatS3S+7ND/ibi0X3woRThkOZ5NFiHTK
1Y1SZndN4i5e9CXxJ797dn6GTC0mIujddRO83a4fni42VTstichBo95vSE9hA9Cd9UoitDzR+cW4
8Iq/frZAN9BvcJN+DeDKvvanhVVmbE0P7FDVorTqiFA/yPvjS+99/iAQiZ67scHbxDi4PQI/+hsn
cXF71j4lCXE8xyDKItfFwMV9VsML8XeHhBi3hphV+eCJNnT3QqejSKScNKeKYS3xhWYock6T9Txs
eQEzTt8sKi5IU6VDY5Lq8jwbClESYC5AqjyF60I6J8rlZclsco/trXf/uRwa8PZ+2YQL66n+Nyb/
kmrm8qE2V8+4qyql+lXwX0OqG7Tn7JUCiBIfoe3iDrBOySDuH7PJJf988m4r3RfUH2k1l6NuPVfK
No0AKling+Xjzkm2oNTSIM/T3DZNeU4lczJkBCZy+nGHsaRzRxxbtm8IYd69HnkOwUN53jmx9awr
lGx8PiCOIXQBp/f0IHrkWFAvfU9ZxpQN1B1DnsDDvMFAUtcGuwYMQqBmFQOQiN2TytHAUo0mzH21
hYG4F+Txgc6Jp8xA/iQHyjy+CldYcJBFaaXEHHhNT6Yp2Gx79O92/5Ym02DTP/oHhdWNUQnxNZJm
WmDFBM1Os2cJ4xIG2y8ZeWa8kCC88FypqegCgqYqX24nupQkuq96lN+6ty32dnHbHBlzK1M3iOis
GZj4gYN3u1MGMPL6dm0aNltA5EWIEIk8kfOSQxiYPBs3OYK1UjxfdbBLUkD+txpKMJ1AM4dkRVPo
R0cFeoyIUFniyuPhbsWi41TfT53HcoyV+Ku0cCX3izq2aCWXCD3wPszO39NsAzqEazd5Lmy3ivbp
gjFHQorxC92OzBjjUPSSTiWwj3Ic/6gQs/cL5NLZGmK8DE+qv2ue8ipRakSXpEGZKIC7KANkEZLG
OxYxcqF8SKLqc1SZHO7RHe+GUoPADWK3iRa2kBElIKdoA2LViqEgc+w0thURFueLKzgUNsuZHPZa
9Yrzsiooe4SgzRACifCG2tAOUf3ygdjJS9lVdS7+HxzwKCRTyCw5s7ioH9moJXGNunqtqiOIyLK/
qou1QRvKtNJgWMHC+PFwsoIJMpSapwxIi+3Xj3N2r+QRLmWZGI69LaFOy8adBdM1kacwBWSWi1J2
nLtFJ0DKUGMTHxHyl3seLK1Cvyht7WJ2SfwJnOJtJWTOYCOsJj5+Vb3T8mb1YYdSmwqI7LLcsOHF
KMTo/Rz9jH64yyVtLJVxAiHChYsByol3/Ud4vND0nlYXGWwKgfzaOJGzn9vRO8DYQY2KGPjFWQwM
lhiJy0jWzf2pK3KU1LNU/6rC+ZLq4LjzLR/WY8eW1C8jmxLs8gg5DxLvyir+RqOvnFf6CKdUm4NV
9Qqgfs6+x9OaBdoBOOBy3ubxFt1Wlreu+07Hebn6eNAZ0C/XFqVbFbSmnJoACW43zJH8FWV/VO8Q
5gh0KL0OSjZmEnNNvRBwv/XrYqEN+Nqo7GO8GTfcC7M6YWCSfI3DuEv9Su27dJM+jWeOHAW6KJKQ
g807AbQQy+CYIuNkRGHU+BzXq5Kj1pOdEx0xGTRC8hDi2V5p6fWfnIRPYWdCDYnQ1BJdeHul0tc8
Eh/9g/6fIDWJEmEKUXsdIzgSUjrt6w2gpDtHrzaNrPZGjL/PAzBnPDPtY5z/oNKUjlZKvt1Kugm9
sCUrbGaHKxO51gupNfUFroGLu7ibJ7rGHeZe8WOGUHh/Z91Q/YT2pwoEAqykQjMTHFF8gikso48j
uA+oY2ZRPAS2l9Rt6TxZSvUeR8jf6MWkLslLYWmMngsx/5qqZuhTZ1wWZGNWPlkp5F9xWOzVmUae
Gyf+vhnTWjW3fNr1EfbnQ+kUH/2ZxQPs5W8qo3swwg8EqyFFK1AlJUS63z+P3hSV136O7V1L3Iiy
qbQTOKLAVazM+3LnrDj9HrxO4egVLu8R0Kfibx4mcy4wojJCTxMZQ+4H7BlDuPAphpdBG2A0oJRj
tXX0M+BfOwcgM2bFH9XcBsj4BpLSq1YFkd9mtMzu/LBQXNqMY6L+0HeOIRQ0R3E/se5VLEjcHpVj
SnUPyx835EJ7052kQgxaEQiD5Ukcy2YC4KSwTuiTSuV72DpmdFyfxvRX3OO2qqovDKMf8SxGi8Vw
Qgh4EG4aia2t5gKsp/nxSUOy/AN3rNaiJoZZ6HlrndpheQnne1RzERTB7PZBCjlgBUMqhdn06XWP
u+2iYUwGysf/evl11hAmQV0kY5vR2jeFaLIrwoAihQoljHsZaMlt6/gMCa9Q9kMlvVgZJ/xAosvd
kLzbr3XRQRUjJbgLHGTPSiBorAc1Y0Qbv5Rdz3bu9HKtv/fr3qHkAcvw0doOU6qV6PRSxCLrk868
QgaFVhtDylCjWYdUOKMaaiW7tDg4sq21BifNYO3auuumh110vFv8q2ssdgZWsFG6FSV7oOGBiPYw
rlz43zsW4ohtj1c6fRT/aHobgVaSthF4N+oyr7Uv+E3w1zy5APXKV6bvq0Ru2YZ3CMQEX3euMkyv
4/hsFtbpeNZUgBrtI11g8Y4ly2dsw3jjsD28Ygid2Llm6USIdjUy1puGC4ZRIoO5So7ZZ8SZMsCK
t482DsbyMpSSLHUrPfLETwBmIL0dzi4KPvVzAt2/l62GVtbLC4XE5rrwGPkQJS8fvgbKNrqNte2K
a/kTF5DzvMBV5/u4iuu5rTZ84VekAEdAoC05SS2QfoEevvqUK6zrrL7efoe3CuAj+6VG9D+SxYcs
Imb236bRzg/fnbDv/bRtM2ZK/vUSA4sYGxNsJFat5lJNHFJw4lA61ylZjqe6t28y3DsN5CEiaQFN
GUU1szJb1JAVBC0M3J1wie/GKK+2TpoFmqqOYOaRP2iWQNN7FeRQWMuJ1k5fj1C4ZW4RFx1tc+Mr
xFYXC+BhG1Jsmr31huemSq81Xcbe2c7m0vuB3U76//38Ie2Tki8Ycly8qYrlmph4CNifqg54Jh56
runfEIIjgIydLqeQChkDI8oRPcGdAy0iLTtVNqWC7GqDiUo8Ao8pa+3/2qY5LCzJ8+B30NtCQGLY
kyeiT9ujhnGNWJKrb0LfrHfO/l+ODq3BVKMrhfz3++qzygeRrL/4+FbReF7OZhC8sLFZMr9jBZdT
qntWglIt7sjzekbu1y6uKBZVKabebLzPhiTok3q/t1nJtCKF6sEyXT3kY/YMCY17Fd+dPntnDDi1
y5wmUUmS1VPGs1BY6HvKnX9X8RNXk/1Lz9WuDUyqGDqUPLhGHmQUReovNXmqa1xBNqGwDy9ViwHO
Z64YmiTdP1wY5o5iRrGOMWdfA3OLJ+N2klrIxfeYUUuc+nuygWk3ohSUfwmDISOkDUAkeEePpc1A
Lfo7xbmjBHCQsW3XS0JnMXkDnRDpyqXbYCRRm9gICn4K1XY7N9vIUlD57YKRVX7H9aNbaO020oVh
fLVzATZJ3TWCKbscblfeiGqYYL85/CNPVPIfX8gXkFGaYhkzLLXCPHvdZKXGXoW7TthLBl2kb12o
guwZRTRpZPntSDqt+Li5x1w2tJ4Nag/wF2yOUeI6gnWXyfhBRsE5ul53e1DjnwERxidAdpJxGJt1
ODG/kuNs9VVFspNc7EMiGxsZYuJH3G1phbfwppK1Q7GDIl1cheIoYtRxJ5IGR0W4OPTKZjPfeY6N
Ku7tCMZNPn8cBZBng8UpF2PgnNHez3MquCkxP9S2d857tB5UCi/HHvAgYzbk7GMdoWcrs4zgoPyS
aAX4PRFW9hpfqaCs8iV8+XkPZYDkHlg9kUZZb9uQDYphtktNa/hTqq5+yZDdIDVTSCeli/qEtEq8
wkD33H4O6dFjDXrL7+mps35LptZhIkMigjlRwqJR4ikFMmK/sPk6vN9aQRJtRkJdJhz/Bc87bLFs
qts3x8YT6Fnwghrrv9jBnK6qeGG7Nw6wI/X57xCeTXU83VWx+6m7qba+CD0Vset/nbnFkJa4qQw/
YVBX1Ox/TmR67X1yCLjA6Mc5u9UZsu7f/GheTnTkbosSLEg5SPfi/btcDCKEsogyvu5AUxpxAlKn
WnAlNcX8oT/qC6OeNKfK4ehrHmlgbHreCHmiPDvs2zSpiT0sXXG3hazDb6bpvkuNiQRBvWU4gI9w
pXfGpK7ZquqCRvgYg2/w4NLgK+jtprr9E/HB8QSGlaNLX3K3e6frpSCxciqijQLWttJS1Y3sablT
k9LVD1+TeKduNVzlA/K2c35Cln4NoiWjFW9E8QusZsauMco4q1WodMDQI+03pUmU3p1gul8YtV6y
ZZfx/LjsP1RcC2CyJ2NdoKaAWb0/6lVkBpkA+LLCU98ZjXebvEU1IDYmPfPlNbE2AHiWoYHhLwjU
fHBnh9qUfZb3IjIPkwKr4QTS+njXHy0rmplCcjeH8DkqDYdJQ0RLKxlBCo8KX4aTfgSgs3K2YbgT
49EbL2jsLCGthy/feZIJ00mR9NOExDXYX+Fzv4qFGoFidP1dAjYkm72rm/v0cxhjc4S6EU75WeAg
+RsLA/viAbSIPK626X09nC2HcPQHB49CDefH+fAzClG2oKTUT8J5JVLRRoPMuZLJk/Y6nngyg9nd
87q+Np1NyvBGT64ECAgL9x78vjWNuWQpXcGCSwYzttZBdcfaVa4s1iL67vtVCk/1CyUYkSSxN9oQ
RQG5YGHGHl+qTVvajojH4X6SNvcglIJA7kIDbLShl1JbcsQmmt79i6XRGyMPW7q9bJ+DPMlw86jh
GJkYU+3PAcbMW8KvPVe0nIVbVHaoYn76cLRgsWLRizhFyb6KxuOKGavOAPzk/4HILtvdSgSit2I0
HM0UrH8OSPFbGdznFC7y0tfaC3kM+7D0M/GkeLkMAmuPwkzYHOp504dndxdSxuvMbO9FR/Fkrk35
h0v3Q/yWO/v/cbvsTRovn1gud5+oY9mB7uoYHpL/Pjh8sxUsEJzZWjgBlWwCsxN3QKyoROyp6QCM
y/arMxv+iizYH96ReEzf9TNOqb8kM+I2WPjcBkNNSrH8G2yjLbDWBd5hPrp15Ju3OJVQMZ8AJktl
NTJT1gbL6sx8F+x3i0CT3gsJjoZlAajyPySXSnmQ6iRdiZzC8RzJPdvM4drBslAZiwv+W8xmo6us
rpFNs83hixH1uFoEDwZuJOnLpIjG8HXArYBkizi00gI3ySacOgcoxFxoiRx/Z5S/fWENTLc8MSjG
cTNusrtty7mHinPgRNrr2jFYuCVUJzcvG/V6qizN5nJZNSAB8n1nv93BLP/D3CzlMVfYoaJAtCrq
tQyoLwcLvOHVN3l4OoxUELgmizLTcnrzRxvxg7OBS31Z2VAga5cpgf2ndeQSlfKzIXQLptHg2kK3
d+J+5OVMayWEPOCOpIjlPaugBKqJtYtrGH4sg0iyQ3Hk68pyc0ym7IGfo4XnqyY8aJR/oH/8Fvv9
gdqP6eT2o6TQgclrEkpvIG5pKrMlx+RUiq8PayXiNmGIvy9L9AolWbo9JyW3YxoVa6dOQruWWEnk
Lpe52fPABTFeh5vA8rDnJmO5ioAM2hD+usetVt0QvbW7kd0toNUTpUy1Wy3kMAREfofX/y6Nka/p
Gdd2VZUhhBn+Cg/WWnp6GcOQTw2ehpuJuMXOg8DDcQMAvQhprA4Suw/lCcC9eBPNyS7PXw74Z34C
slhUtQi7GvSSgLB2aaFrTduvVYBvSG1MbOp+jukWpL4Usej3NeW/4VLRGtbcGskRwurNm+pITYWl
KDSuPqO0DuGY9Xtjtc7w8Yyc0a6poQjItosPFubuQxcOH5mueFjFn6zjqjwouElRaFWttTQ3QQNs
RBVctWzY+fjbVr0hsFa5rYZutp5ix6SbH619dwZM+R943qGs6q8SWOjpH0u2uCoXJKyITcMlGnFV
6If7s+fWtDRbzliow4A93vr4D63c+u3ydvqtouVtKCY/fv7QP0JUy27qmgoqj/30GdOOtFfGLwot
UcBwhk8AbMqEGv09fGbzyj0PwN7iZXYVJ1R64XXM7zoc2qd+GJibAomxxPOEwn2BwkPsqwGO/wZP
WWQz115FoLbI7Ao1MdkX+p17GOD02SUfZFpoa/k6sMbJE9egpMnRVuncwyuEymQ3uEFNVLByrIPw
aX/1dAFVyMl1wmX0VnqTk3uaedXqxenkWJUFcoOCFHpNSm6Zkkl9n9vzznFHAGYNh7p2r3dwsfTG
7hh048gVjtTxFPzwQNLyTTZPzJVz2JunuRg2erUnct4mx6WE75OUhT//MkLsZ8TCQKI0sJYZoN0f
0IXx81WsTWCwjKyKBAdVqwpO/LNbe/VwvAzvO7eXAeJT3A3NqCuLeGYwxAd5wn4MStr1UXOQWRm4
+xaHpDJQIoTfI2jYeiKO4J6OX7Kvr5umXwZ0t871E3gZr7swaUcxVPqJk7AoRdB7pJFpRix7YrYF
7IZ8Q2GZ0n/4HFjILzhDJ2gRBiAxzcgD1Y1J78tXHWlYXSlJKbPVbIWCltuEkv7fejk4V17Aa4we
Bg4eWBVEI/5WCu2q6bEn4eKzl2AYxdYT5CWf+rd6afMB8SpKVXwhe3BPSoh9wWHRgIDvPslnqGC0
N+vLBiX7MF7hHPO0Tc14AgLPjZ2YoqISSIJTSSNDnbyA8X19bbc8afJ86fEFLpdIBqZaYtXq8Noi
zp41uX7Q30Rxt4kTi0avbi8yDjG+3QWG9tqhfIV7e4KVEeQ8QzVHBnApf7SPcQSg+qtpqK+3btSS
nGQ7SViktMfRazSpGJImGGAgtTYsh3PodCFfZTiDmDJXBJbYorA4JHpaIC+9GqBUcn1OEaURA3Io
gmIQOnbvkCq9DAgubrCInu44hxzYI5eGwCJngeKg1UFd8IxJeTKUpzEgg+jh0iQLxi77EhcMui6V
KgzmtxXF05gh7/QWTkstQJ0mbuLh/0Ea0fgl4vEDOVza6kc+64a6/LM0QTiFZGAEK5l4u2E4tDEg
iVZzEP+4U02J0HBbLJ+My07wM1T72OpoO0XwRmZEgkBl6AP5hJa9I1k6fnBW/gSm9PoK/EratBa2
5lUbTctffLaliphfB3vQi35q7bplDsuvCpXufLQUH9fAQlKaoR+YRrV9IEdGoXunY4+Sc19jmv/c
J6HgbwE0Fpe+a7nTCeuDvev3sqzqnCU0hxvVbzRNsu435C7bg6HmgKW5I8/oM+R5Ro8MM+mWaUh+
7+mUhby3RiCUn6CQxLwyUEqHqkbwSN0LY4hr27JuA3uiFui7Hx8aPkt18NQ+ndIdvQQuN3NtRGlG
NnAZK+tbIZal5JbulKTyItA9VFdI+eIIE3qTAXO07QJNO5WGwYM5L/ZNW+if5UnAChjTjQUd8wYb
Nomlie9yVYBhdkFLRlPgE6ZDZPbdfqDkeUS8s4pmDAcFBMRd5X/e7e3bSCM7NaDg7JCH/sZrvcAS
WIG+vwunmqFjoMDAfeK1t0Sa+pGi5OfEqVOMxdkAdVPaPmx9ps9P0H3JDU6yygj+yLweoN2Qyod5
XL/XOCeLsFy1ZGfims1Rcmo6rOFrY3X3XjSvPtTtixAjfMTHBTZm0eh+nrMWWgJ0QGd5MV8Gv9up
/MjUrNhQRy0MMtPHFVCOT8VgVW2bCSjA0UJx7VipGKRya8cAefwyOw7vxhFtrs7iwVSdmLSg3vJ/
4R2gxZirw/APG+AD97b/+CeYbwrnQm/MKKm2ed8v73zlN2S6fv5h7WHlpqmUd+rC9r0mHYQMAJq/
UsyLSW7mKUcvDDTyhpCXJN1BqrB8GBafswG5O62fLnsFGevMCLJhOqy5fImKOTK40p005B8CqUnO
8no3U5OA0hoZI2Edq2uZRaVuFPQdlKZQHtKEGUqDf7brkgM2NznDt/Mx8vtn6+etobgj+UFLskpX
YM1rk8tSigMWfJ/GI/F/w5oVg7l6C5Sk/74vrrmukCbkBgCPjbNvNoe74Qac3iVk6N8jAcbq8S7v
LyPvblYrONoBX5YSNZGs6j+7g68+MJ/z7SU8KR69T9kDl4aFEsfqotx68p9I3XNybx7H7OIcZvwv
5eYci1b/7yALIXcLzBng6OvGOXLFWQasnpI01BMmIVVdMk8F+5DTxGUbOvLXbn4twvDnLB+6qE6z
juKhizoj/m/5FDJX2jIEM3PjNGH0zY9KTxv62BteNc7yQZnMGD2Igo59uuRhFaB8XIu6BonghG4A
nGxXDPT/Ij8Gs7lsnOuZ4tO25JSIfrqTFW430y7WaJZ7GvbUxhFFfA4Teb7fZaConY5sxvMgBHWg
1l4EG2LA32LZyEwPjaz1LSiQPD3uiS3oRg2DoGqMwkWHzucmGdqFaQi+QrQN/YSnd8ACXAmUX0zI
IjAc7EUCPM2gMInHEgRHF4EoJRxYQ0cttyPxkWLnyyktdzSWKt9lOg8z0jz+EIl7oREQXXc/nEXk
HgHPLSuYDm0EP7hpmDFYUVjdo9YMMa+XyhLkqZP3ApEpr3gBEkGINAUYYrY0ptBSq1qbIvCMGF4L
ewVnXCE57THWNPtkkYyAdZlwRaRsut/ZksumPtYQ2s5R4hFAYBqfssf7gJQgTU+n891c2NNHRPvS
3hIsI0QPUqQzCzPkNQWKxXj6z9W3PnYdA6aG0vENmrm671tM79OqV+mLR8gKlLZJFhaBEIlKG1hJ
Ak+IUYxD2zT12XUEHRMgXf76JXbyVAoRxBvPsb2VgF7Pj2Y4VatiUnH0u5X+Z8/KD1M7ycHii6PQ
yIKPcREzZG9Ks7RIOeVQ/1t10FdYqy7gMW488fPpoAtHQC8qr+a7vVjq4lpvavZgz1OYNVo/Z484
byVAZaMn6oQDooelppf1hp7dHQJMahf2haYNloElAn01BUVcBZaHcpEzFYoMVa9LO4KIAHzy/JkB
UT3oOqK6BI5pgkXkiralNpcyjeYLsxbLv1qS5pUt3RuupNq7tOcH9JliRWwIH3Kc3sq+1VGOeguK
7x2kvgtMtff79Dr4rEVZVk09lON/d8XcaV3EyNEqKkxdAMwO6mJERK4BoX0hvz/1+YhItf4dwjix
QpVQzN7Nxn8g4QbTUTWozwfiJq/8rdCaSPdKjbkVoB0wemCVj6Cl2qm0HFJC5VKIHIAQDrzlCD5p
ZN8U4ykzGVocaAERSbeJz+TcrHJfMZiOJg5QY+cOCy8MOMJIpeoSfy8PRyc/mnMPoOoWWNhWFyCW
QUICahSrGaH4PAaDDWCgPozCUZh448+1SSWBhb6S4AN2mqnZBoYbgABesgPaG3YdoDBL9Vbzw2q9
5NJbAr2Wa2b6Hr5qILbkNe4iyab8qlEIzxXn/HXK4pALAVsbeDuJZbC74i7LEgk3KBRXFmUlXCt7
vhcXI983jseZYkiz++hNtV+7LXFXxzf/ODQIMviEI+VapYAs3Lprl114374fZMPxaq5+ClN7IoYZ
7K/ZFExBiXDr+UcFJ3Fjn7Ph2Czquc9SUOibfv1rA8yVXXE6d8f5DE8a0GCAWEFgNYiPT6vrLxo7
PcN0Wnp+21wwZqC9IfNpQ/Ec2CUDBYlkORZXP5Fdg2PFHjijbfngZ/Dbi9Ax0dwC2q1xFtmae76a
6jlYFm7oUXTrna3MWWrHsin5zqq505zU4rJlO2eZ+M7tVuCDWyp8fzcdKwaCUFSPFvrtrmq6aLLb
6MTMkD0fcJSsnOXO1KTS05HIGvaX6t7bmewKdaVBNKmZLdcM+9+8ot3qo47og/BsA9idBwsMvAFe
1l+QmsKSxgTs0Hl3A2wBTEzh1IgvblVrdT0kD1gOM8Wt3ZFY5R0CK1oXLrDQIdVB/04OOTli81u9
k0TyykLb5jTUAgapLelhdTxfbl+tYuSNeL51d74dvAayj21ywvgjxiK/BXBvMejb8XWRuy//R3/P
PPnRc5xOhq3tprFYm6kT4fifNuyGKZ7yyP5KjZYQJICczLoqpTWXZzcddUcOcJ4FWJfte0x8E+XF
o+K5s3wqQEPU7MRGttApzkOc47h7fdiIqC9hyXsx9l1adrz8pzt4CNV+JuzXCSPimoFpifAdni3g
TymQlVp+uhRZc2vkMtBgzJiPYWal/CicvGjScssfJdm85HdFPdJfMPy6i64i4690PFOQkU4ESPYh
uUmPrYCIs23IccdGberO7oy+Aywa4w00IZXFBXf9alcRZyyyoFKKZYb6VZoMMRizb/ZCODf/fPGp
PZfsSkvoGFbGfSfSNmUJmtNL1FYoSj6o4IUiB/3q4LtMhjZp4eNhKT1xuErEIR4I7Vv0ULQzF8kN
HnAy4hWEY0G5FXObVnrGT57qQ6UkwSYJmpgKkSsbsInrj2JLUQyWrfMsvNIbkwj2l3IE1EDnOKd8
zmXE6vTJ2kWJd7FJoz9ioK7lkF6S7/KOzUzO83AKYi/L2MQ9d3sv8XiXu3bQxP/xTQVAmD2ycxIy
Nc9l99L9EqowG/PZkT9edq73YSQvOb28U6NTNy3OVoHxqwRlCAEzKKTN6GMk//V3lPl6so8apyN6
WSSqbcRuy0L7KxAkYZQ1jPEJKK25yb7pcWstQZrD3cN72KvO5bLZBrvNwlZZcwklzzsfpJpSe19E
FbekVIHik+iQJ62B+Y4fGBzSnOKnkOt4z6T8Gm7bnmzqOIb1egUR6nJoKssEIyUT5hXJ6I782PoK
SKTPJd6F2qcaCW8V/Jpe4ZIlwJXzjVV5n2w5IDeZ3Zp3l4/+tz2qq99TQzHfomJMVKZ8SmdemY1p
2x/LnwHr3RJIuvGOPfZqY984dCYuttnsJ9GfXWVF1zeHyDUDjBGnZ/v5ILl40HgetCVLCuM0YNb7
E8Mv3fZ2cDmgIB6VsXoQvgLJIWe/CpPe7aWJ9T0awA4vBEkXMzOKm0cVNcBSxZiEHLZj13NPi16b
+Pb4zf4wbIUMgRktmgnoDdbeK6v+Nai2aLYZgM61/KqP2zQs7CRkEpGnaZVChEvEOm8+9YARxnzY
S/7Jl+s/dK3OxOIvmL/a+l3WED6KWvTGcu53iCLkLS1RROaCzBaio6I99rkG+vPyS6GsMOYBhSFr
c5OqQfRttOQFU76MNtQSiQ72edpkUQlvEt8HLOJk81ii00i00rbchyjugZnhFQaHVDHH8OFWFtok
bxc+13KE9XvdrjkpXwpLcEbB2bMdl9gBX8XkzNQrWSbCgmgeInYU14RdapD79kl35xRw5Xmz2xUm
y2FMvgf2kyRWEKSGsX9evgNRbuLpxdIWvIP1YrXb4b0EdG/hxFeNkZOUiyHYt6qfOV1yJ05Mg0Gb
Gg0Gay+wt2L2iYlp15bBl+BF9twSWSXjutUPX2SSq0vy1UFzrxIx104ZYXP6n63OVvNSRxsYQwgL
8xSpkKa5uGums8+zmpS0uxdj+UV/69rBWGH76gmi4dCujcz0rWGCPv1gBn58PcfHkBO5D42ErZ+r
mxQ12nnz+cOMFW6iOrDQ0Qlf3NLNV0WuMQnmdy7i3E74r1Od4SNaTX70iIa0L1p5zvgUklD7pNgO
4D9WuE+vAYw1ibaZI+guBOs8GAX3kcfXEAL5wryenr/R8XHBmaOCFZKu2MCqBAL3/1tQJNwH94Ij
i+KfJzAsSD6iwd1uvEfuwew3h9ynkjBllyCirpt9I9JOj7hLa6J0CckZURwd1Nru4Ym6G/ZvLzAl
9gvpceKBmr0MbfMUTFM8hvD2c/Q98WmFDlXR2cDe19CKzbh/ML3VuYNhpFC4wv01YgCCbIYUYjRD
S/Ukmc+ie2gD1+iCVn2j+EUr81/jYrZ3SHV1JlaXcWqruJqHAYihbfU2V4qHBwLuSnBy1eq/NjFr
loVgFTLt5BKgriK3hs5tpBNkhT3lLX2LrTjMqFI/wrSxBvxusQB8CycH0muEPLRe3jolNy3mFOJL
wjCOBry4nD/M8sIwE0AQibYgom6xKo/U8oQeGzXjeEUI4syhU2lmEDMxEKQ2LSl6irVDyAoaE7zd
al3fhwRIVOzFK6ESbqV+v8EVg5xOSE0SuGZFq+ws1fmVMpKxD99PABDt4kO+6RWOL4WMczbTuyOE
Zk7+7CI3ZrC4jiPlFZYFUbzZrV3cTgnduKHXipqQYLy08mMo9ghC2DVlGqSU0BS6Bww2ZpUgWhsL
05w5N+uyg2OPGFLsreYrTnUmU/5uId7sby7NTukI+bV3vTA+tEPlwIQ/JrTkFbK7DHzahhQGYd51
23K6RurGdAATO82/Xr8rA9bmqvXYkJ1JvXXWxw89AGNBxiUNYsVcwcNheKjkwpto+0+aMQLljfdV
ZC3Ij8zXxOWASN5M7tk+9lRhblLnp0bvM59mTZjqpZJhR/jTcj7Bz+OfrhYbaMoeFBbSp8uBHcRF
2hEejThl8OU7/ZeaCUV8yjv63GRXVMqWvAuf5oMkvydin/2L5tviMiT0N2G5tora6XRcDjIZqEVi
+NmeWeCMf0Br1LPKFW9oaQVqijxiwfH8lyIUHTqtGJP3s22QaO2bEEgSh/Eg16UVfWiA3Mat2EHl
jZ22LmU5kiJTgzSsC+XeqTtBGrboUwSTKRZdfVZ256cDNEdQl8txq9SC3s7Y4RkYry9xclxpW0iW
wsKSacYAtGvyF69FgH8a1OMwWCc4drFrUuHLHqbP+N4Yts/4F4xqWcfayiVtj+x0yB4EbMgUaBe7
IN92YL788cc8CVMOAB7krQ5Ct0K/ZvS5prZM7WMpXezrHG/YqMT9ZCanAKJFenQayJHYoMzVHXXC
UnwrG8M2+3wmJL+KBVElv/sXOtlj/JYF7QBSaVJd/p5RmB0f6DvUZh62pIoDwV13w5TDBmqYtoFP
8XRn2kaRRiv+xFJkgF8JGC5+ZejNnlCIrXs1BwHaYjz5nwn5GvqHmLQ3hUdntbzjBi4FKUBMyuao
4YPYKC1ZLraqY+JdACXP0MfmPoxOalf+S6C75BtW/rVHgnIiBXnUJqxUZfC+c/C1K0UPnjMk285U
dMqAguzhY1xvaQwKoC4gTSi2UcHLtSV3jIusqd7T7Ib9SNiLxg6Rqz5/3nRVvFo0mfE/i6gVEbbH
jIlUYa31+45gLFOOwhULLOv/3/SBOCPS/vCZwlM+kz+fXkG8dSyIb5+LdmvPe9NjlrI5RajVInII
nTvTJOwSOqug8hFmmzDjdlUkGc64aGeS0bRF1TYe9s1fgSMHaByHX/GpuW4QB3YbOGpZQ1VX7DrP
utFuVa6asYqB/F14rNvQNem3avmwhs8g0hh+NkOvGO7DcXT7eru9rdC2BDp02ZJxIqPa9Ku6PzNf
dmXDtb/QIoHkXZXo2Mx5wUWE4z2iYDynsn1hHOm97Yyi5JKlUVPTW0TxSeqZWX2bgTbYyz9/I61T
yibPtyi0iw9W+VUMyOWwBndbvYb04G3453SNjfJVJJQc3CSMmWQUFO9NjrDFhkqPzZ9cWQg8dTbZ
pcRIKxteruW29A0DbPZ+ckVSKXOKXbeKVLK1l8T3A8qvYYivdE7VqMC/IioZES1/AWU87GaDmisR
IFcI51hZXQewRFk/mpfTNjtJKpQRcCmbq5VT68Mp6twCDrigDavGf0PR0EutCLKhtoBXwvx0zyYX
rvxKpizDrHyocxturf9A71Pqim24Vx1RkJ7gHm8G80rB7CD4QZ4YJfXOpEI9gCRsorrPNl8pgCUP
bDhbTMN+8m72frMQoN4rMZpUBMhtJvKYFtEAlLx6VQRCAq6+ccLm92NSHDPh8KIvNrsTZxktgwKh
pAii6Uf4PxEGAbWdF/Vwehx0cmxkfz8TLzqjQZ2sCTBCbTzVqJDUyyzi6fQY5cqKxWLsYADsEpXS
XDwzZI0v/n76hwdvdTIyVyZMSCpCCkBH43YKMEVjkPcKWoP1sDUKCeJWUZ+ightVJDh+C56ZUEpe
Kow+ukFASZkxlX+27j/FRjtKY/o6G7sfSNWwM2/XDAcX8FT9JM9GhXy/3vPrLRe/Wr6nEdGRVDuj
vutRkqV3GZMD634coD442xwv2/92aO066v+NJEoxZb0OcjfK2ELSawhtvEKbckP3pKu8W3fMos2o
TFOzo0m7rS8A3fszjVSWYcIu13KNE1qvRVZm6VyK06KN1PQksAdr9L9DpwZPu6synLaQ2TIYvJoT
hh7CN9kw//0TpHfgk1YwlMLD82OXiOoaf38u8f+QBuq3wLKMdk0EKcJbTO0PCaSC44onWDCAXshh
d39izuWl+4Fzv24QtnNTl5ks3CSiMpEfY1FVdZ8lT5oJDrtaTaFpIpGa2z/y79O4wK9YBMBPbjUD
ejCAKxB/lmY0ixreAkxKq/8JfgLHFzAoiZWnx59ZNuFgDJbh5ZF60attYiIVH+YVbJR6Ex/9VfVH
PXqpNr6RuhNBSYd4Sz7O0dpj/NeK7Rod6Vdoon/MSBSe6rfbxkwoyHZn0qODK8LnOka2l8q1AkJA
7DuYwIjtNeoLCpy7Rh9KXdk+zY+q8wfXPWz0Wx4TIJGw8izq+vM/DM9f8sJltHgZHGAKPAnrQN1+
1WFvTmLxej+Jz1GfLlD/P8RCZof+NTfI6sy7vTxfoSdHYtxvPb/If8qyz0vBb7X+sYTYBKfeNygD
nR00cWCD5lMXiCcg76eO/IB4cjT2AXKbZKua6cdx8RLXQQ+7AJlzj7z7u0rSK53DgV+ZxjK4U97m
H/9+bmXy7udp9I5F8MhTH/JpXdBIvGNFKWnjDGvGtaTGqGBbbp/w1C9X2LV1pzh9Z6H9TuHamzCc
opHTjAcG5orIPdGBb9Z5t2x3qBn5KcvH0HKKNY8waErkZVrk94QkoU+Ok2cpivoj/FOnbzOaNf3A
P+z9uI81O2ZDTQcjIws2C7L/BzmYOdt9htGTo6nKwxburATyN4Yl1f5nckcqlhqV0gaHqP4/jG4h
/CMD6LtEWj5m7pf86rEYTOKcGZNBgmBpZWOP8KdnmFkTay5L1HJn66T6Q89u4u9CwSia7xmC22f1
fWnaqGaBelmBBxbFhffn+Xuk8+MIJBH8WIGyNDNc12R6UHDGh8XwrksiWIetveMxcnJ2TPrZ5XLd
5L6mmg6PtdvNj5G6gpg4Ty/EiJLHWnefyKsE0ue1jZi8H31Xy0IFYQwRHrvK2MJ5Koq3Hyp8TkiB
TAZtcXx6BxjVpBApHyemfhQEx7+QCCst8Z8dnvpNtFqLLFhIR3MmBaOhEomhlM0eo5yBaP8YW3/T
HT0x+blkIjGje4+3ntNwC6A8YEFxuX4zrxUNFkX33XtGVWjL7e6Ye2o7CEs9G4CGClo6lgDNVlmi
DD2L7dOLzc7zUhcnBD7n6ohB50hKbI2ShCD3dXizWTrVolrAA/UJYDT5XXV7Gt1wHyifw1fAEG2c
gn2eTuk7Jl4joO01izU4gijKZ9lkzETc3xbetvLiuQGIprCxYzv92OAwv/vvmgVK9RTe8rk2b5Lj
mlZBtcPqXfRFH2viyeMLv3zhZJ030CRmmc2WRnXHHq8/InvKccaBzk89aZQRgth3HjivBzTtFxVm
JqA90PM2Sl6gmlOK8e0ABxg7+hSJKHJhuN3M3EUmwEwcg1tcJSRBXL09NTC7hJvk3QRazuEhUO5g
6lzPrAc2zMRNJ/eZuk/gw60AJLZ7YcDYxPpw1IkdT35eX7OpySdT3XuL24WgUbbuSKzn0nOHs4Bx
dRcq77Vx/4NIDwyX9RQJ/PeqDsUqUV/TNQ3UJWK4ELJaugp+Z+etUyEi7DuaVS1CIs0zl8q9L2YU
oSpUB6NhmrmzlZUBoCOxeF7egDFI7HQN4OVOeUSgCNwfnxBpyDSF1KmnSJkhkRwYBVZpiZfq5v2o
A27H6rei97Txx9tKJ/aYaCC3QxYpzD+uYebSDT2SfKpn1jKb1J8AYFufmGwQWnEIl/dUk1ZIcvTH
jL+Duqf4+9Uc9hRJgS9gKM69B85ZzgWR5R3TrlY3TOqhBJqo/KNRgrEBIy+ptQMPay7grBukULQm
KSHsOJk3qjtkCU+HFm2DJ87ODJ3yz1I69yPlG9yxouETbo++RC4f3DdraZOmgMsFsX/ceRg13wZB
PM+iNxDHFHveIX7sHM5XEAw+rwIH704OBSrZXcnWKM51X/2r+QXubjWAIxJku1oJR4pZM41NR+YU
SevxytiNF4tavyyhfLTYMBR/046WNJ5kmbYSu+7ErynXydAQd9ylzBzjwvZYhiljVKl/heIogFhZ
Lm24ScSKfSxfa2WQdIu6dG7dOAx8ozDRlShAVJWUNjsDGyJpnOKIpNxLKLio45OtNnrZPIueM8pA
hTqZ7UXXIDIMoh81uFff6fJ9O2ATOvStBdxrYO2L+9BiGFSpWToYb3LzVotbrFzBByUhb2b6lLVL
UfOP3KyIcYQj2hb6tFu9e9Aw3lI1MKKUdyJF20sYX8tyLCYxamDb1aoV7IpCfhWGGLqHb6pcNunz
FEE67BJiWnvZ2ScybKS8fSHAbWHByax9ISkq2m+cVHKQ9PVeSndxaj7qstwp5ulzIlxiuFHagVgj
7TJioqQ3ltjkXcSOD5IxpCVpltPizBWpXfPbEhZI4p+uCnKTlELc9QujEXVk/GMtef0Wx3F5/685
DUz0wxQYWEy7fpgR343CmbFUdmUJMA0eTWqqdn6bCKxiRfYNvaDcBPVZTxaqXi47Tv6RZg2ZkWd8
Lawhr19WNUE4jgKcfwfWiHGeQUZNQkBM/gX6hmRbDJjaBjVoLkA9CNAVtALnPmqGumZf71+OxOCn
IitbF7AvHD6VwodB3gPEj3dPFf0EuBhreEb/p4LF659O/pPQmYfiQIodGnVsNvKrJgVOggkdmMMj
MJgNvvgY/3SNkaUsSqey0FXpAbvuG8YszyQg0VQ0E0wTlUj0KXVpY7eWdqVZ+xISA1pGhjiQdrhR
sR5gez845jbm/UKma9ZFhtcMpBKh8XAWMUrWEZ+TAblkyoxH59o8HPQr5WJ5u6rtF3mJSfFC9aOp
3Etzt7m+hnUVniAkxf/jlz60/zrGQF2gr9G6jvufQpjp1isH1zsg8kYVu7c+2YTJKYUJjGCMVr+I
QxJ1/cSqzwWo5adpeFicHDUNMER36hiXt/W672LKvPK2u7MZfaiLQMTObmMmCDujB8ab5ZrFzOGP
l2ztYPSakst/kwsuw0w24pHye5JrPlkYqZn2ATS1J/7VSf4YHTfrT+P3mPjAWSUE+acw2tazXFkP
fZOR3iSV7StjjXCje8HIE7rmMC54mekaNuJJ8H4KuHzUENfMWrHpBN3MGxVlLQrLbsJctFIenBeN
KG6dYnAoLEVC2Rxuqv+ctlbfskeDJ8oYIAcUJE6LrTlseWs/JORmJgewrH6RfDksn6HFzT3sQynv
w50TfIgBJHcrMNr1MMS4lpYeQQQE1DX93he1B41DeIi5ISm1ZYWvP5wBiQtub08XLXXt2LNmc9Xp
vpdffAyYWxW6Mpl1UO4sKtntr06J2H1CbrofBi8YcHricMNTotvhUE8aeX49dRtQLupMv7sh3NHG
jjYnt3JT2X8+Dd945Ai2XEoB3LC9U+8pqHG1vrt+x/aaQEVCGCf/wmnxcIbbt0rRUWEE0hekclqG
K5BKHDqXtrXN+DDD+6oyJTX1lTdGx9c3ReiC2qNOyTUFac2IGmAZXUxBNfxUr2nCK8Bdmvt7Rq5O
Rsyt4KbYb7KYH3NMVXO6v1DBc/EdW4StdTDApTSXO/Cy3M//rq2Mt+M3CHQICcTwzjII2hC3lsIc
RbRJWQqt1enqgVHWP58EgkVEFqkUnTKuegmKqE4Owe5HC/IpO++Qw/aIKces/xqqROCieGBVGIwS
GXNa07yI4RflEbyoCslAdhjimzIcJClwIis37WgrAdbw//nkyoUPUgCY47vYpkKygYsU2AH4QzjY
6kX2ODMXsfAPaxG9S9SbXr5/xa9Rp/l7Si8ihqdkIMmUUpoq51YT7FaNoDkSGgtp0nYYd90Q8NGq
lqQsV+jA5B1/Yysp3AsoAn2taja7lgasS2y2zh99F71UMOx5IxKfi6Pr00oj7zOuac2VDy/z3OFQ
ch7xePttsiErG6jT3bJQISbvCD3Cdvw6nncBezWQSq06/NcXjLoti5Jwl3pi6jMiPzpFJb/QcPZK
DGu/larNW++1nht5t88ya9dBMK/xZQToKX1OuBgPl7J3IQslrzaNwa2bNLiEH6/UzrM+rktQs2PH
0Jw2qYlAfU+5rAhbWHbT/SuoIuAwI0H+uzw0g9ulmrtcqwRzVsLm6yeAEOy8j86lWq5Sy+/L5Fhw
y/iL2ic6eLZcqJDjed3BPjOQoP06CJcaUIJvfN8JloJX4zmQjNrV1HNqCKaAIKm3uBcQnLMYD3op
/Wg41r0V+VY7Sz+wtAwMTj+aq1lwodbfWiCHl/jyDlfbBvDyDTXLl68gyWDbMuLESc2rrQBtXleX
rsTB5S+rpjEwJ+3qQUD7n46t3RPfNjzA6g5CO/WaARL+kliYjtMSWNlxsO7CYlFkxXGjkHKlueLE
JC+yl2Q1pSYDYORuOz3qR9X5avUKWFcsB+wPvTsVa4KQk6u5UxHcJRNpqO5oyZC6vLGOHauBCoWp
V/4yAHDkq/aWJBC0jC5z+PiZgMXcd3F/ofaE4WVitBrQkFutRu5XH9X04gDUCRISeXsdwwoLqSta
M/ciCH8DfxdMd1ElfvMVLAYkQC1ejVpipe/KJdUUtEgnlAYPjtiWyaj8NTwJqTnl1hlBeFI9WNKB
RNceh7uUfME8o4i4tW7O0qxbOrmBa8ZN2uwupdvEF03J69rXxjHv/mT25gX0zpCjGbQDcSciUGfZ
HwteK0EFVJVQxHflR3dNh6xlFOESSQFNfEY/pEc2fUFUxWnQE0Qxc7fm47Vr0f8FEZMqpES69M+W
AvYQZ6LJHpOmTjX5h4GQgDkrhhuHzaphrFpzObzT40FvniyuVXKaBgEi358/ayFGkTYxNZTQZtvd
Kdo+N/D06BCHMTqimgfPST3s7Pjuf/jk4LXY3eo9txotzSYwdLTDKGXVzIWy2VeHQnNKYYs/Zhkk
5WMGw+uKkiy5tRYBtcgcRfp/l0XRzr7vFrNOYK4pm0uPPGu5XVb19aP/l8HXTU9wEVv+894nWyTD
hgikxD6aKzKpAjJ6hwR7mWeZyf98M4b4hSnqbPtrdDWZpdrt0jCNuf7qryRvmyxVP+gwNREhaX0v
PPF/39wvKq5bD9OxdjbPyfFhXtj/v5nPX/0aybuBqfoCYlaBxPgUQy1xI4iBXW9Bx5VHON4RKFET
ZE/PwlqdhnBILHehiLMlOrU1fiM2h18QSUCGcBFPu5tUKaIiWmPPovqx/NuJIUtoYbZZnSaQDP3f
pivtFJr+oH7Z+k/5/0IyEqMEQi89FeeKcBA3P7bKcpQlxl4HPVmZJdbCvihaK861rjcjYNGnpkOK
jLvcEvo5Dd7863jnX5FySnGMFkjHAdAjm77oVXub85L5QRww9Cg5RFrd9wo+lI+3wd6vpcBZeis7
pB0prPcY6hjMfMZiLd45pV72OigLwC2wFVIVi/eNf7Ga6iqQR56M6JM75enp/buHKr43ZLxkx0SM
UMO9nb12UROANzRiQK3U6LuSl3ZYtPWAddtO0At+4Luom07xNyaN21EvlcuMGxJ93ov1NSM2IVW6
nGHd7iDRrG3bgp5Pf3W/VmcIwzrVAyDW8xb6oKV5+rXGVfS9tn8eylHLAWoH7L2KQSQwEB6lTwcj
v0bgRz/5vDjZ30K+vYH6p2xOjlfVkE9br/G516v63EiDIbZaOLQ7iHF3E0LJgytVMrosQ+zBw/Q2
LVwMcvjRDxkhSAGK1yaMjRw4bLUEYpuB/w/OLIpS8lRkj5WNAI1u0CjA/KbEtxmKqGtkHkoEROJ9
RqGqLJsrT/5Wi9r3k8LxHjczDJ9YmmVj5j3nbWQG/BS81SjAGLGysF0X5K8QmHzOGCZruql2jZs/
/oqMn9hQ0SKH3l+CVL28RPpltGRxWuZ1hmmWJSCLmyRD328iF7dehYqYIvOTmcF8aF8Ob4g7n9Mq
AGw5ziaBlCJyvp0OHX595fcvs0fRywvSw/qH7WLE8NU7bDeB1f8klInlnJdQLXnVPiRBK8iC3MFm
ZDpjRQQv51Mt63iZ72w/qhf8bdLZ9hdmxwzpBiiobBcI0QYFWrnO2pzzDxHhAPSE2Cgr27qLNUTo
k61GU21Bjsci6BeBx1rZxket3dyo8FrvTstgRquSxcOR4WCeCG5igF4UZL/33OCmxRJt8VhKQ4kT
JAzF7sM9mtAkwz7iyxTxSY/rWNLWx57BnBqZBZpxQeW6Jd6aZiyjW8gAw03b73w4HrbEueJ8sEKg
FWs24mCyBLX+ZheWa74a2Yii89rQx4VSwCTuZUojh9CgZWJev7TzGKu1XauwHjkM/s8Oyr+1ZiVy
+ndrDqLp3/RUeoC/5mk30hAmiqNnoyGmBaOVgitGCloQiwtKoXXetzoLg7D2Koqg4rG508N9bhTV
039i4wlPgpBKgKTHHaM77QBZX7Ou1UXlIPzocjXQlXa++bGaObn/GYJyHhtuO0+tWNhyNLwW2ZUp
g5RhnpuJV7+Q5gvp7uYvUNAEvfUXReEcBRIgkht4IsMR3SE7kjfI5wCyqPgcfaQF8PP1xh7xceQ8
UegjFUKuLeZUdEDPZZyNvBUQW9OVb3bcK7bo0SPgjqCakK+EpIOI/qJjtFPZbZMz1co5+dc2Ff4k
gHnFtxv0rzY6MJdVwSYbGLwj/SUTJadSPQaPtRLyQB8kYc7wQx6A1mzqTmRiMXtL58tXILCmE/4T
LpEEsgkBV21gDmQHxSA51mFM97y0HHkLizfDmTec8QuTMKQ/jB6CUI22rqqiGXnDUVDGiZ8fF5HR
cBPj+gCt/QUtiiwbSF2oks/fYLL2IABZ1JHjhjSJ4AqdWRtO4GZW7keA384OjX2jQI03QjIXsYlD
AFC0kLrlvDjr71uHL1MEbeROy9wXRn2HfuyWb6OdM0kLL1cpHWjDRGIjbVhzRcICcMgtB1UQM1ky
WSYa8c7suH4xjSbY9Y8LC0r3umemhiUOyxl3CT7d5boBFHT8H2jZa9qGulYaPIBoQaVZMABzyH4r
quzO/4vLhidL9FrYZPa6YQgUT1j6y+f7mrnEXshrm8JpbKhPUQcDonilLDnmjz9cohGRndL50ZaZ
NIbLP4J9zi80faB4fOEonhhQKNh2TSmPYZ7Nn3JRxsXvY5xetuxEXRh24gH76xT9sY/5NVI/pZKd
hc4bZagASzrgVLSFoNVHqh9ggscdb1WWch6xpyf64BrNzDWq0J/PaJGHIdpDx0zF2g3aaCWnefls
YkY0MgxZsBWCimPBeHbqHtEVTT4YFeT+KNLUve7Jx8WUiDBYgM8rzRBH6CWHp0Bx9V5enDQICmVD
INnx2cWI4FAMf3ZJvI/OI0cjApq9i/h6FiskvkAl0q07eKy5k5M4lKfY+VER2OGiLdJvLtL8hbAx
cEVMAEv6HMIXzo5GPQ0qQYyRISXRZK3YbZ9HFykEMLUD5JN2UjNZ5po3Y/eSczhjePg+hIHpQlc9
fyHYO2B6cptIj4Q5LKVwm9dB8fJphvAZ9p1yrsi75BeYPT6l6jTGqr0D3gyEPuZ3YmEzH2IJfhuv
7Gpwuom03Mjhe8RCUfvgCQnA/Mh5Mh4hCsC0QJn5fZ5wvK4u6sRs7D28TrxAG1NwencigOrYQuNW
lIkV7W6+IuFscYpykf5H7Zs3qFysfj8km7ejrrlhITBaqltr2GWnsXtu7GEIPs4AAwsRoiFhK15R
D7n+UGCsPchiL1sgC+m45ZmmPSGmMUD1JqeB7Eo1gMqafjopbO1Rynk4tBEEDm7muZOJoatdfWp+
dKYpUvurXxKyPQoxNWFXLKyd+sToAnzcg/yBGdv/HcbC8bos3xcaN4DTYHDFLhur+mAPSGAZDs3D
VzTg6ak8Qq89KyE57ndrma9mrvQgtZAp3HyFf60aXZ08VRNfu8CinxQfpAdAwIo4jC8KAeoWABM5
3NpobpUyqWXgRSjJLIuWd78cWP7ZrXxGRuKvzLPVcQ3evpvHeS+wGPjfafF2/0rT1lZHFzBn7hz8
F14bRgJ82NnWDDG54dzHNNIomW81+n8Ro5ogiDKYRXOF06H7I1SLcVhA3dDvbTD1LSVUCMtNb8jN
AdmEJ6l0JzqeYYEOYTf6R5RV+ZcNO0/WfZQ6kowJ7M6LakPtIJMikF+gu9vcONM8OblG24JI7UM7
+pWMfgXmpyEzSxDbcyElvDPeR/IUGaBUMjIRLxOWBOVDbAP77in8fCsTc372GYzVykI4YUIwJYqH
Ii0S5qPl+lAieCi+pT5Ns/HoMOipVG+VCdTTBLvB6TPjPNdW7C3DzPv05wH3VOubJJES8I1nX56I
b2+TRxOLaQ9UyG+hm4tCVbPuc9Nx87tWSIyZgmgtYs9JPW8orijS+rW2JKzEL3BfC9pv2tDqcywq
AkOksdZBvzC1CycraCkGQzmbpw5S7PK3Sf0nfua5fgpehnYiIK+a50qF63YC/xzkxDApMz0h6Q4J
7hVpfQMtZSD/NZRUNb4CuFiWh92x0oXpTXtpSC749yZw9DU3F+7P4M7pVgwNXffpCKJd2yBroGRs
LvxXY+L6usnHCr3Nr+Vyvz/OAn7c/JzPamHSyyblsL+FhX1KET1uqpiS2PY2aIBOata+2YjbjwcN
Hz8xWxNgRMW4Okg90mB8c7tCf4CoDDFnX1DaZ3/wmKrmZVmUqmcuYiGtwQnRGEaxMz9k0uVu82wV
Vgrc09whHimP//05HuiM5PwoSdn+sSC2glvboFLGB/dVJcCusrD7ZECkWOFauUIJbRrRuBSsyKzz
fFZh2kThsZyEetSub5/SAYBsISB4C+2el61XUOf4d1jzk5BjljTiRp85K6nEjSbMfltMxxRh8sl3
vAhQNGdO5ppmea/F3grfhIUWjvVFllAdQYtKC4Z9KA+tar4OW6UJPu40c3H9QEHbUiCRPVXHqjUw
X6ig+nwzfrD00hjTCJji42YWmsvnjNsA0amaXn0GlDShdMw7Qggvq4AwW7GuuJjOdc40S5lkqzaB
laoGCEvcWlfkDaq7XRIw9n5sG85M27xBVgdcCeGDb4O+p4ibwUVvHnSalUCBYlv2ofNEUzo4cFgb
qjkXq6Q/9P3R0p4LoC07gcp7do8Q/xR4Iy4y4BpYw8KFLOpHI+M1dRmVmNdnh+3LwD4sQGUPAKLC
cPMT0lfLzLjMjNAWlUlJtMPWVjHPPoKNECcVrXh8ec9tWGBV4vjf9eU9ytRyJVLBQwJRwhrPPo2G
SxJQsGcCwZFO/g3sJtOulSptCpqWvT8N04WKrwM/5Df87l6Va+Eol0xGKE/DLqn+sNLfEcOCcTgW
DzFYyd646e+62hPKN22q5tegen72XqOSHyn7uPZFJLpS2Tj8DxnwxbLPEBlXJEbo+jY0o5ruVTPB
nG2opu9+li/OTdUh0yszYymwd3/vqxNVMuot7s48nPQcBfiv/LokjKVU6wJqpFMARX33/ByCX5TD
Y+CnW3rKVteKhH9cGz+wbrCNI1hq9pWkkuY7/wBf85Kryj/fAz9Jvp8ozL6i8xAKyicNB8fJn+cs
tdCT8adfab10JwZ0Jm69zUQKCePNG0CQw70R0q0oTwqtil6rB+RtICFA0FW9u4lGSOpnyte65XMq
tHn3lC9nQt9yx09+7sA1O2DKDPzuBS3BzjvsOtlC5kZubDDWZslnOl6Z1gKsxgVsnPDpagocG17T
iEnGm4azuKEaba2p7uRmjE7HTLGPMB/Eys1ZuSbyVLvQ95SxHfEnq+ekRo1c3vvlwG8TAF3u/l8L
pkfdIn+zsnOPP6Bu8z+vb5C0js7Wv0/DPgw0E74g+Ab7fT5+dGldvOgvDIrcgPOXs8ycRFoLOAJn
WjhoVkcgEqKwOLODfDKWk1lIQHNJrYkNTRqIFQoi7Vie7++nroac9EuieMHy7Cpd5SnNyqNeunzb
jvw1gEZyOaErf2vw4IrrhnA/T/YJl11Vxxw/S5TzTj1j7DUVid9Zy3/aVo+g7ITwwBL0YzKiiHgp
dGh5zY6BraaqUhVQtd3EbZes7Cny6wt256ZlrwjHm0zcGVtPcMPXxZiJfGVDtlLAzSpwjtYBiKDP
gYW3aXTGst7KrLlyiZNyqmJbqeZ+k3R/nRp6W+JyCTxXq1qtXyrPk95iNqmk3BQbu6+2S/EK9xMy
0jILSUhmy8jqhxwG35wGy5cwvUkPz1rRpQe0Rn2v/2iP/X+ebL9G4X4tc8afYO6nZLYFXfkdEeng
cqmcQfMt1otHZyeV9EwKeyhVgPgcYj+lg3C1ScFw+vU2jv7P7hNHppPW8rom9Vc72ZqaJTBCtMAJ
CEA/4p/46I7W6btgKGOx6okDmIhGUWF3NsqwpmIIrX4qzzqoj3shi89SUIeYUaP0STYocrLOQITq
NVa0m0uvagPQy49glrT5JBIMnYaXi2q15DBSpoMIgMYrLNAGqeujQ7aktMT+rbDfXFjO+/DFZB7n
WeYyDjVOz3U2W8Dy7QMRJfjVrDQ/hmIfHgW+xCwtLJOf2sL2MIiYNKaW5B+hWfp0idiVp5AAqQ3P
6PqLiKeTzu/LjD+QCmFBKprPpGGkuwumMqz4Zh585pDs3lF1OQsMcg0fM9u8eUzxdPTtdrLCQgW2
dNUJZ9scoo/F/eZ0Lnopi3L2dHCI+BOQAZv91DFzo/VZJ5r7XdrJdXhSnbCY1s3RMQuvjb0bTKex
ewWxweU5H1f/wNDEBQRlUvYG65vZsr05tq+oqy+5dXc+ioHb3O4Rofc/Q12bNfeh+7ZmCRuD+aiR
N4wIQTWjJ3vVLb/ji8McX6ODWCM04p/x9+DU1D0JU07e9PifWs0zjarZws6rbxal0pbc1ojTIuZm
PvUX5nIqLSqSf3cpOVtisPg5xwmf76RBiZAyVw7p8TFwYY5Jam/RBVahipLDQRdp/B1X7w8LPnpw
XYjnj8fiTmvHxx0xKajzZa17qbezQKkjWvGbSUegtm87veg7BwBjF8PqW5pXFgfzgkQag6iy3Abv
XFtddeU4CqVc/j5NHIhvFBwXD8GzFXfyauZQt6raBXlE8E2IR6ahcIhflUadtf1G9kUlv8/SF1RW
CexdebHfN/Gew98Njl9W009KpuA0otAeMEocU1huYFK4qXRrGDhXyU04NfU8xtOF0owm2PHvm+OF
kGULRW/OmRtLpcnZyq6FoJpqryReccidR+Ifu04LvQPdUZH1tsl9ckfbmIO9J4F/31IG19ctef6T
4+qsyZ4AruH+OKIamK738kBtcqh6S0F5X+wzERtLtoLETHq0kOtlRDRLPczo00nSgNwoLGOTiCb3
e8U09onZmX0lcc2roGa1gUBbzOMF/ra5EycgFOr5GgTI0c59y6wRmHSRV7vICBHlA9H8YECiOYTE
zpvDJkvc/fQqntSJGqFBUCm6B9WIv+mfMmEchghRM9E4HdYUxKVtu1MepJ3nQQEKihA7HbzSd6NY
/x7DaG5ifcd6IF2mh5ywfXqhy6PFkhS8HZykw2BvfI5GOx1GQhBdP97UKKdG1Gw2SrPnB+ZdHo8D
ns2dDkWMjQOhm6SWcEBwxlOqZjgrjwJrpfEY8pXOUtjIkDyn/Lnsrvfiz+ryzmt8X7gABfUmpA01
qkEX+Jni22in1nteh819pvd1Q4+BQmLQlyDXP+T3mBQfZbhZNvyck8DuObuNUUfZ5Y54knHxz6SR
fLNgZ7lcv66XsSAA7ZA3OXbyzEPoGullfe59fcHMb3xTd/7Skfk2uuqZkxOM74CSgyvo58oiC4gz
HC+gmMLEm/6G1Su7Tq4tTdoGwZ/YTLa2bzGEKAIC7l1okChKR2z2npiquGGqD9ABXS6qMBBONxv2
iCYJjdIC6t7PCMQ1VtN6ARkSAYF7MxdxlPBbtQ/YLrPv9VLjYeGw0Hmf72ALKqT0CfSirEZifnhg
8hpt8JveIsaNDm2Fp8opl9Ubc4T78E0xeLqJWgHd+X3OSuieO6I0M0rDIyARalrWldjKpK78TEFf
88oZbXYqAwPOdEJ8yQELYF+j+Yntp0RGegRYEtvc8wvd+tAa4cfwGEJrhzRZdIzeGUZqfgVtJgkp
XGvtL+Vxow/NmF44aFd+LJD7rv0oMjpkjRtHGJFh2ZGmSp9SxcNLPv0RtuJuxKtf6yuKcVjYYIH9
4mFpdq/0BXoIwaqkcBWkAFnt/7MnNEZ0bKxKTFhLDYCf+G9uApYQ/288i2Z8HQTYmV6YCf1uR20m
uL1lMtYDjAMzwoQyIT/YXnzHAnmNVPqgsKcgKPh/S1qtZluvMIbObeUPeI5XWUQ9IMvkW5QDB5ln
MCwPH6Wq0Ip6oMCHBdcYNvQ0ZGlHvKTv2qgBSEjbL4oazpwsqAPp1eHV14G7UhlA48n8D883QhYV
bvo4KgcL+nEVyxlsdTvMwAmZu0beXSyq95xicuG9KAPbOvtqRHpNTuw2vwNelZuytQznGIksfwvV
JFweftUV2GKu0WR4rMm9agOPYm3uq/XRIZNcEAMdxKh/dkrQG8/XjQR/bQFWj2nXTVtYxxS13APg
aX05oswrbZcy1KK/GfMBcshNTj5WWWaagTXqWJTpSdjWg/gHdZH7uDRMVU9T6fXX2+f90Jo5EYY4
EHy9sQmomwJMutKU4XBcwV3YmHgnVpOp6ZZz/kcNSgIwuWs7gqI0bDuh88qTdVNIkfVZKxy/TnkL
vf708rqi+x99KYbA6M4nbRzqRjRi/IDofz28D/DyxRcEfEbZAyByegRKJ6enonM07fXjEoRxGir9
LSgg20C7UjRGO5v1bm/CjFo1aA+TJDls+Spb2QnI59V8XDxrSz5/drA6+sCW2Yp47uhL6VYOT7Pc
nUkKM7Dy3kZkj77feNhFTxX+aIvAYBXOZGAAsZIKmwzAbnIGDtBwNgzIyIOSiX+3EK03yP8H3Fpl
mbUfyHHRG3VCeUErRqrSyPVefJryddIkeAjJNkKGy66DRi+ovIKQ/CQmgcbaR32cdXWGSZ75/QDu
p/VodyhbYPQYm4Ej39FBmPXPBmQQkV3ZtwfBT5qZAYVO0XSJnOjXo+NCsL7Qk8B2R7qUdmY0K0E+
dFpjV2UEaMAN1hDpIosRgErPIWzLQp0HgLJnOWlcDjI2DIOTe8KRrv8AChlL5JgTiA6ig4LERW94
djWthY1X8ul/WddY51fUYklXSEymT9ab8ZT0zoHsk9PVB75OcM2rcm+DX6iXip7lqF3OrIgE6ZHn
M/3iAAS96mrnuE/b9eEMiac5LKhQf4K5iSro1Qg/t24qMF1DXDrFu4vbIxX5cNtOJOcglj+Lw42/
lzqfHfRHksNfxNxSDuFm3+ql6CqPviVbyy6KFd0ZZd4yXGlJ0kGEbq0hdVLPrgfLvUxu0HIZbx+G
kmx7pXAldy+D3zFbzqhJytPYNBudiXXNPvJS2cAohR6hGFIjvmiMXwlFQZpZAYfsy3Q9QhCbsJDw
bXOLi5UawmZWnB97CtC41bDgunM748UbWfMgZYN0ALK7cCzopAJ5QjIEeZ3bqeSNOwC87ho26ple
reBCcOqOEOrwN0aVl7b6uze/LA3/OY2Oy67gVimzG6c4RHtu29HllbU6ED9Nm5sYudrc1ERapVvJ
BHUO7GdD3iM1ngZp+yTFlA5lmSpaBkzqNt/J6WQpUfqF3zjGScYmbJ8/jLTPvhXGcY/XaSLYqDyU
tlwi6NZ4JWxXKodKNC9USG6SIVFb8BQvINIpEuukIIhId75K4i4zOeGMQzPPAEeFUeDPM1mA8jHR
Wfr+3sQQPly8bDG5KzRlK8bNaU9uvhjFk5K9t4CLPtahcJsa52NkslBI3HGYL0BGNBGileTPmnzj
aet6/ianSzG23HxY51j5JoedeQ86OY6QJuyQ4vtOW0Gux47Jtc9KqppB7F4zz+C0KhS0cIaCMd0U
alE8pFSIzR/Uc7/6NOQUg8f64nxXKJhuk+O7jdbmShyfO0CUK3fNnz9ZsElWcef37gGlJgcfgOLQ
34mgNgcGtKXhd5m40hy5jpfjgZq+ofxHB/mPbqGh/WO6MbeKDUmGjzmaILieto6ibuzJfjvRrmte
6L14bygFm4BaOH1o2vT/xqLcbC33LYKxBo0uCH3r0+VbOl0qHck+5lzL5L7lKQE+549o9r2/qxzx
teNanJXA3oKOlKIBfpkFiy1i7ukYmM8cxWSKouVpP//KyEyHvHNjnGTode1z+c+FtQcbBnS7tkho
3y+3pQoVtC+rbaLygfuVmRbzsgbkHeK6sIh0XDJLTN6uujye5AxAyL0HEtrq5mzDap93abauqJkr
4iXYpUKJZhwsrWarjBsVHdFwN+bQ/uNrG2UdC0AUAdiBpEEBAXbA8ECYvMhyZPU73egx7fgR9QjV
yndJA/DhkvboJSPTtDX9M1znYY4Bo9scOQFIF749YtSk6BeH4XSRBjLLGdnTE8JKGC3Q+uvrcmvw
VwdYbRcY9lQ1SBiACUUBWhvxgi3cIkvmzC3ZIjKl6GztaIs92RndN+54UcUrVTZwq0Ur2VmqkGEU
/iU8aZ1APa3D3UpLhjOMCASyDo2aice+I6wYrrWc5mXf8IiYWUJ3YNJsXE3SsvGhenioplMArwDA
hYGA+H0N2E7Et+OWpP5DhF/oD3ByX7T7uQVZYZeYXC8N7+GJPzQrf2fa09n99tEON91SvevkhEui
1LstDv3evcDeZh+PZO8X0Eu+iMV62nj6P8nssM6saJ54uUTIXN9WM8UZOdAu+t5WQkCIpwa8by9p
DkWKQ+ZqGu0qnK3VbGCyfOkRYv9GAed67Q3kC42jrrSyhC/x0TNO3EYU1s88uI6ujgVNOskM9F27
ZupQtv+CaHhVRkQj2bb8avk5D8qk98enXbVYYrkTzhjWOaLbLUK06ziqp73lys9clrhJi2c/K9Ka
72GZ8lQdIVbOapjT5yElg6MyPpCM0E/AwBgNf/qfFo9oU1JGzMZu0lxuVQ2lFS+FKVZZg5FGPbQV
rgZGBS/LTyneCL79MhQeucJQhHrIN9ey5kgOtihP/nwOj9un0PqQ7olFmq/jATNKz+2IWE1Yerws
hEXS3IaBEIBCTm2APBrdHxiPdUM98TWmkNpv11eN3i1bzxArIIWyR3SeEtptDKV6ls3QMEFyNAxJ
tSdFQsRWTPQ9FyfcEFg4rkT76uzeouDlNCCJ+5c0/DD2n27F7mfEicfxANdNFSAvw6G1kdHZeLxH
aTzHIp4ICyBSL0Ug5jB5DlBi4AB+lHByKux/ULwAYphpSURSW3AsHrIpm4udQJsVBXiiFFgOmxDC
CPPgxIfPxbx09WpTk0YD3ipOeoLFdQNqMqMMrm/soSO/Dtb5HARquIjSKVDiXW3IlvdCqlejE4ka
uWfOKJ4TAbJ1TJ/IzQ8B04m19202g3t9SxXP5Eq+I/Q6Kaxv6YH+ZHrQxYA1ZFcPgR05rUuDqUR7
3Vf3x2ROJBcl+6TOZLpWk5qPaE521vagMxAVvXOgSkkzaPOBVu1Uy5WHiLve6SxLwwXCT84gLUEZ
lytfjFLhwaade2dbfj2FKVbWWI4ULCV2LT0+umGy7IRXPid+r/7FCS30/U8NYnWq9OskVlpFMtkt
Fo+HBI5PbZuVb2B9rIHNlE5xukxJRSCBmRk5E1yVdX+/9+qMKEVKxxbzZlQ9FB1mxF3HLaJ9eMVQ
xY+Mw1xdgEBIfTtVb9nPRwQuNyDfHOUeoWiOeFIvDMwYjtVmgq7eFzyhAAqIj3EuzZLMvtzQwrQ7
U2n6N/DYkvx5JA5XVLnfMkU5B6m6F41MZHS0JrgiCmEHeQLJtSf3KTbN7TVBU/UYEuHb0Gkhzu90
77EbJVluGLYWpGX+/nvVFjvxiEJQB+7bfOcFQowJ3t1b6M4Ggc9aUb5Q/kmX2b8jxyho5ufCoqgC
PQzgbqZ+KY3ubzLEVELGn4Mpr+KgmDcBjKeMfXPofCDgUm7BilIsavRbgs1gaXFq078VtUm4cFo2
PUD5wzc/e58i1EYrB5SQHTpeaiNXnRaHP0LZ3yYkqfC6g9wEwgMSt89LH6K5JfyFm0g8q0YzK+wI
WB2rk4iwTu0sIY+fUqqtaqThXhZBoUvK6jsEKBG5IlAR9Dlfq8lp/Tr+MFrSrhgN8tXHpTIEJ7/5
XAHxrEtBBEgSmskbkeMSF8CuACH2lpfiP8BE32FZrqRKQF5y/idc8ndPSJBqCFS2Xy5Qg2ZSVTLh
lU0owzDU0r72was+WWUsG/bOhiji4Dhsu3uwbKmE5sTDAQskpvya+d4FWeWjyX8xj1IolWPzijXO
7ZyYr92qQ8PEDYkjSqD/g1Frha7RbnwO/KH9x89Se+3xWZhw4T0zOuppknssB6qDN2WDM+LSqa0e
FovtC0m9TMnv0h5euMiXVEp+s0pj8rJeW5ZoK9bQrf9EusJhWD+dxmPwzkg7+fjKRtYe+TGZh5Yd
rFVR2jy9denulQiFXXm+L/qnXd3TvrmxKoFoHznVvySgOLOeTviRyQrWbcdbCF6cQjHDv5CPoEjd
NBV1/2kw9FfiJUJ1Uc136cTu5qCK2MkckQ/ypQdlJ//PUeNQAAkI7Ds27Fn8LHY7LPuja5mujEMx
n36D4wf2vVTHc9oSgJUd0FJ/VqdnfGj4Dl/aLdErTwNgm5Ip3yEoEElkC0tD602R/xVZtN0x/5Zm
ZLXTNunbvRdoz3zwZEh3n1isiHBpu1l1ECKoPK66DoSGRqPUPUeTpaSxq5IaGHN0U7r106scrNNu
45pfUuyg9mHRQ5vxAl4itGwBwy63Gm/ObEPvkSIvoZV8iFptcIK8r794Gdq7GgxoSTFFSIlrXOuB
7pABBVLh0n/ANMw0TFWELLxadqj6NuryoCyAX2yjwzTJYyHBu0hoz3SHbKP8Sp7VY0nIjWnHaC9n
QXZWBIKG+copqMEXp0UPnl9BFBxRGyJU7c5zJf0wFhTzgcx2a6hgdXiF/VXuZ/fAxaI9g5YSDXiB
6WeiMFDoNOUnIH3weUaQSnfbuclybIBOCpnfsHgHsvT1KddTdIc1XtuL857vwL4B0110Xbq+lDOz
BE51U6Q0NJ74oonZ+mCN3iJHZWiM+pf0bq/e2k88TA44xVp2BPbRGwyCmfLODjig/FpAc4Ly2Fhl
zAp1Lyn6vMg3eOeFhR6UA0ba1J/tbmFxyQvXosz7aNUu7eP4OELDr5fqcWtIfWRFkmHI57QUGE28
jbss4JKmjfM/VIKMJctv44OjFR39L/TaQcBk2Af9NsWAfm8F6EJidQsMclVqJ5+MTK+/4kx/CKPe
zK2o+tJ2IhtBDa3v+/5ca8OdetoBymqlUtN+R6RFXXfRC0WUDVrDDzyHShcczLy3fG0a2MlKExGK
hQVSdzf+6ffRYEW39yVTz87s8aeq0cVg55FkxsveVbhdLCDDwiICrLz35+MR62d/g577kjYrosVK
eRnqhgMwqg2HKPWUnr9+D1N80tUEUCjr81aL+a6U5eWE1EGC70IpqSUwcn15e6lSYaJWoA4RDHdL
K8ev3zA/e7/H7C1eIptZoq3SImpTGvxzAB1j6V/2yT3z60tZ3qb8kMDTJznZYcB0pKkHCoe0bYeh
w+Sck0+7450vI8O73kEKdY1XaUVsiOK2sNs4D5znCaaP8kFsnwWvIkHwaUc7xXs+iJglPvY45/ls
tfwxp4mGGu0DosGppMZ0Ia9nFhyrr0gQHNvaKRQZ4GpsRXtFNsH0VXejePemGhGVi84nLlFMqXFM
KMOQTCbe8hw2sYALECps6UoFGWQw2pf5pU4EZzAj/KI7UARYM1+Uefw4ci9Q/A5CTNt7K6x1PwWR
guvVWD2E5x8J+2im7xxyPuzn0B3KmXXlynfUWOH9njS1zj249cGAafL5eHfHJZv6S811EzJD9Npa
2TYfkeQctHTu8WZGJzWEOxVvr517ziHAEyNqkB9RJbcBKxq2nVIXBo3LFWKJUUIuQjpsby6s4Png
uks4sbKh/JBB2lN3Dgi/Q2LOLe2iN0PpNH+52ZulpCKHcJGVJKyJJdYBE0dyLFRQ5CkIj3oxZfZ+
xZchUyZOqsQY0v7sjLzal/Ohr0xZUWsKgTfAh2aJnMWRpuEZm+UFJ4kp4dtjxoAhdrfa1fjXEzXl
Xd+YHcZkpiKc2uO935JssJH8BU05LhP0EMYsSFAfAoPqLC440L6B/WV6ulZBvgwE14PwQGs8AinH
GV3LsVJv2mcPcILC6E7WDRB+Wog+Ri5nhx8LzcpjnjBktFb0v2bngPJEuChtbIH+uuAKkYFpO91Q
Qp9lEjfxeM3BCPFfNok0SfCZ5UAqbGfP7o3AfDw+RqRfcGpFXiEQrJZGvkozI7knV4McN/zdO0Nu
Xjl1RiAV36iULQMc+9GHXgd82JmFydRCD126RIhdXyRQ43+8m5QA4q6qml5yqcIMPjw0927kEUPz
hkfTD/UmnP35diMSHIdG7gQlcZmGwO+ptBnhetWENjUMHIC4tYIMAJTi1cB0eJsWMJS7o8azSaHT
y5CvUCGnMbiZRp6qw9Uj6tL8J14mtSlEERv8kH81/qbHk2TE2/ZamR28Ce3oxV5QcgojeqITzS2R
iu1mSsDW+jAYvd+/vjMLWvp3zBJ/HXPPR2RpdpgtTHibbLMyeQ6WHsbBq31xKrZ/7YzUNGydFhsb
OEzAuO06HSzeqk/Hy3msrBjPgb2hKeu/zFZt0bcxGV8LgXMpNdKj+98GWHQTStluga+AfWvBpcJr
xLK5JvScW3BWCBKBC/SJhwcAvegovS/B3z8zCsNKfrcgH5DuyQK9dkMncbiHkCeEdMo+fuxQYaBm
nbUYdB0CEUZN72P1vgDpn9p2ADLWT9Op6Q6a9Q+h7Ir+wXwIHoqVcO38KIwI2CYFPpWVgB/DAU4r
qR6KRiQnYBb4KGAlxtiH7J7fdkJq5MRtnRaRGnPkWhJdhcpy4K683AjUPkli2lDFkWTCEKBW8d/N
kGKKHv4b+7DoyDfMuvOKETagS+wyUAU14icv1t4eIdxMExv+d8zsFxAdmBmpKKccJg3w8kh0UfNj
tCVojEihtmjuOXxy2FtqTM+hxWU7zsp7VQv8BCaF/53H1NZf9KoMiPV2lwrGxM/6JxuexNeCeRw4
FEjA737J+qq3KMIk8vRFtE8LoMTkAc8KHsjli1mXkoqDRZcQjoWOrtmSg6gaslDCvUmTE4gKZr+z
pPFBdNvtP8MMa7Of3cXjg/G01/jFdzhvPgU57x57aLKk5SQ82aqXlYNWhR9I+4uS5X5zO6AfJycz
z8bv8jvBHBkqDZAy8SSo19RGhHgWNQ9g2Wi+ImtRNeiyXtRVPzXIP3sJwQRUuL6nEMgDTHEeokZh
eybXEtdqdVZYLmqlpnmae6YSAq/V3YqFCkM15VyQTO/kfhx+vkTk+jYBUJDC8zDGvwxoq6hM6HYV
vXGjVk5EgZsbDA1WIZv8v9eGc2zsW22jZoR9oBkrWv8+IqqYX956aeXkSEpjhAxRo4O61/VQMe57
BEnL8RDgaYgNaIVtvycYBAEnTtgOjPjecVjyo6gFnWDbnDaSA+IlkQMW6ul1hdN1iifye8wbOYME
k6p44sZeX9OShANpQoVurG2mqI5TZPpmLbHwasyEg1kK9sXFXzv8yltQwvKTAtmHZjyNyXQ3cq7O
ps8D3uWOsiRvIGBgNQbz2vzAP47ocnHUmg29p4wfYvaHvxaYhnvRIXrhf9rUFHteWBgP9Q88iTl8
V0I1FWGs5weQWEM39GrIyBjV64wKwkR2HuhIzHvTULg7Wn1z+OSejA4HPE9wlkLQGIA5UjjLMw0E
ycHVzoPefIXqaPzEvPtWcAEVgcWd7uRy/HYVyQAyOlRe5pkTE4xoIqsYmnsEZ87+agPG/i948wij
ouszXbG3uPGCqR0o0OruioCITfvzeGSSiXYwFabtPjj61q7+2XMc+hGThL1603WuS4fOsNF65Jz2
gHYSNyGIyzJAhnt9mtepGT+J32yP8KMXm19Haw0N+5C/D3Vn7x8zqfb9w9p1MP13IKZtPtFi0Nk1
yUhcSTnisQFGlIy6XaBQ+E2XAyuihRk9hmHX4zfH50ygR5XcN8LW9v8lBSEqBU1ENM2Dy+PKvTVf
MJO8Emk3YQBL7/jep22RFEpngApcjG/tol5Pzy4BD4l+yUYakcL/nKnIa0QeDAjATMQq1RVPDMGR
CfYTJLHIKddH6nSbdTROBK+c/2blSuUtI+hTbjMGloE7nRKH3YB1nLhgUbpncxmQcMUsZyUp2W+j
++Qijne/7KKe+yJTZh8TZYr9rcSVOU6o/fPaN+W4HReGX92P/5ZV+NYwfReww4w/6MEGxOhoHX96
vu79Tp+9rIYsPmAQE8dQzKactcw4L+t9y/08udugLCj8GSx2aVow1LMAzneFjBCKTLIDP/+sKyCf
z0QOvKnBdYWAPBTWOmLHJwijRCec2DrJoB9+7FYJkhJCoAskoS8QcIkHrJKmnvoq3uJnUlY90U1M
WFhhE31u3IWSGtktmLH9+VXF2pnj08s1L/Ed/U+ZmmirgcWBDfVN6rqoZhU9OIcKd7CHvL1mbRbj
w0lSqwbpiToS9rW9JI9R1BAlt0vBzq1tHvAEGoK/DTTHU0bg0WI/ZklSnRrU5m+IvJH8QIwwp33N
YI9P0n6K+rNTrE5YLndnLY4+49+tgmgZI1wPeB+M6TI4pZFoYR2ocdOpHH6qZ6yW+1H3/HN8HaYi
uLlSNM4e6qyLyOscHUiEq0ryKv+/mqhwD9vLNVg38pOaL0mEnKiYGYp6ajOnc2B5CPIT/KL/YYDo
3vzbZkof44lB5hqiPM/0KX+y+wZz3j8XraRvAPZGhgivvK4B6M5BF4XCR0JYFvTqLvfYZX0Dep1p
uuLl9JMRlzErknwN05dsw79ebNcMEZYHVOekiIk8UawQGsYosjYqSMTqk23fexOqveyNMx43atA6
RDCAZr0i1cK5/lAzLioKSSb2bnwo3SX4N4C6puLDxnLFxiPEXVpxgUwSfB37RxMVF2EkPJJ128Ai
HUjoOpdpRTlMj/DpbxcrY0fMuKixRzs6UhjIfKXUbo5H9wE1Qtw9TZk/YTml/6kMMKNZaAoRro0x
Ea2yL6R15EDx6yxdwsGLxYGwC3G7wTb9mB3uhg5ydZx/YI1BL7yMuuDbeuHMv97p2AJTe9OsdA4l
T/o8vl8laFxZKT8/8MQVVNVuTOIE21/I//iKOzLpO/8G3gssgHeQ8bxl3eWixM6WpvxRI8dmiKM9
zlp4Pmn4IpUS+hBaLi7GM4NeL6Oo867P5FiBlf7uKUpA+x3N4bOO/vjok47plCpKJlyLrX6/uTTO
AXwWT2dbbPOx/VXvf+0EBZC40yFgbDetVx23keAwt/xvHn/xTolFmo2ycX3CxlWKRsDBJAOL6Gcy
KxS74d9WAYSpdXInPRk6qVsGY6Ke1c8ZK/rFaTjJMQZ2/bO5RMNz81kV9snv9QDqnfEJ11qhVSPr
uH/TpSJ6qJYh2iEP7+SXTATIAAhXVGOq3tLhKsBSyagpt9d2hAHW9vIggWZlgILPVz8AJ3lQ6Yql
fpp/mfm7WLgNcdMNpo2EAXDMnUuZU0a1+KQ7DJx8qigddiaWfBt8f9LCRQP4duE9jYK9vkQbZI1Q
kTvydUl4q44cxXNAkCzVTaWLWTTx8hAtCsEBNXgrIGx6n42IUUOCXGfYUggSaa9As1Zzus4yVL3K
RIWrllkmVlt1j7QTfTFj2Yu79QgZhhZNDrbJQK7iOGNydJ+xJBjb2syx0mcUNnU/PoaYUnJ8Rii7
xAiwGQ0OJDNP9szk2PNxrqgalyxJKlmx/tMC7h5iN18ipj9dXQxlkrHELgGZbN5oqkJal3enJBOz
3QJ0wKEzgT/C2l13QxfhgZ0DV2LoIy3mN/XcKOJYSxJ+3wEOuOJb8edrgGvtheei0L0Tgl2IwaSR
AqD31DggHD7RUslPWOBEYKyCKhBybYBPumJXhg9cRskymqIBJlgnhoObs5Bsn/1DBQ2AO/0lIr4g
LGczy9zijZT3iy7N6mXQ8WbyNeLK/Rn8J8zv58l6QLwaLS+PKSHSJ7jsWPFh6vczIK2Ll0cNLO4f
rwwg4Nh9YRcBi6XDYKSR72JSEURuJEInvtxZNeWD0A3vpQk6bOGZkcnu+2oqW9HGCtOae4yQxhSk
kzYrwxlAKnhoM/p5YDgyukf28dqHYx+peqgrEZKxdoCn8RxPQeqgiS4Y1/HLzqesuO4XCmwiQfGI
nSI/jvb0gV4OTkeseSeO7mHIoIUPha6LjndCdb+zI9vgjqLYNrPKlOa+dBaNu5ANqUjPObdRz57i
aVS19CSOKkX/CRdYdJyuJ09n7WcUuQWvedeOG6z7bcVuDJSY1L4NzBNA4is6UK1n7bS6jz4famIz
iOWO0qBXp1BAG5KuCBL9JSVc6x5CbcGLT9XSbikqVyG5BFAZjGJdiisY2cNJzQzIHfL0dkjBhLDl
Qwb2LHS1VyrE/h9RfwX4YK1WduMPY1WZU1uKQ/4FdnV2drpdntoAs9nVLZ8O67tVhvCwZE28oI99
mCE8v84jaU0yXJXFh+dWJBJs0FVs8kvOMuqV5Hj6Fgz6HuGPX3Dpmu8qwxUBPBdkU5HnhowEEykw
aqQR8z3YfKA6SIoAlbjmrFcYU98DLBpXyeg7JfnScGyDYl/qiApmTlLFYfy1jCVOT47jvha0wyCZ
tfzJB1GU/If2v+DM0jWVWQtHQIOPjcmu3SC5lg5PXB5Qt1S3gT6DzWYqmcCvaPTsn/WU43wVrViL
/ZHJCQ8SvVt+AHvVm5sCKxeuVTfycPduclgLvBWs19JvUXwEl9Daf+lIacQhv2w4JeMiVOqlPVmZ
o828BFhtMID4vZmD6OCtvMcUb/VW9W7JZe7lkjVGpPC2eqnsHs5/htGrRId9jMUphJCuwFUBshwi
sVmFIF3JQUx9GBK48RM0rnLnkJaqOyZIe1j0GXF3CQQ2xs4BYsElhO4W/HTdgGy07JegzNC5mp8a
bZMLZZlmJrexvhB1ZMVmgPutHWBJUcl//ZbBm9vk3QVGVmAgfKfWU3WVDyvyep6wb0Hov7zbB59G
BB99ACCYBzpnF55IyzBTnIeRrifK+Czh7gjFJWxFBMftmW6WpU9cVQ3GhSphEFtavy58RyCqO2mu
gJYoCJQL7lMHCPOtpql3rQGlkL9312/vxb7118L7Up/ZFW+jZXjmaAG615QoWutuC3lIzT5sDKLH
LrcCo2d5BLnpOb2pGx0Etuot21631/X+dL0hPN2Q0ph8iv93qjpXTXM25K/KAYpBgBL23s8fKPgp
a9YaMz3me57phBG/W6jcCe4G/QEDi+/A7HqrbctWZG//n16xaK7eYu86MKTo4r4kQKkYovf8fCVX
cTeie6UZecop26twap/p/gQ3PUSTeY9RVK/xoS2KuFfM8/XUCNtC6D6BBj8aFxYWQg+ueKbgrmIx
FW0f97O7CaXD5OBqb2vTtkS0dHp7LgnqeBDfU6biIZi04TyFRUOy87OeE9HK9ewjk1RdQ7FxC+/M
gqgVVUyfBxth7xLFq8J+09cq1fcDTJDrJQrvFg9UT58BglkZdRXOoS8ekkqiY8fzCJyQstUCoF9z
B4L4ggMaM5AZsYXrF2UPRYj18i0Xg9+56HVwrSdmfphrTI0AXyAvXdtC9YilIWnBND84sjO2JcS7
QnLdHtA7fs38+0wyPqCRuVi4bneXJ6Z0CAvw2J0kl+GwkFB+1h7iRw3+flMHsj9PRndHTw6W+G5A
JkAfxttZeWYk8+N77RvfkhpYNqjhi5ijespHFhwsJUW8qHoy0IM69nVEA1fUuQOfFfW3SQEucFTR
QsAsRpyiJG7Z+SC/Crh15njosf7Dje9zm4acab2JSC/JJ6FNuWMfG0U514t5hRFuGeZMTKlGofiz
x05atDgyrxu0P5SieHjnmDRHzFgOEtOReK8/TF1JvHKKlxPolmpeUXj2HMwCBoG8Zhqm5Q2woXJp
gFYravXUuAIHket4YkFRJIWJxXEia6/0rk7DQFYIeuM3T5KMv/pvAtAd407WRoTWojO6FX5MP1bL
SmxP/h73Qkwsxr/MtLchKgiMKAuVXI3ELkhGk1x9V18CD0+zv90ni7KVWPaBR7yxBCFl344ZsLZX
nDdCnaNxdHeeP+k6yIQVAWwxOA/fYGMveJkA3KAAe4nxiWqcrt1KQPFdH6FnJtC9M9hfxfrk9ln3
gtXpU7FHi86PX7esOLQNEPboAywb2s8NByDYaIAqt3spiVpVa1z1CaZLILocuixcZ+15bYGOdtU1
6b4el6i6E7edtE/ARF3bV6/6rtwWDanW/TxQgiZxya68ecc98qR0I4vCjeqq84fd4BDDI++T9yx2
auvBxOwWyCqwG/vQoJf5dhFSwwx+e70cKkigv2M84uVGYlld5yLj0rk9RVnBwCBrRhyFtDbmv9ry
E6uQG2W5o0QGZIzru2hQ+Bv6KX/6Fq1tQioXf1/508kEdgYx4Nz0Ro/prriB+GMeOcX8BBk44do5
lO19LYy847GkHRHyS31n6bMrj1COZ0D1N68Tsr/hgX3WF99+/5YZoC4cGX1P550nV5y/iVdUQLtY
WDJSWFtrGJxpsVKw/VDoX/iVtHAt/T5WzM/gAdBohxD8doY3NnF7XjDwjWK4slaLYv7qDQ/TMB5O
LtQYGWGPvhKAjRAvBW2E5oO/1zLdDKJtkCFQIeksJzi4YYSpOuk8+WNacgWarCNPKHtxDTEL0DZj
qU0OV5hP1yuuDNqOKwjpebY83AcFoF2jr5Bz+qKY7jFBSsynznxOBjPyeXAhc5l/2Un9TCa4+37q
TUUE8hjaIyF3M57A9WE89JhV5zGLWyCL9+mmEXzO19Q66o6WEQXHX/uI+sLu365ZB4avXA/zQONq
vq6YMNg7k6rVf18oh9CQcJReYeBVg/ISb94Sn58B1/7Sid3y6oMvZSFFLamqHHF/LJ8VotX+il+R
NgmsOKOAe4v0nx/wSG0+5DT4lJegGoMCEcreioCI79epxgrIkAq5VVnYF01G3PT1KWts7nXWvQH5
8P6vOCzsSsBDStiCbomI9o7ctNlz2Ec6T6SGKS+UA/UZUJuS2eIYar+7yvKoq90Z0gsoyvinFXZB
OAaAFq3ZVi3BmfRwueYQb+lJM/0O5/GPU0ZHcEqALQhueVwRfX4oSW1TsCPukg4/TZ94g4fDOGqC
Jx2Npap1e+NbEFnM+vuI51TO/X0qsmytPi19I1h5vx2Sec6JAIZnPYSAc+SXn/bdmrI6w9yRgx8A
B/OgFI5b255CccQlSRBMe3Ac6UN9njZeFCB2F1GFtSZ8ldHk2YMI9C8ddN4GDKSBGCwKnW9gr0pH
0kMAdKrqU1aKbXkQZL9w7+EgVzrF65mJiqAH9b4LlhIP8HOQz+4QWGtc/FkGoMrcWK4U3b4GaR7r
nFCILGrteamgsZuf3o0Yj4NUw8cZaXARhmuC1Ad8/07M/PmW2A5ASESiQop/hNS2ma6/+rJwWbSD
OKnVAcD6rFMhO/z2B/wlHkH/KipvW3WxppfKjOVj+z/IFvHcS7sDjMF+pR5isrxs/k04iGiSHCjE
jxRcGZ+2/FGclTkAmZJI9XcDaQVBuzltHSB7pYo4lRBsBhihJiExlr/8FqL+wTTbugDk/jErulH/
hwH8BHF2DdicEByDn2XZ4kmf9E9kYqE6OnIFS9DQvfVgDndMaQhf5EL7zNlOtPqDPbYpzYwu+sUN
jyGWm8ksbow/5cz9PablFsW7Z+d+YY5SQUkhaA5LGgDufaS7UXzoWU94oUEne2+j8ALsq3cVcMQy
WkcrVuithiMdLTOm0RDYxyXR53VWYhH6Ro9tq/2Rygs1KR9W/fy8ke3158dhYtdG52l8IwTiVWgH
Ms8M7AVjx91ToxmNA+q2ZwTDJfdITSeFq6aTxAVnhKhsfy/zurVD5/YsopKuwLAHANNIYwyj6sIL
kXVKLbuRCqWEhdwcKITbU9bmflDXkxDDast4h3SQEn5oRW1cGzIIihJGDjIyUGAAEYjQccmpLf4B
TUplqhgsiogzlQi5eTVXvrMz6htlMoWnJToQ6219IvLgFmuIO22bS5W78zlEmKtnfvaA4Dvq1+Kw
OMZxsD4YDXOawQ03RxcCAn1pT/bF5vbKcUsGXl/3r+is4bi1Acr52hbFOuKcXc4mKPIlc0bgeQl4
pe5t6roNDt1Hkfzap/fHGV5iQbN3mRbP7zCKRntTNo4SQEqNL/G6T/urjyfCi9VjdGgF7cX5W/Y/
ORvh6R/1lzTXAC363Dorq/f+nm1Es2YQJa7CHknULxg/UuLNpPWdg2IFDoP6U7+ZPwpqnndyYZ5W
OqIZsXxCfzfIytaU8edjb/CnRzurMR+pyM/i4h0hDT6lhYcAChjHDyhZSFGGxBjRv/cw1fm5Djqq
3hXlYqWHohiW19bPeI/k2C9563EdC7EYlhMfJXcI0VhCDFKOdWcPLIMh/5CRPAGqCGCk4oQtYU5C
oajukugCfehC8NQhJAC61aSX1b7MSieQZBDnqNaU0R2kvgv2HIZIlWg2ktcjUCl4WRyzCTSbbLgY
/uoAuc2FVBrEs32RdwHcjXojZgf/NL02sBPd4/zntAoi+e4qwnw/roPwgf1cfoUqPx7R0p2Ep7nE
ToAIYERHV90iARUirvZsAi21hjoolnjydphVaVgnFNC8qvmmwgN3zxTpHFdEN0hZiWPyCGPwLuv9
M0GHcnuU2rE5UcCnTvHjNFnNyiZEak279sHrSzq4kHzSZm8h4yI0sD/0ZM2/ZWnI4vvH29nKJXdH
4Q9NTX4eDUgtdZDsNPTuAHak9/4apjiNFhZp8k3LXIzslMtbArA33B80LTxofqMykZCJ/OQuNNRH
gik4KynisS3oZXtmPOZlLaI2FOyYMb2WyLZ59AhtMTlEeRZM3zzdFVyozOuixrwvdex43+++ebpE
bp6YDnJAdjQxksyThV5eDmthXYof4PXxpvhi/LZF+ZOwXL/ACP2hBiM29q9dyKyc8NfAwVhGcGKD
7jCsqtkI7BoK0JfWFGpUP4ApFJKYdWga2Ga/rz5ygL/fgD5SiMzG9g2i0Vkx1sIkF10n9h9jZgLi
ZCcQ7ZB382kZyhzsypZPzghHrr4H8iuQIwC45K+zlPyxlczjAtC+16p7j48OB7qVEsTVd3+mu0/r
MR2/kGYrHSkVcBW/oqh21oE8Dx+Vh4VzOZtaHjf7QLXKJ0U7UrNPy3ZImdI9Ydhuy8S8QFms4td5
Un8I6e4pAsslS4VBFAdzVySAz1lmhjBBnLBugGq68/Ng6cSkOZFHKAySIOQlZHjNuVpXMbNMvzQH
sMV3AcTum4Zkor685+zThh08CldFgqleH1cDquOy/8r4aJCr7D5L1KSyaN8Xe+9KWF6ien0oBx+l
pKjONEFuVRKQZAMARkhi4JJ6YfT8q1L6XgXdsxR6ZqgLFKjqgAfWDyL5f/xYS53JZCvK++9sNpGD
Y+RRs69JcEFmyNK/3A8FmNWQwzFFz7Hz7WXpFutaFMmrnMuC4nxkAYGuG3sVc0IeviQuAPLAsp3R
XSIqOOkALaCUyhOOzFXOU12AGI3NnovFGROtIHowXj0psCMWbXVenM85pRwBeZ9p1DIkEH+Hfdm0
Kpjb0+8o0AFv2S+70TOb9PXW3I7yN8pSI4XWCOi7nTY66R1rJi8gMrZ0tVYb5rCJrGMRUe5ZkEW8
kSieuGOclFXAV++noUloBlOOw7b17WZPuQmyLe7qwowzx9xHspCUTvCNRkgARiP+FT2c2p8I1bgx
e0uIo7senUOTs6DnOMgfGJcRzbzwF9wsJ1luE7il/Q2y8/6+Mdgn9NB5iRPzrIeUpUmh1MNnrBp9
+YN7nGLfw2W7ocLZp7MPRIY+qKuAe+YxTJbp2oo7QjvTTxQ4+PoNS165lU03XI1LU+xEmuzf8Gb9
qNcChhLC4TqwDzxx1qeLfsesdqdmOQe5BsBFJE0yrWI7c/BzCqzICaP3ZFUQezRRf2Db3b3kdonD
0gY2uYMQXzKYueA7kGoegeI+NjyY+RjLpJVFWyoH0RDZyA5Ha8Tuuzy5MILWoSI4ihVvVLh6+t/K
1ArMBWhGtNLH9EVp6rPKaqO1MTjoiwqQa+YBP5BiBAXIAI+skEZGB9obE8HjmhcKzI/rQeKaskIh
MQQppRcKOuwv26k1H3nmF9CnHq1aGdHPwJADxrjfObiwF1z86x1MdDtYkulQxWZdIRkYeBeTbJ4S
Dve4POtDbz9ea7ETklPLwnL1CKCOZj4WoaT426mZ+aqzSzu2pUPBlDPNAxV4nrF7ku6jm5MXVQWu
uIYmAmzem3bUjNmBg4SzXu/pHiUa+BxMDTY8B+um5YbCC2oOr+DoKJHbWfijjhri0wJXEh6wQiEw
1EX1sUMVFtk4nv3m+lOX5EVAYtIezIExzg1osio+e5FV7m1M1C/hLOzJC+fQKrnT6KZFEkNHEktq
lCmvdC+cDMPvDZrlmL+o+OhijcyUhFN1B+cc8WJRw8sGnknTWcCmu7bG9ku01bMvngoJ/Mxd4yJz
pNJvyFPhzuCcVVs3H5dFvPYoWKm1blgF+M62Rax5aoAFV48ASHsV0MEV7zr1hIyZ/CCJoByH2e1k
k74ThYvk30by2ZcGLM93aEDHFmt/0vzhDsZcYbTrZhqPaG441AjnS+PQkPuXAblH3ETB77llaRE5
8bdhtE0e3Ro/ois4w5Emov3LolvZLF0An+JJSKqOisGsQ5p6CvBpJjQp74romal7wkJI5cZSjOhW
yVdafT/gUg4839oz3onOmyBgR+TwqZIp3AAAy7LSOI4wMGUwER6C7Q4h87KoKtMRzXGdBTUN8BcE
5+sCrP3obov+aZDD7m9EFCsf1rqAw9lWAZSS5X+967eNG/TdQHrLoB3PKmahnz0sAuu8U0Gle8Rg
5ERFM6efusgDzoJkBqGKulvKM39lX9z+s5AXKwqF33p6PXz2HLvHnErq3t2rtGKZDNF13FkhnduP
DzM8QUNJF5CTzAqPaXfTloyimnrtIXhW2tkYs1w1b95YdN7bcnwVR0+ask/tM4Rz8flY5ElrUBYY
gNfSj6nshkpUppGkNkhrhoFATKC27V79sJ5haULA9xQDQ3PBF20PMUu7NFhQ6EWcLVL+BVVetMQR
nxiqmKT9nGtRrvY8shfX/oY8bOUGf6yk4uYwgk1q7G6jjYBSN+G+A4J8DbolVEw71VjVtL1CRjeU
AMLf8ncrqk+6Oa21dmu3TzwVSMuo9XaE8YbROwHEwQQjLhHmPQMWFokzib1Omc7/ImNnROmFWLIz
eTV3cjaoA6DAw4Kwv3C/OCCbsu+Aa48eXDxdiv1plXKynFz2bpllbRphZATBuYFGlNlQ92fL/h4Z
ttay09SzI71OlclMQvwRUF9D+Kp3oEDnKIHT9d41TLQRn9at1nEU+RLNV+GVvW/DWQJT7ao6olHI
drn5x68RJRvZRfIFUVtyYruoK/HCTtfhwcicifu7mNFJsL6l3Dja+4pjTnENduny6N31b/VfPmPy
OFMfRDNFGB6Sek+pNGtBLky/i0vgonSLNE87t/NeipunA4iIfK8PqHGIrAJNZccO4lIzXtt+bvhR
JGMlxJSyrK7tpr+R9iif2wi34NQq0+QO9wvzLvD+vzdEIdkYc+dqvqqsXonfpf8V98OfQuNQJeaG
aWLba58B0Fsu1xZthwBxwCIXontLNANEQzI+Q3gPyVWgwHiv4rrTgyYTrKP6PIAojyOLVaxliVMY
n9mk/vBUeFyQXqCI2qoJzKWiYmFB9Pdv+TkBR9c+3BASbuLM0VJwC/mN7ONugOtI2hxTzZwfT17D
gqdOaJOzaOwnp8nKpGJC5v5Ft8cvCbavEZuT6Vr4eQEXfrp8P3snTwEK0eovnbqSV0j/Tu+AGZcy
8FFd0wp4vNQ3Qp5zVgrSunvDrhmIJNmsYFGwpVuMkYmnt3X4CYGBNOWzZfTs0r+bIdCbT1oqnmH1
+H1Gr3HiFSwrA81t7qluKmYma1Yeqg6wB+T7Jm1lrc+BF8dZ7PR6YI2kpBuZrBkIcmCSRw+Z+ujA
/XOM4I7Sa/MP6M7IUB8dgScbJfMHrTgRDCdGE88GTFy2iAbEcrahrCv1JW2nYpvfKrM6N2zcsfWa
9zq8U9ifKvbnWaQySK/e520iZb/DzoWE2y24i/DHKWoDFas2OJf9SQvZcgfA8Ffccsdk2XbbluEq
FK9r9kF2MkuacoRX1RvBJ4/C3Q6Zg93dmwXi3PoWxZh75Cb+RxgBYmcywVtJLvswqZJQGObXUKEd
kR/ip3690UvOTPDpsHsNkDvSKMkoDLdT21pzaXnhNH6FZX8ZYOYTp9PqrNiEuihpFdmXPkyxFlmk
NDH69c1OkE0Nd+HbCr/030DvCz18PkIaXupUKJ++0NaSvltxgU40jPxUp66R0M7oP1tpbNcPCM3M
8466SNTJkEwkmrxYRxm4capRpk+N3scrBYetYh0WB6FaDyOcS/Y7hcAcrVTxqHiF73ce1n4P2U5z
Th3uq/nZb4+/7NrUz6SFx3FpvDbUrkdZsIkddAh1J52tO5KWd+nZfYYa0MdBHInODq7Q7Z7faBnv
mOvt08VJFzgmHko95FmVDzV399Kf9XWMUPTCpd9HIoBD1db7A+8kEtbB/pfBIdwbosQsHZnCYKq/
+YBYosPyLfcXsArMwUviXJ45oJI6QCqpEDyGQaKPm28rlVkgvjDRr39oZ0QOz/ja8Ehb1gb10mRd
u0k/+a81eJun7SCPN87GkWcwrrWJcWE15omQ6/MyfSSaWUW4xVsiFc3JNgCjFNinASNUqaz1fRXp
l2y7kYIAXzsUtz0cfxye7oBbbMcP5nq2cWrTKb+nMSVzSpDCWQul9vdm8N8ptfJiYnF5kRn01uq1
PxlxRYD2s14bBpSwjbUURSPHRovlqhdBXhbdm/MeyAjg8tb8mIgxB0BmvCB12B6mcNXoJYEzHOcQ
IuCrYeIQPewDuJk+y2jadWdJGwZRUXws27wdAp2oKh5tN8XdfpCWYFk4auaDwILrMkhpGZIx/L4J
MppRoIs9Y1Sgdu9k3kq9ixat4OT3rWkjD6PVrCJE2nlNoKTPIZ59xpeRbOC+D48q5OrfDlolePTq
T5wFh+0dgCqdNghUojzy4LCCbuX8vljge+YVoH4TFHKTMBPTvMOXt2mWiN2t15jP3kpepNI7yn96
MC98qtQNuOgqJN0OHmL8FwdiH+6BZqqvhuKeOHN456c9XV+k3LdsKMCHazi23X6xp2eO2Pj3bReD
zaT4c9g+NLuPgMXqPkdghUJqqlBI143YFUraLQKeX/FbLnydbg0hFSopMQf8J+2HcPPaZZAQ9We5
x+Fq9QYDRni1h0nUFZhtf8cY2R1mT3Wjab5mWQHwQslLzN6OXFzV1loCgpIrwwME0ftpRMAOQKp3
Kd5EJBDJpMmy87/Hhl/34jOmbF0EnLSWLX7kQ4o3ZfGZ5WB5OR3gXq9BX77X3O/+GQs3X7upChQH
LJwz0PBt1EXYzhxdY9nXIVHpKm9jETMGuvFYHlzRDgDyjNQsf1b8KV9sngAkeI0OmvtKWEi4wAXc
vjmwx9XfQcxnO5+1JTQBsKZ5F4VAaPY9SbDEHgKAbwcGfevw98EVsd1/JU0TV8bG20DmvIR4C6W5
ciiqLgFp9EvHzBBzWs1E1gzDfTebyUZUqc6HASBsxJlTXF3NVMJr6wRDFud4xQ14+lm/UXeFQmCM
zEZXIjlq/xg3rQnFP2mu2KqqxvIB3Jx7T5I/TTPvT8VW5vLDYU5ZfMDBLgbLyJ02hzCFetFUKZ3Z
D7K8pkQFWpQMc0N80/Fk76yKrbVTKoCm8P7Lo8oXaTo29hLilYT9FwWOxiNXmMUwAl846fIQhQRS
xQfZYXDstdh9CSaykAaU+Mb4u7tyQPMMpxqykihvbFx3tzJO45MQms9INE1jVbfvW7JPg+niEPua
nROTcfbQrsL9MyMLDFp8yK4nBzGuG0Qm3zHpXQnywtm7OR7KIQLf6hTYBsS2FXizVvtUbnPTkjqt
tzStfL3DhIwn/+wLtPVYOVU1vTBKC4jYSWCGtwuWgapQLrIvZDukmyzNxUY38QfWbe06r4VcnzG1
91Oj9Qrvl00rgFuoljPeVI7tMGGf8Sfhmi+wAx3KdGvIlbxmTu2Cx33koHVr4b4jbV3/1gu4yluh
5dUVMdY/NoizjrnIG6g9ewdkbUjpXYRLmhpN0F1KLY+q7lgcP/TwzOyipTG6H9PsW2VK7UeTyRmM
W+gVDmK/pMBm7z7vVCVKKA2nbLh/QOjjkCGMHII/08JgPu+MW9w+CO8bK7fTvg59D3xX93+sgriW
2u1M4/dS/A5z97NAFnXaRhOPErlxwT07PspRKJj4EJ4f3y65cQKt4qAyGEJzZWAMwyNmZWexve7B
vGxbLF5SvH5v/Wbn8pfWZ78fl3v5exyQ7esDdKMvwIicPxdLwiuZNcKyMQJMc/tJY67/yfzL7hRX
Vmz5R1X9UVTbi63aGAgr0gz8StKaT8Ag6u3Lh4CjoAXJ2Xdt7HhMD179Nk9+VzgzgYiGcxYKGCnd
hRgIsFxRrQ1p8j8GL2LL9ime67kybWdpD1N0H6pk8W0sfwjjJuFpCQc7utEi25qMlSM7RBKYNgso
5Kyf+ytoxAms0ASKp95socaqzjKVYUBAXu/Pu6flA6qdtdUZ4j1a7XqaYWnv26R0f3lB+ZaLgEFz
jEzqgdKQau34hAo/geN0X0/rywLBoLJ4RPI4sHety9oswvR6umcAb5XSxGaPufvqtyLB1z3K1oYY
S6HALKfZrtxxvcesr4m7RMzAE42oaVq1gh3bWvsH7fu/1tYVljgQ+6NuUdSxeBSgzTKM6k1MqNTi
02AQtDNpqf0twG+MGWdhmCGk79daLIFXlyyGukOVlUTYllsaxFDbYQDByBBkDXepDZdvbx0f6wYt
Fd3RZ6WPAZx6yqR+x5sm/4D1prJr0GJmD0XWVU/jiJhEf3pKxNeTjifuX7XPCLcV6OHeeM/TnoWm
3JMmHg8cJTuafsXHwjVSuAu2m7m1CgNz0LZj8RKt+e0xo9UuuJZbZ9jiTWRx9r/9EcTeQE2dwsOp
ZuCSX9sbkKq2y+dHe2+ZD6atU+8zj0mWnSyPLyfFBcJT4mtSqZoW0MNjQSFu6OhY3vN2+3vR9ncy
K4cMKfhqILJRs+oV8/hOHqHXzEWRyoyrm97uVa8rnGJbyzVZWTXSO5/s+sH9cVwfi6HpjkI5uPvM
1xGraFilVEGz6HFC/2CEe+5uRzdArp1c7YZ8cEksTlwdo9Ybk2NSlS+weL5itL6m8QQijPqrsMKa
7HjLBMYtrZyLROCL+5Aqtw0us8X7tu3FzhDaL2KgIvEU7EjC7K3e8Esajr6TDi2lb8/XuGIDiVtn
vcadeZebTGK/ZgoQfI+IvbnnMYj34mBEiP4eFSyavV2TAD3kLHzjo4Dy78btpFelYY2zgoBd95Nw
XXbECXFzgORiC6hT3ikskXl8hWD008lCLdcIOk5zfW2eQSGwU/awOOM/HHCTzTkVVmNXeZ3phSiP
U9w+MmOVEbW2k0klrKqUDAKrJOr0rUJeTmo0DJBxFKXTZIUYYX/mDoHZldaLLpur4pY2r6/t7kh/
wqW6oVVwo108xTawFts0XE2FvtgcuIiBu4rbyvQYuNzUdwNzeJLPNa9DmMu6Gvg0f6SJg5ukSxaw
+eLD4wjnWlSs2nC9/wC2mdOyKvuviud2/YxWZr0jqL3Ej18L24UKVIktM3mIJB/cyOUqYofQnp0h
Yvu7gW4/EtNsB7CAbjbeOK2HNCJgIWSJaCfTS5I4bIAoMcfSlCwCxPUw23VRrD5bMcpEOuJpVy1Z
VS8zKrZmY37BU3ibjynAGMTME/LJ2OQ4E4YI9uLda/sXWjfSS8CrQQVOsTAKiu3qRGrpkVgh8lER
SFtnkvruOMb1KdpGbxbG6fUK3OTwiRl6DjzMc8vU7QvMtDNjfAK4uvm3lMzBPqPmv2ZLf9MFZLP0
+kfdgD091PfY7qn32J1rKSphd/zMD6Pd/mxJ8g21dIk8kiRmK9iCiibvrIR4MPcKGlZdKDWTGdbq
JNLhiAUvhQEmkZUKyOoUUwNYJIBH0S6uUEnwmht2S+6rmrbUSic8LGza+GuL8jb1MW2FTlgfIGiJ
35sa5Ac3oXKGf/Nh44a/shSSWlaimcVOJtgkTtZWl2/GyxooVuNyK11IrM+Rl00HVCVF20QWuJQh
WW0WrbozMNvTX5fcRMUlJyoJls+C7zkjKl9dBYFSuR6goJQVBRWPvyydFTZl+bxxVK5PsY0V3Mqo
byv3u1c2/unRK1l9nSkEKshUAztjpgZ8q+jSfKW34obwO0x6Bo/CfhDQBUxVneQ0Pd2Y3BzRjpNC
+UwY9eOQRzxMFwWslPoXLh0DyvOeI4dtvQ8d1/it7NDfBFNUUuS/hxx4Bd9iDnoV98SHDwXk/KSm
vaI3/EWmlN4I5hoT+N9d4bOcj/ZQ36tGobGf9z6dRJKeUbr1DkiNc0DnBAECsZRz1MhzlI5cZ1xI
+mft/hqvu4mtz9IDoJ/LYYJ3JZTm6F8JJppIYOMkBHcN0XDbzP8y7FxXAPpZBe6oTu0+6viD4fjx
yVB3zFcGFzhoNPWT7N/5YDJQjMBR+lYdWE2Ikl0bconMA7JruCpFxgQLIF5k4gPQwsgcy9FnUKCi
0InPLLhWHMfqFOZ4xks6x4f28sXSwUwTZ/u06WcWl7rjAlXWZg5yzx141aiWMdsbcTfHWFsUZ+ri
6Eu6pw3SWiGU1WyV7LSoiLElmHk8Kua+O0+SENAw0OAGPKD6SJXjRcwWWyCLJn3eG0NGjukB5MjS
GqVFLLm0vzq6t+m+Q3JRm9zRoZ6qPPIVk4F/BBK9PWRBZUkUQNXMEtXkPWtXTyl1CWI4aWJqfb1D
0rR5DFGBZo/XHH/AxJ7WCYS+tNAWvWCMWyDSbLVXVkc67yCm4p8AtXXC6nypvzROzxcYLUx+XD17
yGbjPR2aYgWm2Mm4CI2sWyQX57FYdzeOvSULbgTLhHUMAgjSAKTeHeSkeEuf93weSvn4JIJYspRY
Ted5u1cFVvDNRwqlj1QGnd81zyigsRLrsaKddcbWe7I/bprM0Iw5ugny/iLaNIe2m0juR+WGc24e
N2xtIQ/hlguP+GKSzq/GxjA19Aod6VdRZJCKGPZZFshLT2i+KlmpgAB+C2cg1xdAn8YT59R5sJ0+
mXN+FuayXLWPfRBGpV7r080MaLpgg02eVmJo8SF9W6Vs3ITlwlM1DiLtPRP3PShMFLGpzFqrIVFE
nWrTgLWLiuQ5LB6F/SUpwmzOCl/y2/3spRrDw4jG+axHmIGzlO4jc/9KNaZyv8YOH6mgOQLdrkMP
7csAHtwBDPpEBm2wJCc5wbIMtXA8BytiZxg5Dhf9czFYOtdyhYw1jiY4FvTq+ib3GluUm7qgzzrc
6lklWvXrh6YAbmYYAHLXrx/atGppexrDnrEhVbNYqz4j6yYdH8BdhwaHU6riA6Gz1kkMrtpzNnHI
NOLE9g62thCWP4vILEqzqYFOAeReP8f6SyQIZJ0KfnJcImjTukHOu2kF8VNAkU8ZDOzb90rx5eC+
oq7AuE9ERQF/upAgWPKGLTHDXSHVCxWf2Cd4O2KGO4uGjUn6Z8/YYZjPiySXGD/9EwbX+RwKvEMk
YfoIq3WRFi+vIoThtJ/TworopNOSz5MZPBy+otUH5oWVbWKOh5m3zWuo2FUor+VvCmtjI9NprUnM
gN4FBffRlJBzCgM1cKwWKEVyaKKiewbM6aaaMy9mSRqjLaZYmW+OF5CX/e5fTCiz+zgsEcYl7p5j
gSLH4wK8S60hraIM1vols907X9RJjJah9QamvWl9bB26Kgz16Pptb+loRo/dOZvjHtlXMuke55Hn
ZnvKekd2mRjjzL1g6GyjCtBUO8DS0YLOg3DK3ZVfuhHhp9d36AZagGx6WWizSsrE7wUtoy50ULQA
Gie0tu2q2uWrFVtZuO2TewCXm/sc1gUEuSElTTuMCtzLIrFTEXblt9+WZiNedYsrJkiLfMl5ahgV
Og+Zh86weS7DeCbmAIi0weCVMS1yeE3iaOIAcM+V+Uomfawmx/YbPCWzh4ksgpKaNzbfSIHqcpz3
gxf/afIJ0lEx1eCGNe5KYBHcyFFPe99uarW+0/o7lKTy2a+XcdBe/JlzSgm720b+EGgQGEP3fyGC
YllsY1hJtisHs0oc5psrY9VjBcQ8anRvMK7yrFXmyiv/xim4WgGHsK3yP3yWwrMifcSgvWI+bsbt
TiwrsDQT9giqChTCrEdy9JmB+EG3THB9htmMgmICIPWSG5E+1eg1DADOffH8dlYCnxPrh0TkNjov
TZIbl9RBQ+i3VXhF/cBwwAwQVAaIn1inIdJU6LIGIiGPSWYGutleHyDoE1dPJF9JVZnoahw84Oo6
6dRGZmEh8JrQpss9yn3LOOxc2/wbHU1RcTaB48uI+sndIBTzHkal6wlQiIQJ2NASnwCOe1FXTre6
zD+iAuOSJR6FX0HwD4GzGdey1n9mXuSVR1MLDPZk0TRw7/SAPV3beGsfcNxvq5c7eUUx7gbmznXl
UejhDh1DQUMoIAJziwldvqr9hSijyGd9XwOQ0TfqXi3CW1zXIvAjuOV+pdMb8fidgXv86cgvuHML
WnEd8c6F4APvjQHoqCMLu6Pg4mBssA+X7PxQwQsv9GYi0gHJo60FdejUZve46ifE7PABlbyOPqZm
j8BclSw+PvHeHHqjxOJQu5C4eqKBKKomj9F+o+j1T38DyLUtUVXzPccFV1Hn/NoXFrYFic2MD08u
iCrHFXPnWpLpZVNi1Co/6xpLYANwsb3gGvHrxy+mboKhG0r8HaUOpH7+SK9YD+lvWdE06veN9M8w
ukbObZKXI8dP3naaqKy4dpiyizkukz+fn0aAWw8lbTD1XGWaEeFNr4nPoFLDyWkB7nCfK48Ydwy0
aHdkyrtj7YtqR5sNPn9/C29TnLiDlhXlzF7Bi7PxKUSYNa6ybcgyVxyTHeRnpObEGbNhCel0x7mY
qUcRtndWfkg/HnBpZYS2VJ7UrjOXkpW/lmL8r5W0WrXb2uzDt6jEBhoC64dzAzGD7VHFlrv2oHIU
5ElVhMAJ2ew1OEzCZUYNLXgFBD09gZlJUhARTnzR+3mRs1p/z6Dt0T8u5WoRAkqhD2w+nnnfDSf+
kGq5uKPaLbM9F9dfLv+y4tcOTIuzs1Egz0hxJADwFAJ6D373jAntqaiG47G+CJpxTt8oKnvNrVpW
s8WXEH9Zn7rFRq2iPC9zTk4fdO7KTGRGXz/yi2imTsCWnLfQwU4Dz9HxqXNq0r+8SSEfRjfrEYgQ
SdD+dxM43JSGQnV/GSC35wq5bGmeEHIPRSx+tbv0mZI/lCsJxqkzRAppYWAfmurNe3V5eHdT8gNl
vvwqqIS1FsVPLnVdWdjpX92DdFQQd2rKMd+kvKNmS0tOs99FPkWOJpZxUWxrGmpfuIULNz3v/EfM
CNxT286oTZNUZm1cALko2voihr3GWgPSpdkbXQfrDWoAKk/oW+a7QFx5W8hEQdmO03HyPKsIDvvE
IeE5/7OXTNVXGAhQM3loldctthk13AT/VduFpyw/yThXdLCJeSPo3kCqppajSkN/1QuARMeW89jx
oaAqNMJOiNzZ0MUculQ681uxmnO0m6x2YqOZ2wPTQZFo7J4m9SrKJWhAKlCEpN5CNgAxSu5O9BzZ
T7PnfowAmvjYu1bulObejFIykd/peapnrjfZTcY8XD6lBEvxRxYlUpX5U7wOibgGOcvUDxGy01ye
B0oZQEMRhILcCCwN3dnf44Ggx2ns2iCMZpQo6Mr9WWVvgeQuKQceIkqqCtBk+5IAUQK2QfREZ/ff
yMqRX6H8xmYIS31hsHgIsrMECrNrBaI7UiXyHeQQ+YJXrAo92LEYDkJzplzQCV2TUbtqD5nMOoi7
rD1tf4/M8uFNLz2wrnT0142IERMMbgGmOmGbQ9n/dYf1xsD1xnLcS4n9ocuBEVV701Erq6PTAPQT
KGKf1Wgz4NPTo557JSQztig6d5A4iBEHBKJf7qA0ZP56RDOdFmLO+pX2B+w/iSIDUyGDMTZN7d7L
QO4yOIioWRXa1pGiRHEcvhVWUbh00asZMCxj+bDohz+hpZtE981/VerbCMSdWj9YBvptabNQaSJq
BsB9OLRT/4BpDkT+DtU5k0Y30Q7hVh0n82QXlwPxmgu4rNmdwtOxy8QAAqki6XWl+MrvVGANMk+M
rlVsugB7QVLxsYN00Vchn8ftbtKDj3jQqlH5AkzuNKT9QlIWNxFJ0FUiefmI6OCFPyaT0o/JzTd8
tOnuiOUs1umXSnuQZUborjMcuc6toK2OLuTlaPm3asMnR4xke+kwrf6bnybkUynhUTdjitfeNNmW
UCtk1hUc4ZYWZwCy7VYztcbZmzZZG95XJqyXhbMkhkII6AQmolitKUMYLHPVw8ftd1G6dnHN0kyV
YDJTL2DZ2ps7P5MQ8MUQJQC4piwACW7lIfr+LiTLTRUIP0ntXjkH9OM7ufVVd/nckKRzk97a+24+
A+wAVKFiQtfzvul0/wuMKoyjw8rqGGj4g7b5D5qMxvRJDnt0RWZRvc6vfA9EH4Jvr+rxG4wiZYAz
ZoxEo4jbhVXbqqfBSNW5IAmmqfLvXY/295shfqE2zMG6yKlXHgPGjq3GxRgwA9AJNs03rM3/2Uab
eGcRSc0FF7tFqdnQ21J1qURW/ZUUSp0aWf+PfzrkpaOkerd5wg9Xx9oiRCSpl6GpmeHAsTIHAp5Z
q31VDZr+ZPdPmnP8Blo4PXoSxmBUY99HLUmkAfNDkmx8hBJoy+ivgtOJb4PhYkAbKWnL3zZR5Nmf
ULWF7DT5INf+5OScbP7WIJteUM0L4oTOhKjhFNY7yaVsnMYFSOt+ApRFAgLqE8IroRHnLnlcQZDI
9KCHIOckr6mo7J3/JxMMh8GjYUw/uczlRmti3Nn28wp14QCOQw3sTazzr4skUPphbnXgrbF+wiWJ
ZpvG/lywi2A9WOV2316fCqI1CZ97ZH2liRF9XSL4GOy79qGic8OogFlSXIQiCFydA+T2lXTyuIwo
rWKYi4UbCRvy2HTYRzT/YbRay8jZENuDahSbKxI25rjFx/XMn4ATdeHncJ0LFoMe1wFxafwS9SF6
FCM2OFVjly/W4k2+Ocl42+tvtNZ0ree7PhG1We39x3i+qkNmyJIZSXjGxrDJzLrQrZp96rL4oS31
g4qrR1k40W1xqnKak0pidoKVnrSRVMWRbus41AWL+71XQGlgDy/q63DK5Qf9x2xqmMfIRRfPRokw
wQ7TGLa+kYlLBk+Xnwt8htWXhxSgC2Ia7mX4Lo1u9fmQPLft6r5QbKfximiYxZ+dGfYGo/fF5gvC
zXKY+bN2FgbIIa9VppCX3XhpMWL2k8RIILMUDbQCHcgMrCK5539ITog90TIyv93CvBKTyCzSgI1k
lIvMHx1uHlLCMY0mrNVqKJrYQeF80h0JwMvC7xfBQa5vYPfdMoBeH2kvZtb+snjuKIiIIVT4Ruru
ZAiOECHOBOO8ugM8r5e3ahfzrGwSYdqYKXSRxrIgKyYqZ/usj6LALC04SzSPKTkCeRMcDihlNZ2Y
Fv9+3ZEPtwdj7EFnF3QQXj9mllCwhNMEZMSkc6G6nRtid4Toj5Vf4SkuC8FmKeJnFaQNpZhVvOxf
KjN7UYcaeMhdRYSc4cvY5WIQ5M7MoqIo0FN7RYGpunPX+nY8p1lQEkVIHM3K+JgxqzNLC1nXRI8p
+pKAAVQGUEN5KUsHhmeu7LuLUAMC6oR2aLFbWSuHKqAR8qEPky1hTDtFOm3cOVuuY2SaINI5q4uH
AQgrElUblFnFQYT6pj4Q5Sc6dHPnPwWk6mMxrg4ATmoC20MrnhojWl9N01rDJgY75wWmyDMd+Y0d
QUP0TUYWGP3ysdwQDB6cY1rV6kfr9629VYID4LiTxIoaMA+VmlzTJFG9d/1W1gwN5BvdubnkuvU1
dsUNwvxyMinZwUkaGmcv5lskBZ4bYFHerpkiNuJT4olt2OrC22omp8a2PFmRqPR0QxJA+wbmZ3Uy
Yxgr0I3KjUH7zmoy0szhAw2CUR8Z6DVppNGFNj96O1fLFLjeKUNeECOXYV2Sfyp7tW3rN9YN7wej
1aQHkF8g4s1MCDVrpV+ZO4i+ulixhltZ5jWa4+OCochbqxLa9M9jI75tdpFbA+vGwiDbphyhpsvZ
VRi3YVeInz0JjwzTxcFDOnoaiaIUNtgENXSfkB3cEr3lt6jPpeTidy3o1OiCO1SbMfoE82ZHlT+0
tcl/zY1Ezosn3JCz9Mp2FroMzeA06304ui1gWuy1mNmF8mXCn9mnLj1YFuTKfbjYWls6U+yGzF68
iKVxjoFe48mns3uNb4YD3Okicw59ObT2/HU4XIQ37UaAeTYI2zib5UoZocjqR8cqFcIN57hDZvsr
eFvVVFN7t0DTLWclqkB1+Ju3Kb0DETmShzP0zbLI+n91aM95CEB7Q6NODm/QGooB1hyK87WPBm3/
gky9OU+BG9dV1oeGIvoJqdlZSLcb+PME47f/ts8xNzdkMEHEPSwTe4omZxls+uiuJYc4rcAVvyoF
28nWYQ5SkPoQWOsZxs/I+qIJl9eE0qbjHViEBOVeXP15VRfN9YMG9MPmh8+MAouxqaqwCz4sTtJN
XYygr9GGlYYQWZaCAgoWEgNQ4oxbY5HDdKkTUBPvRVHXkN0oGzFf2A+u+5TcfP4XoCoMbN4T2eo1
EjYaHNEnaGOI802/WxiDPfRPBzbHkcj+7TWv6bO00oXJqxdPlxWNuU/AOMAaXnRGleist0XimCQs
FuKGOzdZjMkBQjAlXAjHiNpeml4W7EBEa1YZdWcqYhFQeUaeO2HcR4u5zolhtuvce9aU6tmcXbMF
b6BC/Zsyyu0EXe9YmCNllslRHYSDZkEs8hYZVpFE7Tcs+FKN0UlsWDQPmD9Z28SWrD6xxilaXk3X
eX2ruFAsI/b0HAHyeyFOs5LKhF034IZ38Gxd15+T68ZceAgPjAbNK7IC+k8MejC/Lhpmwy4xvVgD
rurp5E/faTnnSxILfSymfLv3m/gi3noq8MPVslks/yYojLbodpTEBEedT6sRv+zTvE3dt8MCptCo
KTv+3JM8j/E0PsxnrT3Mn5+CyE7HUyAR0iNnEVDByn0uTKt7rjyVZDXe0Rfok3IBZCZYx785uhqO
tm6a74CHZJnl3T17BP/uuwJHExAZMp/Q5b/s9Fjp6I9ji4zjc0WZnxze/3Xob8l8D/PPE38JsF4A
T87IuLE1sLBdb19fMPAjCLUJ1TlZxZQKbjAlL5BgXl7G7UyENfRFqO7/hCdNZYV7gx/2AhLiPLkO
QzvMBM8orCH4iQoza0hE4D3EN4BzxX3pfOwdW2ZD3MIp1OA8kKunls+JVDtL8TPQhwEV0eWTAAE3
psHDlgxl/ytqfLhvOUnNmnJaMEDgIfkHOIvfOx/a6kxRgMWbnvYxHMH0XHtwD75lo5VLtLjoIUL/
AjsOmoV6yLXvBrA9tBqbkkhuzanJTF5uM/aq3cEViWscQuETQ5fv+eI6FkgFAt0165doLCAHYtPV
ud13gjgp+j2ILLc1vquPvBGCFvGFPyg060SCAVFDDLeKLOosYHOCDO2683zJDfrFok0VC7hQjgWO
OnLqpCBqIQJQ1QBzA22oVKWBHY/VTRdh8YpqbJgFt9ReKndZGCodTgYZMT3KJuE+HEt2BxazBWGa
RaxocpiS/hSAqL2QxNkAcTHrq/yHClJiAZ0Y/8fjWUz7I5+UcBr73O0brKjw9zKGLfkGFnulVOGW
mIwlLG87WxmzMnNELD/7cP6ayiXTKA9WzJfgSquVAbaCCzbA0KJXLGQfoI8LCfsLMm938VajkZYm
fmXfvhJct0hEge7D4aZPAu5jqDCHgg6DDDMgz2Byr1oJoAtMhV3eY9Eh6RAAYuDg2v9neoIoYPGS
m7heWLT1ptg5c7TVfywzP4pe7R3niUturNypykOUicaRUbFZuwuCGvMnKMngo+UqsibQeb1Bm63g
mId7nYfHMq6jX1XkfF0x5V4xPrv3GwesIdGxAdfIE/98MlVNaz+YR4A/pHgArFNWp45p9ygpYFRt
mweYtpW+Ooqz2uFu7kU55ky2SjGsPSRobeAxlIvmDcEMXo3BYvXCBd2X02WRG1LTRsfFjDBjW9pH
u46CXHO8Q+ukgXYzLfSbuP6Yp1qQjTga8zQgx8Yo1XCnrRoU/RKgnRMXlsvUj0Md/4w0e42Wz3CU
XuPXGZ8Joqhi60y7q00S4POpqjrnITmdVNXdaOQI+yXSWfJEcGDCVIJs5XUtLbWYEUhEG+vnPIUc
7fm1r886FmaVIIdcP84xLqr/gex/PL5rYWkLIaBz8iGs/Y9KhLSLdaMTepLWP3PnEu+0CULtNA96
S7G4xZBGzbU02PzL0Dsh75GqOGobMxrpacZ+swscNxeYR695xiLqpd1DDbJ2lB4UXt7fV5n4Rry1
j31IdaHCe86vz+5kXxCAwqixsZcgdNy0qeeibRY+nUDAexmubR3Z2LFav/cLo/MwLqx4ZTEpBSjp
V7FzBQ8BuG7+gYNPXzisqJwL03pyVgVkEErHurquJbcIqPUjAVpb2dmKOXolShK38baiVRIaRbQ6
PHj5BZG58dYKUfD62hZVEX5rdM7eEYHA+bh82WzGXIZSGM1kAuXFEAVoYvPuyttJQQpYzEntX2OZ
a1dmisPy9Q1P9WZ5HOcX9CPtqJmTJ09MUgLo1vi088CqWd74L4J0wNmetoBKYsA2gpAMZkGTXlkW
u+FS/XBaqsX6Qrrv4qU3zlJy+6PfdOSguv/QwsHdI0bMNV9pXAepFV3ysJPmUnnMdz5QJM4O4k9/
/FcHNWRuLvotOcClMG/nW7Q2ZJZMhLQSiROiCUuniDHVwSfVMiPsBSxoufRUGn7tOyeOhkTa2VvS
C8iZ8OlTIgv3QDsBJsRLG6t+jtqZXgHVbHXVh/SeBoJeLGxtnlW+bGEmLMel3doobFSGccazUsSf
uEL+ONOgRhq+xWVu7VmrDCMEplyQNdVfTPxv/Fw7OqxJ5wchGfq4Pm1Gxb+GEtzwigqWo5MmFFha
k5rhIDfvD7rGo/BOYGe2WK36oMRXjKPanxeT5rpnAieESVxNU9QNSzyg0JUaWXQ6w8dqfnhLtldP
38jcAwHmRAhdfZutfjPlCtYrxNbzCpOAWJsJaWPgTtytPP9GJ+EeEhe2F77u0jO5fOnJsV31b2Fs
l1PUwQTq5g639arDg3IMaA4tflUHBmr3oSKbdc9fl8KWf5wfNNZo3iGMyHFWU3oiy0FqA86w64EY
oopzUMPsKZuWT2o6T/oqx4NDpYdnEF/1+XkUdPybT2DUgo+Cmkj4+AEjvQG3JovdPtxB8dd8Q3zg
JaLTQvVJIINUbpjtHIQs8JE/dx0lopA2fBH0ODT4kbQbgG14VYpa5DeZlzZGV8qy345ZQnNfJAKf
EJpbjNR48uxREaZJVbjRfEyT+H+vMq8K8Cv1JsF8M/BDY6U2wrn8P9k+pH4YsJ4v0llgc9UUNqV8
EybfSx3drVpUDEeIO4GkzOnlcs5wweJqBjMdXUcZUkm1JeudcUanCPdQdqq2rQOYrvUC15A4ePeI
qm6h+eIY0ZO32PKw1ZJ0P0+kTvKE4890iBz4NhoY6TI5OV/NAzh3c4iKEVjHGHwK2RYRF2VlHwaZ
OyMuDKi0ViRSXx/PxXgqBgAIInOqvOYNCVppLSmGwXd+KwerSpY/4wZKabhVjv9M/nfb/OPLlovV
nZd6cAaBPFGAF3JxZNqFBY+9UoGmZKCCOYobMw5hjw9pe8yllyDsjCqxoIOblW3NnJ42DpkEEyGs
7/qDG85IDl0kev3CtpvWnv6Ub1iAF6zH0IkAEl5LstXvgp8wKUw4PgAPq0wfAaZhaR4ioA59bgAI
4CwU5g7bLpcV75mIljkRDkLGQ844B0vPfrfLxowKwEtf0asebbeI+uIsxt+5QTwF74nDdqWMyK83
1LL2cSbUDy9TIZEPxex5XtUs/jc+qGeu/NEqBmt+hnIg5kfBBKDnTJ39kTmGJboUDY7z5jknbalq
jX1NiegyAsqQGYYbPRJTH8bydI9xWjPLfTkHRV7MV7vhGDL4hejeTZLeTjKTN8tXElQNRqK47YfA
M7rRoBMhZbMbV2OkX/kvaecS2peKsPLGmetcow0/I1OmoV/yAODe6B4QiYN+e9MsQWIBy3wUJOst
IUCahAf4KXTsmvGmmIzVwa53B3mevnZZGc8zu00Wtimou6Ng+iiaDYwpFnrzSZCz6Mwe2QIfuRAS
ZJkBuhduk+tEgM4qA3AR6oeRgptwF2YqfAaw4RDAROJNRlSAQwzLpsjY+vNdMW/zRv9FmQfuzC2U
vx4CnPnOM8SCqt8i9CV5l0WpHcR6e0rVxcaIp309/tESWIZOHn/hmWMnSU7hEHrpnfp+sWrMrNy1
rDtIHr9JCs1TljT/a0zyxxLGHCu1kANYg0817OFDRPG7Q16dlaXi7IwppGRwTZ2HtGiXtuWP0cnZ
sCzjfQD+AkjZEPzVt7hZqE7ExXMZa+UrczcSnrSJk6WZOcXK7h4ybkx9EHe3chqHbfn++aEC8aHT
SZl7qUHHao1ZS8fRBMyIFEWmBdGA/YwNxgJzREUhUCkU+5vq9Z5zDeH1KzFLDMe3dtpPnx3Y6Fxl
smZGtM4DTWLizMTV9Pn8WIYK5utC4e3GdCesr0qNLzx5+oF3yJiDgEzpzbZFWc4Qg31P9A8ciBYR
SCm3BLhaOFOvJidbDnVEjbtbl7EG1TiyvKmSk/kN71XdIqnvOrM4A9L6UA2VvRhSS8nJU5Ybwvh8
7gRt1KbmeFEXoPByBFNXIwEXnPt3YzKYB9zvV7MW7AaoutZlFZRjd5ktpsjSYS52hQXeo2UJbqhq
sRuDTgJPawi3VgGYuk6e7iU8u0W5joVRCjlDcKypU85DZKrnHnUWLv2BD9y7TUw5CDiC1dmbm/SN
jaYkKY8LWKAER0SDORafoqrHQa+CeNebvwuA/efHipo4A8EjH0uLuyQyZfunULxm4LNhZ7wb/xsO
hCL6mPmVlh+gBoItfRSLFDgIAjdD5Di9AWNaMG1FQpwRpsSogh1JJdi8L7f2Hb7umgijFy4PJNGh
ZbE2AK5srttSYSDoVg+ya9lw+sSM54SbTSZaE21q6ohk+RcTxzKqGd7nJsWkgdf1u/wCNAGpfo2s
4fJnmHCA+a+AYrXrMOZawYh83fVK24SOKeRuGogJNl2p1fTrGblHYihIyoA/3CEJtHpPxeqNVRE6
8QgMhuPL3FsoxPyRwDlL1Mk68lD5wQ2TXJ+UfGHsKNUBqzyHEpMmeR9n1Otl8qKuP6/EFlKdbgQK
lc5jZuWGJmd+58u+p7kewgvBcGpp57E85aYvYB2EnIN9q1BM2Xk1MOeQAjI3fhyOTAr1LB1SfEoW
ESCiFEEwOYWFHZZY159yuzju2JJfGFwV+/NYKH/Wsi1ccoxfsT20+Ckm3/lxPXi1rrc3DYwUgwxP
SeFhSh1kvEBitMB+ZATxK8XBHOU0laJkhUndsayt6PD4Lw7YgWNOCcv460uNWdvzt47mot+Do5Ui
7f/gnvmwju4sSc9JTA23wpmF9QIkXv0gFnZ0Dfb+WKXbujKsK6tBoFAwNeaK/oFPZ33gfJc8tqdH
fZuy1Ei/2M80ZZl2KkRE0p+ekHCi7xNUC0KrBCJ1k6mU/EBPZyUqhcd9qJA884TmfmBUnWhoQoPC
X9frSErKWHZVFdLFxNYyZm1k07OryBpa5PvHIspnrMgCo6abuPxPC5Pa/TypTU/tgBuZRtueiMzR
Kj+bT88j1YYxPpPfV1FI5db3vGuHzQAP8t0uUnUZbfdLmK2M+yFJpGHnrq0+7lZKTeMlRGK35WFy
Wq8zYz6f9/Wazshg3jHkwAk/bQBFv3/SMpE6svYbpCvZaYbWm9F3kdGQMgHM5VER/2T6ZRLGi0q+
K3joUQdfeGs4XdoRTLqFDtd4nZLJi9qjWWkY75/r8oILIDNhng6is1XSzdHBaI7rubbPEXAhuoVZ
PGgGF1S8eHaCOdA3ZcsIJHDqNCHep5fEGizhm0HxZ4qR7KkqOIQL3oJ0PDkh4pVYX9zMBsuln/nR
/BClON2bMIBw8LTK0GdTXXBc8AE8pqvm897GfFKhAnUjT1agE+CaLFPhY/p7Wntgbgdy/tJuBE7X
eZSol28iiln0ZCflG5cGrt89hm1DuKN5jjS7Tr0EyekPdJ5IVLfIPNKfS5YLhXZL09ekxTJ6LJIJ
v4oRj7FNCceoQ/kKl41g65uTI04z561/AMQf3kPQepCekGPH4FiBgm4FCT8vVBkTV+YJZJgZAr3K
EibqyZg0FtSDCwCHRpIkRddWIwoB0XyZnnz7enTfPa5dZG+HeifMdXx58qlHTNXD+xZjoKfmDm6m
s20UAC+7nZCgxcJgV+xYxfXE3ieC3VldzptCi6XIUYD6X/JYEvsTcyj2JQlIrZgIvE4VRzrMZe6H
oESk26IQkq8Bd0Kn7AJpU2ZtPoQlP8oSUqaHqQTMCobz0qUQxv88gJotF/mOD8GMHBV45SY/RFHK
4kNwViDeKbI9RlyfE481fy5robYR0OvAQ726CCrou2M4N4jAfE4gGYsFRFYMJXPxjQh2uiA5ut6Q
UJQMVyiAUHgJLzo1jZ8IZLsSU9BSz49vu70vW0njnfZOHJ+n9YvqA5DdqP6Mgr8bHRsYzAFy4dkv
bobNfgzhuWPBLELwLajVw19nFK5vdHF3NgFJiJzZAeCmlxcR6+LUNTNG1j+yCpyDLjZySSnm14Mf
khyKgcDgDt77DiuChgcNdiO8TqO2AXTwADr6m1udc/vrGiej2XKyFh64sAP+0rHYs3mJilrTGxWM
Lxdy2FbWAFKCPX4lTngkWIpcRncbU+aCW5P0mBdrEqhkcBHGHj25Hvu+HIpqiAUFbnpuir0DF9Qr
D5HyuoOdId+gqq9NAy22mDKy1zkBascoGaaeXQVZAN2TwxAjn24Fpk09gQBNuo5n31+Roggokq2r
SOMX3xVWO4JPjl+3eB4bidLfngmUJj+9I2ttAMVHozJdRLcBDSZuyY6U2p8GDqyKTrrBQn46iYVz
Dam6T7SZpH75GWZCCJaIDW5/Onwf/7vzRNhY8C2CHLkENtnlhTEfbKE8dDn0tksyPVkLTs33D3mG
ASrSHZLLCrwlX1neTjiVOc+hF9+0VHbuJ1cZYM7mZphNC+YsyFphiIg/e9nHCP+xNBzRTrUcu5gm
LBKjgL+mSPEaXzfy0nA0x9vjWbNriuE9OBTIjE7J0rYNNFkDs2jPZNKsvc336lMCQvg9HH5C2/8Z
yVF2bXzmAt1PTd4C+Hes9fK1uo/kgGn8pN2uWQ9JjBFkbGRmUjyMS5SEcHJn9x/pjlo37ctqyQgc
wdY/XPq7st8lN1fP+O1FatK0E5bUuOo0rYkX3yuj3d5rKi/O4BVjhQXOtcj84J8/FTNreF1LzF5K
8LyLCQzaUF/Ki0vvofQ/7h6INHFH1BJHuK35TGZlCoINWT2RKcG4b17qAUNLz08RrL7Z+2bgRVcd
PS1DC0p4YJ2yCZ/utczjPVMNIccONYQRuBXyhiuAVuvBxHwz4ymallWijXlw1xbJpFlf2BmdFAd/
9XyJ1wQgOXdDOcr05WFLBD2JM14dFI2NMT05AM01bY7fLwqMv23LTm1tUxS7wYZbZFsnxHkbmOFe
sQlpHoqDtgmNconQFQLAThAcM8bk570kH38OJ7/fiLp1zW8OWvWxypYuCImjZx5u08MCacpFL57V
GvNaDBRaueMwYBe+kDE4iEEWK6muZ2uJ1xkyD7njXeZckmIU7Aq5/H3fFOFG05/cpkXk2neJGA8a
3iZWLPdnEec1LXGSpa04G4WgOGMl52wmcaiEU4/cV8wlu3CQZv+7BBd5fzzs6McJnwsMWtZEr6N6
ezI2vYg+ISlaYiCQCCrZU9WxioM+tWaUDUWOP/7fT+UsSwMLSHtpqhpzga1qD/Ts/RnN4PJ2yrPp
8Em/16PKhudmoBcEb96ytbvGACwSZDQJyPq5Vt+Y0CPcKTcbeHfkkNxbjiMK6uq8gFjfSJrtQARs
vi90GH/v9YNDLM759n2YSNadD8CFEP1GOv8CEz9Mrb5ipr2Ih3XVqmSMPgCqpUFt658QA6il55pd
FvW1+cdJ4SF54fkalmWt1MbWxvp8BjSU0LY2nHgSMXSty5j6yckj69lOsnV6ff3K9bEJhr6oEIpl
SdIKXeQjUHyIMg8s8GImfboW3o5P4IHKBVt2z6onyTNs+TkdOvu6wzbHZAB0rijLvz4O/jE9zIOX
EzPQuh5OUqD9TltHm7OgRgZFJKP9FfdFoiwlQ+NFE09me2Ij1PIKLoPzpFEfYQSobJ3488J5Llnz
ywXT9tZuNnV5hck9aM0JG0gm7zQGBGpGDBh/a9G3A36OHQOcTkZx/bcc56NZW1B+jsmRUIF0kp8c
M+Mv+H+GKEJLDrsuqv9pV0GTsVDBJSUmtcHkf7ebXgNo/l5TZVdI93mPgYhyT1nuNe6Ou9po4mRr
ZIAaBj70gnlj0kVSPui0EYoX5RsaUXltUhabKEpqY6By7V8W2xoJCTNuCVKn/7JENWPeBFP+wGPY
OiJEIX7mattP63KPcKJFz8fdOyKu2sEvqhwEVVoTBbbc+hi9pZ+YB+dEAu+HCrfC02A0U3IBoJxQ
HA5o9udB9AlOz8YDdLp6YahnCbEk+C8TXusHGRSGgjsEswSx+f7MVv29deP1fRKR927FqAy3R1Gc
RVK/M5h0RoI6GEfksLi7dfKWyfHMHTJ+a3c+sPHR0+Qithh302T+baxpowq7tprdzLdgZqmJJgyw
M8PElsieAmCMvYIdLUdTOoSOx9Nbfqf6f5JVNjjvciz59OH4zRlI3GPPzEE9V+QR8B20Ajsv9Tyz
TVjGYktKdmGmy7SyEcPGPKf2NdDUB66DXmqb8BJA3dYWnduoycmoW49U4xoLUIlHEEG8Z9gDw4i7
82B9qICRem7BVf9XHfQ9ec+hLDLUpyIf3GmJyRIZnkGlBvAG+aRyY6SZOdIoFWXw6zcnWwkamCsQ
McMyS8CqME0bEPJtfVvAZVWSqrkCuVkT7/3jt46C/3eMG0auzFtJh4ggE+G3HDTYJBUFaAtcGb5j
qY7eYuCSqkyQqzFMa59zi05WeEGkBepPrVfhi6mAVI2k+8AGpJ/uQOf0xdHFga3uNeHqWwQCkGGv
2fcJP4JM0+2+jZHuFRfu0q+MGzYFzMCREuW9DLedRVscx5EPvRrrUeddVUKahPRTMjWieuzqEP64
cM5OgN00MLmsj4dAcmA70HIALiRtZVrX/ytBfnnOYi7+lHDU7EKPK3gfUXUpus4j8Uy+zAt9WzAz
3xxL2NxrDpZA7e2cpuL8pzWI7I84L/Tapk840tKJDmTgG3Q2n4qBmzR4o9wgCVm410xsU3Ih4uu6
5E/UkSTt6Ghx6Ne+vN1yRCFa/dboipo1UsYBSaXLAEzWG31OkYOZQdM3l6FJ98juvvoUs2OMeAYY
Vh/L8bNWiy+E+M9OYwnLkmfEP6M5tJTa80o0MKkKA8nXyRgNa/GUUgjzRTXOIXIQwXfzl0rnTgKE
a5/nVl8JWijXfRjWGd8T+eV2makyeRPK+0wyuAn/2iOZVZsWMm+yoBWmNitDvPEKvXK1lOVE/ao8
3INLqeAta0gThNbf7Y12GEWhwCGawvJyFwOOYAcguBPOfiBQe8l+IVlsfDZfg0i8xshv2oVdRwV4
id1A1FbH5BIdFIJqOy+TEljCccYzOh/ppZA1JdoyGJ7JhgE1dJa93cVj9j8FTQ5LAfPORQs5mlxu
qShPvWsqrgSU6NGdrtMBeGiojkbmWTf2nvBcx2tbo+7KrCi6kBcTQcTEytdcGbJZXHQ51noYz1gY
kgnRqmBpWTsWSc2AjOsNPtFE/IChKgckd2GlMwRjRkfouvB5akZAgDSDWHPPM3exAmBFmVEkdJ/p
MeB4tHNC5YV9WTBRSsqgz9x64JmBrDCbOEUU1gJW0OX0M1fWwGjSLLezrm3AIR0metHl76Vuf0GF
A/Ue0eVLRsjBSYummyez0co6GYWYGE4fpVu68j5FYNsmPYLYqR6g+PusI/o4RUaWt15JezBJmZH2
t2kMflJ0HLDYjifkoO9SSNmdPww7IQoJyyHsSLMaBXPzX+ltmgXnejaToQ+woPuLQFKhG/y6ac6L
yeJI4R27Qt4KdTjWmU1AFwwj1NxEK82/lARGxkbVnWCRP/Tvr5BjZT+VqGDcXdPI6egOnPnynGb4
xbTH8baTyOLSVIT4d9DMkxl9uBYe/wuRJAGu6ZxrZG9tnvpGsChbrNEMNNrQ/eqgIUBGqc0NZkA7
MvXDX38OLzzOOPBL8QiikKNHbU5yr3o6n4O6K73mmwSlmFCF5508eAM1UKwvcnOlfdB6XRiKI4za
uHTdnt9Lw39IM8Yhe8DlTlGfW3koz3KSmap+vCUETzmwi0pD9sFF8wKrNZNtjDsSGyQowG1CSV7R
wFXqapWtrdG0rYjZ3Kaqvru+zwhL6vCIur7FCzxZhwRDCP3TfMrF7+0XZJoq8uqd8mamjgG1MLp2
V+KklZTk6FxpttvxAHf1maeVqT1YYGCpCmTU+CWGJBR5pMOnacJibW7pTF5aU9oBOY80m3Sz2qQO
GG5M9dY8IkQIbB4sU8Jo58Ai0IGEc6Bjzhncgk2k0yJpLjWnMi3u5tEjhUhDyNj+WhOJitUtP/4M
bKhboAOtPWFOk0hj0j4KGOGU36A1oSH9scvjTQqp+4Mvq4SDLzj5cpQKTQR+kxNcZ0K1P5nTDkz+
F5hY/PapObliydDj3y/cPMxdLM8ZmyB7vdWMYWcD3+M5qIkwxij/DNfx1R0FMPCM8BsFqRFF7fQv
HUYToMuCNBYOqLJ8TwwGThKc/dx4NcLCmVE8qO6+UNlrshOnkf87LkSzZHkV72CJOmi756KdLwBm
OefDm72S929+3ibvoDsH1GhsDvXwEzxRIzWa0+9dvRFrDP3FdDAw62Wy//w67/0O6PKCuvoCtOMy
sMF78ShJHLmPL/cUCE3yk8Er9ikt76XsH30tVIU7pFyf2EIWlUyWcJI9SIWpUp3rXMOqHlctAkr4
dmFiWmkv5Dto0LaLPSg9LMVpdb4CJM+aFctoTnlaFmWhOjxeXcb2LFmIHkHxncaH25X3taJsMS77
1SvQR3I9wS8YxeZ2JsHWfpQKyD+x69LvDA7xrvqrBF0L38j52UxZV7dqpltNM8hw8zyrdkmccgZS
I0UxtuP6rJLCVmcm/4jj/BbkMXiZocjsiENlkYLJBnzhPBfE6PVByyo45pjAHmdMzr6C5sqmyC/3
g/gw8VGGJ4575eS7Mxeg7gsXzQBIku2cadGsguKUPNeHgQk4TgeatbsXqtVQhwDYAqcxuzUYpzwo
eBc5WCki+rk+crfmJpb5xB14vcB/+4z3AIqRah4pzcodpHtRyGs7dbM5/B3WACeuUqTInPeygMvK
38uLDTEAWO/ngpXv+NzziStO6k6LoaFvtvPL/ZH2eJUNxC5Q2rv/tuCgkjs6Y70UCtHIsMZ7cU2X
B3JfrkJKKjzliU7QVrQYaTDyGQi4S1b/mue+8Tol7Not2lai9znoFbdbbC2rTAvoRVQCPngxV8q0
LdNg4ps3MgHOa36+Yg4CELtNdbSEitxzUivoXneAlfcZR7OOizm6A+Iu+ydejXz6pRdno2oYFLO0
zCZhIk4yyDZryNMb1oMHIwML2IvhJHwHNDDZYp1+0dmqkQEnvW6svlwFo+nJf4VAxwRyNnFUq1FS
jrh+6bOF8vX8fdoqAqTckLTiYXjG9mj69WkxPymLz1wOkhim27QDlKMqz0FpuCYcfo88P0FFKXwb
qnY7WlhP7bwlKRjon3tndde5Ll/674gRxwevqNVV2+ecnCIoPGFRff1vxqLMPSNZY0MzaSKbO7Oe
5rkWh5+sYqia7a3Yg7MrQdT5Ds1Kx8o3Yj0R3Epx4o9+hlAOjCX0CuRx0ul6Zcw57HuVoA1OjGCD
FFauLYTzHi1eIqdc9Cz36Lh+M5RTW4L49eywgYa7N89gW7VMc4T2turQHRApg97szxLXzco9S8Df
SP1GMhWxVnTrEnPMtY83K9v1qf2sI/Bwa6Wl/FM5XMVo7m1cDCdlrsTxaYEeiCehk6oFSxFtQi50
OYEy+ssSj3/gTY+lzFStE7Xhvq0tRA1UEe2nyKddpwQRfwGVkdag0GW+/8imSMY5UdZnid7AyuvV
YTYiXaUShWdGUlgxz0D23tHrEMFWWMZfulLnboSjWyK90JCpqh6CCZ94r7crdTwgX8cU5iiHVt5B
QIyl+ajJvd2mXe+PrXLokr6B8NUfujaDeVhDAy44FInP9nFi9SjyjbnqAtO6wvM1D0b/HfG328YT
fCziDqQHJr7KSoSwQfnia2qyddhOqAJefGPB/lMoohzJBbm1nxQUCtb/3+CqXK1JpTmC9m0OzXxI
P/bQ5wscOjVzBE+ZsLZ+22yNZV9MFqWpJmTBdZGE7uMIGSa3OcsUNRVF6i7bhu6NA53lbnniWJgX
XqkkyX857pCSS5sbnwwpdGmsfeY9aL1cR1Y7XvCl5g1S9ef3hSPR4O2uns8glV4sV8zYpUDA1BAF
BGf8Z3cuTSGJqDyUyeWo+RTU57MhfR3qCBuvGfku44uCXgwgtqD6cryKfhGXgmuSMM35mdWCUNOP
3eSXNcaxInyJkyZzo2fN0yzhN5MlB3ld2Q+WbnXSw/O93x9Qi5bVT3AH6UjcHsDCXFtEm33EuWqL
59fdqLpM8RROzTn6QSJ6h6daO/LG0EICmJDGt7S+0ZniA0/o5psMDfwF2sK216aYi+I5Zn30+i02
PKi2QA2ahBm6g8Hb3AfbLHYXX3vpzzVMqG07KoX96zStZ741K5pOSJYAPuG+PXCfgxtXJ2vjplNU
1YeZGh1zcgPyhwYxo4MPEdxlQ4Xd5a7met19/GzDd04Kn84uQOHMQu8EQy9G/23iltVGhozILOBx
2tTng1nSzAhTB19F96thsYiHDbLhE7IUBuogKiJhBtqEzCQG5sC++xwKFG67jL2rQ6kCSknzcg2j
xHeIOU0wsVZttJaYi6pxJ4k8UWegAKkFnJk11mIkoPlHMJrT8JQZghPZAINPL2fSX4xV9aPzOMXU
gqvdRCpzqibLATaqiIaW5aZlSantS2LHMDLW+gOpiqdOVWmEPfPlZvEzM81EmAs+3qUqc5hz7F4a
cpfWdoqMd3oQbDDFI/VeHqd5RHCZ+3IcNRsq1Z+dw+zZlW3MYFqAzrW5RjPSMj/UED0VSuprIw24
zjikLIHYp6x9Uo9d99Jlq44r59N46WAha13mT1angYHqniHwqemMS8+ZIQVi+pzSvkUPxMrXFsGV
Nv7jlt2lDGBzWs9SDbjrHOUzrJy77A2pL60E225MRMj1lroSaracKWFF0brK72dZwNq5sJsrm64h
T9zHmWf7BibsKUXonhJbzm5yydnM/8ZbWkew0HfjnzegfAG/14rjXrjETZJkTQqdGYxkJxi5F7vg
eiANxeSoA2+/H0BAG2e83DtL55+UG35HIyeh5AfLlfT1OqbQZJXc1dzVGX0EpRl7oY5wdzRZzpzc
L/q4MgJMKDcuDKZcADnO6u03/NXfdjcK3kryUccfenVIIYPYoXPezGWb27Uil1D0ibtDxfrigSbS
8qBZcl89fmFEhNHLxud/EyCZuN+1Qk7hT+IUDs3ORyW6iazM/h24mEgjo164hWiW0iensu2GGIJW
r8dUNCgl36WLcYAPJt+hFXNPWCWls7eEDmRvfEr6c8XolpuVYzmXhNSDcfOdSeiqVYRAcRquUTwo
UrYXzCBfQ1we5UDLjPo0YI20XqXJF/vpyin6aRHoYQ0Oh5JdtEBqZWqYzwXanyx6RmdTSQ9bqFrM
9RcJX/88T5ohquDd8kF3mfT0Fq4r5/PzQKv9zdUGYa8YyvhmNDxXPlu9NwII2V7n+7873puWoQbD
JSiEwKsMtvL3CGDKQ2LNzbidGbgPGAdl649mqiDEdCaklb8xdwjWdvhFVpg3lR94nfDSCq4NOcN/
CgFPiWd9SzVhCvazrAqpOC1DK/I+2s4XEZatXzkWX4Sn/WaFIFemdlxYlywFb0XQXW43SNciRZYx
6PdcUf/KDL3V/L9TXpuJdgmyzgnEhteRScbHVsnmfkrlRZhT1aFiu0XJaDVJEv5MQvoTvomHcaBW
kOXVmhXd77QJOyCwYwAGL+74nS7nfMpLq3f5mNgbCrvmfMFsz6yoZmqmhjq/ykwGfhnu5wy1jxMo
g19kvw1pwAGFzDj5gpl16QhW3UsAiQHUNtGwEAqcsF/BIqImn6pbdRzcmY66bP01iTIxyf3Wmzg2
k+Y7SOkK98KwUewU9qQIci9TY8hq3wW+0GXwsOkcIYKOIABxoiLlDCMW+Z3tCYBySIyRzz1NKLaV
ImCNNv2u1NHvUsSEsjlZtZLlv16/WailRkPDyCLdLnnocndEO+t9sHwZTqd+dgYXWfHD9IZwRBkq
KD/GpD1MgzQT/e4lfB9HgJY8gKQrQIyeS/swddUNTLpRAzuayJsDPgDruUS/VEWIXQ5udUYgDZ4J
YHCBJwd+8F03FlzMd5Ib63y09wHIwWi135REfo65HutsTtxykxhZZLBMQ29orbKO1p91XaTzUOpb
1lXKKRCCWBvu0pKFvRBszIsKjzJqncd2q/bfrYl5f5pHVtkpLRzxJ+8KuaXZWDYLVBrB3SSADS7o
+Z6jO/iy2isldoQARkeRQZf6iAPaTUd3/qyIgl1rwdoV+LmpDZO44j+PBfUHfWIPzAAh6urbQLiO
Rsc8F9gc+/gV4hicTUHT+eHViAYp95xTKndk8KzLEuC5edr50TMN/kIDZxf/ufImiI5GG8necsAY
ioHfrr3vpZpwjM8RfdREWDGcrPpWDlIkXeCabqthnVlHPdj+32GKJvlUkM5mBV7pAJgdwy/2iMpK
rFcFXNqm1ZFYaVGU/c7vvnoRpErGLwZnS9FKIKSxX5pzjryKVcEqtehYN4P8w4xiDdim0PueMJ7F
SsNn9RoBfFhC0JUEj24a1cze0M/ZGj/YoHeHX1Sg+NMbupmL12jC/N9Yez1QwcpKJkuJP46cUNVS
nSFNgwaxwSIR7lTWL1vBdT7hYXXPQHoEW8ICaCD9lKFau03X+0LaXKw9MYl6GndGsZk/seHc62oJ
lduOZNnbVTLW1t0rrGvD3ZNAI1D7ldFvZpb6e8OpT2zQx17h4iNl+OeMXNMi1vpYWFmdbZcCq34y
RwUqwzSk5scb0ccRywI2ot66gVW2uRnU9e4gVCJn7W3NktO56FL7EeXJJY2ZD9kFUrMokRXwv1zv
/FfMqEBZr7ZFnm/YsWWeEUC/f8vn7qmJgL/zzkyqd5jCW2eRIf4XGJZb5FNFptuKCOWyByNQxKMC
QjZE6MIS4hdh2i8UEufI4oADulnUYSIMdRXpUpTQwpV4AeKBJi+jnhTanvJiuxXX+drJ+7EyjD5c
gs2iz4WD5OPaOy4BXWZ66+q5GtSOEwZUV+qXPcIeLbipPVBhn0YGI5hNzucxDZxzbhbnrBCUxa3E
pjaCrbhqbuqJSlsQNz6VTALDqGDSfEwwEahRXYmtb6ytBusZSPioFDFvmFlzOnlnn1uK5x75xYOc
uddDDSqUm90zMjevfyl+08DiZ8MKMr2unJ5XzBnRnrlCW5vtJLE5wka/6Z1yG0nui7MW4npets05
d/Rk4wtOFJpM9bZqI/UMIkvhC+06a+EiLZDqTDBefeuXfhQ9v8DpgOYpwxBU7ztbxmqJs+CHXFAX
erYdvMrQnqikrDTLZdi21G5Xxyc/86n08ek6/XmkaI0bIy5xcTqQf84I2Vsu1B16jJDk71MumBoU
KXI9DQ21zymmfLGmvGHdUeg57uh5yFFJtrWPcyeLcsQbw+nwiJP/Kp5bcjv+GPTWIHsO6M1OR0Ld
ZZSjmRtuCnpv1yRwZWPj388vKBCqLAEptRQJu+3KY9Vs5qKS9/QAnP5WQE3Xv0ueWvvXnc5Empy6
bkED21Q5a+rqZI0X4a/OdpGJdGHpGBTSM6sYoVJEaxJVbNZrT0SQByXhPh5fK4CBpvFXSHmd5bM/
dhxiWQCAUtBaG9UhSeaLExN9HFeWwQQX04W3B78d4WAZi1Qff5fpxwSkYXY+ZOl+dzm/gdzGcJSO
aE+YmWzI9CHecuewmSxPjvh+dDxAswpAD4hEuwArlFpeH2sLfbiH+CE/q1texvZMFkt4biO+68Pq
JOKhtbcmLaOYRdVwFglufaZVd+MH8jlHC2z4n9ovpT2ulf0BOABS379ZLoYKTIDVIrmL19KFasSF
0cliw5c44UiYDX9izR4WxD8X81+RD6gzq3Y0FWrkizQCH+6D5h4VBlqbl+lDzvxKN810EdzG0w/D
VPZk8b9yHvq8+a3/K4cKl4angdoDYZwYNzTkoj0Oo5ZW6j2CkRmcvNFgB/F9YlLk1biYgWmblhJX
0eiMT2dj00yZZhuNerda4ICK1rBbf9npBdJBrDq1jPJzjE+6AOzOi9JbD5GTJebx1ypNgwAc+cT+
PY1UYhZo+H8AiOjiC+6JWgtyJ+qiyv61trQPPaa15QKxNSmfwRL8xozha3HUe+X2zAu8nnMItF7D
/yhp7DOtTMEg6XXqCvYjnN7GyxSY2SzN/e6EgOM1KtjOblBYxkgz+bs97Q8Qfr0OR8GDQY/apa8I
uMiYrLFLwp0hSp2NiQV0nm4q0eWkKiFYz3r7Cev6r/zV5HLH9pggBrnV9rqJG7P4LTEqAgE61p5m
5pchEZiXZ0fSf6rG1CwlL9+bvoqKsYX0w1IWMqyleg7GNI8uphfi6l5L3SjcTJ/W5vMuEoS2kpkg
kMQKg6EB79CD1UzUvhu8sjJKENdZMmKlX95+YchhCEgK3BeDht14zOCqE2CB9BEloe0LBmBvRqcQ
oi05Ar9iIx3eTBKYJxclX1zQzQEGSQZb+IO6+IqN9s4AW4YrFqs801lp/VsjUruzSl9Lmr6UZa51
o9oPlIz3K7rw8aDpOgVYtt2aBxoKigDbGr4Yy1RRsTtIINkx7l6hJTP2fphaClOvc61cfwzAt2mE
8sazXS7BCCkRtz2jF5ouimzbG3z7T2VGMjqkWmcNQbmgJf9Pk+nCyv5LdFEp09x4P+uW4HEYwYUW
5MOh0mpVJMAxwY2OfGx83uCjAxOu0QZf2v2tEGijNQh7UsBr+GDG5JUGm4zsj8qjWXuZm6nLvPTw
BVFeyMKkTuowPYbtjuG71314N9lrAmDgnSRW6l1r7UAZAB0KzUii5A18Y06hgP9/86vFsqOz8fsg
JruRCah1fSeG6VeMRajxXKW6Xcvy2yTNL40WIUNrUr2nR1OYqR7PAGtO8YVUTlHjsTXq5HkElX6L
qXEEkCsXFFZr86ryLbIEQLkH6X5TLx5BQ32EPsZINz815bdJDDrk0Xdv1djEbLOCL2iDs9w42lBy
GzNpvSRXcGesDpXGJkZeyEA/r8xuG1b89FIxKRrSJBB+ODwIuT/vOjoD1DCu7waElrADj97C/EuF
8gR9EAyHTUuKrOxrmcSB6BLwKWJq5uYq8bYH6040nebQU7UVcC80S8gFX8V6pJVkWVgaHNtxYfc/
xLrMlenv6io9PfCj3N1YUK8J5PE1Wc8aRE5Td4DgjqfnHaI1zYVT4+8pC5bZBVCpPAUPeBy8uSAz
xawO0IkwABMvJmVDDso8pseaMTv8dtTQkIsZPu51T7Q8io/9G5K0Ielc6V+ntrnFJWYxxzAPFxnH
MbsIdt/rWk16tm7FSCo0UixvEK0AQ0yuDQUJ/RRTMzxwEP1ml3iKu+Ao91maR5WrMfFPb3sc7t9E
kajup4WtWPfWx2q6Yowh1uxclz9hcWdOgtoSYIOH2rjU3Su/SvDVXbB+19MtCAyS2puBjrKWyeop
P2UHzeJ1jouc1vgYAY7V9WvFpgnqcDfEmfi7J31k5gzca6cNkx9Q5dPpaBw/inVchqqefISWE0z5
l6Ts5wowb4FMZcSo/Z/IU+PGJFY4RhtCs9zzTiC8aTQ9F2pozdgqF/6J3X3k8W2i2YrzkRIzOR4H
x/k8868x+Z+WzYFeRPIRjxuF1PlbeoNu16zDEuwEnc30lfR3Jws3aX4lt68MtYRFW76QiBJOU5FM
qPP0wGlYcxsy+2KCnF7kFjOa6Zl2G/iUlWFNOzUWBNoXbRZjAivbRtPcWT6lLKfoc1rjZdqMiuqs
g4T99mwe4jM1ICYIOtHCVDnHJq0G3dYyx8AGsJ7DXn4uNrzmf3L4VvFFaNZpBpZRPGYm/pGrH/kn
lHgXucrZhm8BqFHK5RWsOEFYDnuUq825ZV6MyJj6uBGxtr22j90ywknz2/yN7apSleFH5ooUe4Y0
7o9ec0+vJnrLKXMOw5oezTqiGhgNdSG9oArp1bn2ldZTYohMZv2zEYHbJjGr7q6iD87/9xUTiDTs
Yczm7ekVgB4f6zKKUD0q8PI2gGMnXxaoP1Gi3puB36rydrGcXsgjvQRO4OMN+iv4/oKqO16M/mso
6Kuoz04q7JArGrAoosL+NS8PWrGY5tCO+LP+v9bFckOQ845O/H3YcerBrLXtpG0qaa/4Cch4/TQ5
kLPods/1wx/MkHvwBkatRAnkHqQyWaiJZo9eVmGNPxQEZn9NFbNM8vEkxjelcDhfsh2Emid3zV7x
F0QShrasO6T4wn5i19zsrJKeHcGVScVRv4ExkOfrklSO9QyXSkBsd/M0aRAtGAQdU42ufbrkWA2v
2aqmBqliKq0MYeffEXTcY4wnAybh/9CQmnGQ7gptvOzYqx/oyg1ECcHtTtQxGXNZ3EKoldYvUU+o
gqQxtp84XX0twRsYlEeFCwntI4/aZ7I8uMJMZmsEo0mInIHccm/cjdEk7A6aifOxbHcb2pzlJGnC
8xrJrk6Ce0XY5/CjsOnmfqUaATeoBY8BxHouffhcK1Nt9VdFrmvoHk7yWkDkuChw3yicPwZiVQuH
aNpkDb0v4q/psYMplzBW8VUoE9dQ7fMzELbmGFSIk7j40ONV9bM8Vd4FHFNzKErCdfJX8se9BIYK
FpoTpJVSHtKFQ3klBoAJp9gvJVO1JmAb8KVB4yHrHIvK0ihwUb0FXO94sQJ+5xnp7Erk49RqANhh
fJSfh/xfKf4pHsgZ53leJhCn/a6E0nEd5w8dr035gkHC91HAswDZtZmb59NXTmcrUwgY/c39sf1i
uXacG1r08re7epr/T0tHpvLodnB0CB3YnAPE528HfGXqCS5YPu+SMRzyPY1qmv5qAgHiuN2vy6Ln
MKFBZX8JcGNjRftPjjd3ubmRSah8DZZyEjsGk7IREV8WByyufIpPjM6oAA4ud9aC4otZRDALMg01
q2l7T3G6i0UI8xAoj9RUclmTEf7TzQ9/VlQBbITzgb10P5p/knuK0rC+COOq2ecRbaDpAOLQKMNz
HjqW+ZoAb0YnWJn9sCjNzp049p5n01FkBilJtbJ6IkRxPQofMkXZMT45gZaNHhrPfhqp108J+Pyu
74a8s5Yu39y18OGmWgtMA+DOx6qfkYHZfyGCQtmBc7DjSB9LMFnlH+RsiLcpCEZd3zz/YNPVQDrN
9+4ayE0pcH+c2rTOYGsk/GOLkHVqU7AkR4R8/jFFU8F2xtTzwfyt23/dc5hBYwDKeqjcX8rnvxGH
LsowSb97OPg6YDFWiY2EAad5V4zxh+K+qHh1da7KVVh1MjCmG/mKypKjQ8DeKuPKSaGx/DzsAnZa
Z6Jd1J6TRjW0vOeF3Q4uC5bAWui5CW3/xKTHAQ/A5LEnBBCwKL8h6cznoV3kaIfZecQUV+TmOAeN
pDZTNpvR+HvmxVda4TTTQnkWo0os0eif5oryzMtor5Qr9do6+qb8fM/n1hDtnYr38x0inr0T0Mt3
k8n9GkpEnmxeq8GL4NMYA5YzZZD13/sigmcKvtSdvAPzArB7ph9ZmYvtK7hVv9DgrTvOLrvtOl28
O0Bb6w/KIpWhPQZD16d1COc8itK0LCnnL3hWZadmpVIJigpDIlh7ErzVsK/QThsOMeqoOY9vjxup
rDV1OnCJwyOb51+I2x1NmEReQODsuVRTHY7ioT1699/Mo87Mtse+JnBQmQpHWYywQ1q6KSWgVKh/
WSn49mKqGG0aZ9LdUrJ1ljcdivgBeBF08eK18Ztt8papVQP2pk99UbgU0x77JQw2A9mwpDOu0Pt4
rAtx3zoNePzCGIU5Yp1ix/QwwyQA9eZa4k3BUCtFOhDhtFvQru2SfggCBX+zBpClmdCGcWZam2RO
1+7Rip973BZrhJmuUUoO0oyt6hMpR2xQAHGaBk6+XwXNynXiGLDlWmWHNpMPchaliNKmNZDunSfY
GNOcOpBpyA+0ZIF5kKS4qX9usqTNvRoQ+W3PeOW0CfAZk2rpzRADNtlKS29RxF7Oxy1Ev/0Vd8Ww
wvgjgUafYnMBDzeYk9EMJC7deX3lPYmgmno11SoqLtgkIPLxAHJBftBub3paHMUaoruEgZjtvOvN
+ryK1STKp4hmItDgv0yE5Lm5jcolr9wwJ7TPJ0DWVyYYpOs5tPomtkKeP7pZjgXHT9UrLXGzC0KL
m8eC4Mc7nufmUpoVBjjubKHtto7NDKWtAtMxTm0q38NhpBktb3GS6LQ2BvOtQnujsxGjKxweNynF
s84u7FL2GRixpvt2iIp1qHPManhkvaKjW/sDNL+E0tl/MydEtqVO7Cnml1TvsjOU9QR7B5gi7QKJ
Vo6LI32ZgI0P5VzjsUazualtJ14gmMrYu32d4zpAZFtjtykAND9cV6+5pYPG6P3YPT4i/dTNaZ9x
kNXkvies+ix5OoWyMGs5zzlN411QCiY92mv79YnL65LLobPPs1owk+lE/ahMekl0Di5lJiOm3vxT
XK3dpWhUgnt9TEmpN+Uch5MUBOQxe+hI//z2J3W742BXG7ruJbkfNI/cPOnhp6ZVEkpMJFWTiNSu
BEDm7jb6rrgyg7YmYOqNhQbO1k05NavFhnBfiOBBtuMrdQzZMJ8xKETaTWyDX+MjLYNYDEd5TYp+
Sh47B4z2hWcRvmPsrki2QBjTzoQQTBkOR23X8ycKB4fgnr/5iFqCGCgz8nll3RAEnRhbhQidDwCW
pTc2ou5M5VcPbkJinizmqJ+CyGkQEhJw+BCTqDQUlJg32iF53nm1L0grP6d695wen4um9HdILf3l
Md9Mx5jVyHbUrHSGDHSHAd9J73y1avbak8ZjGVxHCweVd2k6cTswihtWhfkDfYKyq8wfOy4DTVSn
MfopHgFSOHyfrFeMmAiBx6Qd+NLAWvxZMz6wc8WcK2+uf5QbkYuuvZPQLkINKc4sB+Q/ZcetBp0F
ahm8SOKHeMfGlL3/ZJP//ZNoyWDb08U2dKg7lG5GvntVyR8qJgKBdXfflUGzB7jV+Bq7t/NHR8Kt
GFCCgRf0P/w3bVV38lhwAtQK3WvBaYcvTFWYSaJm4eOnPR4Dag9C2BCpS19t6qjzjolHkC496AaH
RPASg3PF5gYa2LkuFAAkyThAQovpreF7SDQULGKqDwl0VUwStDNG0OFmTeYx+DTgX/T9G4aqHSJZ
/OeXxqmLQQHTN8S+JQwP4gqn+aMeqgmLsZc8wbw5yrEYQsm1Lhp+3HHxb7hqFBGiWwJPQWi7vdR5
32hty92HggJn35Jya8oQdhH6KGecB3oNK04IJMDIKNuADeugjYAhm/AAmiVx89nqZS1V68VdbO+0
pQb92uREfLDW1fTYXbaBS+JkYSIEeyccsw6QZ2h0xRAMU/XUFpHRMauU/6SbbX80yPdVU6ZFQnSr
XJ5JSQE6TEHN4t/sHZC7g1aJtQ8EJMPf+1UYRAA1IKkYRX4512psFnarn5VzEx4aCHGHNPQAHaTQ
WG2NPcN7nI49pYxwdhyTmltswtnQVA0CwFa+W8X6Gd2zOFRjPD3v3+ISCf4lv8zN1DzY/yvpLhnf
gmucGxhTXv/xBsUHSdazomjOTPFkWD0+OkByyBE4czF84BiKaKnDQMrVBqmrx/674Cx14ct6SCnw
mGCIg/GlKWfdFeWF7t3Sv/PXhDnVEGbxXo9Zy5h47BTm8mm5L2KvZqSpbNNlmg5U9oBnjugi0Q4g
UybNfUXl06PDEx6XlPSCv503CFP/opB3MtcF7xk5Jyh81ohIygm/I/hJIAXzNtLGBwocCgPmT+HT
fnpYtoxyk9VHcZzxckfxuG24HQq/QyRp1SctGTMUpmHpq9Dy4VWPu4duzRx8Wg9YHa788YOW6CR8
XgqML9ezXN3xVUZeyGy+rLBKNGJfAYPH8AegTuOsZp6sZfCui5fHPzSQuvDvisBVWBjEI4peGvhN
SQR74BN412I0meU4LkJxbyuWv5FDq8msqZbNhB+56Cx4XBT6HV2yVFlqHAk3Yc70O18Wz8QW5anF
xE6HgZwS5TVjNTgihFAirIKBhsxluuIlratWuySwlPS3EC0368TMZVIymcvOcO7hTRVVmteA6oyl
vx9hQUXUNT7DdOEeKTcNjsvVppiDNFdEmfY2dHBtxqDieu+2BP128sKs8c9lk6DptPg+zatCyokx
K41WraWOFqZUtjS9yDqTd54W4dYJErX7HFPqbzH118O5hP8zBu0tvhdbqb+ngc/c47iTBQmWZtaM
+vDQXtvai4KjPzya7W8PnAA2AJ9g7gyYF6avsQDZc53no5px3BzmIFYGVJnld7+Ma8mqhJwXfdOv
obSJqRS46LY//F1rA3g2ysKrpsFwLs3wSUPGtFMMyrCwFUE8uRd6e+HTtGCWSFxMW9wpIMR4AAHe
/lucJcGtUhVxgGXATiQSVxEI1JQnp79pTJaM9dvPvbzFIiRnUyQxtBm4ho27BwncRzpglmdQGzkz
9qt8GIVpy24qVlw9drpG2II6U5bn8Kf6xS/pBexzqsQhLesVavckez/uuHFsejWwGMlL9Lvyva+U
vuhaKsLOvcfnIFA2jXXMHvGnNYEufgn4kmcLe3sTKQbsrG9xXNPoKXkAhKkDU7Geop4rObrqyVgz
WuYev3jhG4TB5OvK6JsFw1HglTlCfm9dUJ45E2yA3Q+kFUbzNz0NalPlRnpN7HQbaLKWJWfaSAYG
XJ+bCc7FsNiEg+q7/jhOrymkulB2teseilvENGdwk4x1+i8NSJS5ncSfBFag4f24EXG4Erb18F1T
YFEWIt/JzUgIiLIVQqCizES0qENJfmHsA9g72z5MzsO97ozVQ4sEo1DM745p+X2W2aGV0FG+CMXO
p6TDg6n4ZxfG+dMgMpRFnXcAgB21yQmOGMna8w8kB8Cjw6KjsVOzPZL9ejwvQPNMtpm7kquZ48I5
90gsq636jqgWEv+DAY9E+vNBlSU56QqUai903W6r/ycKF8Zy+Fi2edSKW95AFel7sq7rWy0jl9m/
Us4CrjAvEvx8zoeY/2cajh/w7SObRdH79HWuDG9NgZq2lmC7D8OZC7oJA8Sz6hJm3Y/PiMwaxQAq
39myvDyEv5tDc3gPSV/0pl6uEL2bITsaV+jrY4CCFiCV6srSpnes6DwlE8Siu75GXQT62Cv0ew2B
tw/L4IV0EesDJXmwQ0YKBqEK/tq2fnvCwv2w7vCoDOvd4PvFBIq7EFAkrR1NvUvJd3dITfPMGiLE
Z7/oJr3lfju1GoZIMeGEP6y4zijyQ4YK/mN1rNoSI8nL64RxuDlVnXkAQAbJ5ismgCfXijcYBBii
JtqRuDEocjj8ntq90jJBTN5S6z2W7mEvPwDnBYeyWUqO8voAyQiJ3v3HhcfpUPBN3wSoYqbhda5c
YKSfqDYHEIU5297SBTY3DBmix2bNJlTc7fo/cigE3thogU+yovto5/Fzh8p19OT2z4ktpBgwyg9c
FJgyfHwBpP9Q0aBie0FWAeAUrTOZsc4Ae0UZhH0dDHHEwuwZtkbVxKkTwhsmjqBCf7Dn1burcFgf
1cTJxqlkguKA8TYvEbmvPYr6F3vc8u1iC4naH82u1WWWUJmcTe+nj+C2tZMIkvemF/cXQJ8FgcnA
Sw55ihC3DD47TfSRbM/ix54+ciAhjuqPJI/HdVJy7RDlbYILVlRnANFTC87PNSdn+4FZetOaaVq6
33bPNOMf95y0YmY43VFB0BtVatFifpNEJN+ziNyeu0MIqeURffhFF+MGKi2m3J/YOpeuOygq2ufs
MBY8VvyR8xPH1axbkjpFyiPZ9I4lqR7fyLQ8/B8iyWQYSAKMnfW55Xx7koghLqLdHchxlqsKV8wy
RuT2oh0HThrNnh7NY2WjnLRyXtBK5TSj6h3GCQWk48fgFEDP1bOH/C4qaQpSGoQnDBaAMSAZxVis
pSAmIZS4Wly5dGF8Y6z122lYA0hsmSntwmQbCVClJuyiO91uZ3UkjxT7TZn17JuAZ3jYwGMFTD2n
fnQv3RRdjWfhxrV05qa68aaOP8D8fD/gor7GJpZWA0OjFFPw94XIg9iIPchqklWVZkFp2IqFM0hY
6D/uFRnGmNWIVti9BCsiA2moeOUKaWPARm6ACoZHHAGKUFGKe7ERwK6UJhTmI1zjdD2gSSwIX7q+
gNKlUlZ94ab5KUvn3nO8bMztkSpTkN/VUnSGIwip3s1QXgkvQ0zl8wJT+qhMyqKKC/LLpE8fvUks
Hlhv/UQ+ec9ispX7JbgGb7SCZgtgJv6BedDpqCGxfVcXQYgy5+syHh2CMv/bwktGZwcui8kaSevO
Za0buEfOI2/FCOBEp450YpZLVq9EekOTlzLrgfd6WE57CHzvZ5HoWGyTcX5pF6wyjuii3lR0gT8g
RDxHrFiMqMUp+tCC48gul/vA/FC7becCzIPw0NIXwkxN+Zekj5+MoYDRP5FGG88GNGRvhzG8sTcL
35p2HzXPXm1cLgIER7LNrrW+BCcIG6FBWTa1zcfljQhszobitUGklP4vnAwxMOHutvy6TOBX8wEw
hiayHjblJuCDf1TcNRTRlidXCSxOqGYfepgSQYFp//hJyE9FkD9imITzA54C76LVnKyTzQWlpmlI
UjEU+a8AC7D2IWCqJKpaaddHiliIZWoz4VOD01IX3bXqWVk8ZVMHvZZqZYjuTipVEAP52DXaAjol
Ina+zhE1FN4dSMgsQw3yg0QJ82EG1rGX6cntb6OQg7Y85zJ0Jw4BrKk4FtDREf4TYTXG12ceELHz
wvsiSyx/2l7lMOJG/JcIEQqPczpXsfFkRiVymn6Ex0iH+EKTlcQDrWnqebcma3QO9C+Vr8oGqkN+
7Vou1VVSdPjl2BjkzYYi1DCDQAPg6kp3e5HR0IJ2CTUDBYYOPQuD3O+4+eauqDN62CECMOcVATE/
tQbGcEMAiJrzf41Rk2FrRyw4vCZlPushOfwWanCljz6B+keDxBCGKOlc0F2mnRKgfSQE3eBOec5N
ZMv8SqKmSgzWwqwO097lNlNpnQyuaoqVQSIwHL+ca3r27P4x7oW1UiR2m789Z6q/zdnGniu0IiqY
26d9thfCqWeD6cOHRxxWxKdgPRO2bTWYfGvoA64M+L1yYi1z0LQJkYp1s2X4pSBdbO5Be1DTQ9ml
6ACgE+Ag66ByGgKJqIOO5/cg5DPEdgk6G6I5x+O+AsRHDvjesojWXs9RcaRKmiXITzCd+SMDc1g6
6X/4XtM6yeoOwT/ErHlqEGBivJgVzk4YDlBmwFQ9fX+BoVsj8qeSQ0xixtfBPVtB91/GTmD/KRVU
JwQDB4rcSWA2W3OoAEILGotDU/QqjbCykrJIe6GQWvrglCGY2KYjSLAvDsqxG62Ow1eeXUsBuHuL
xXq9e5BTNXxrwFEBBE16IfSI/H6uvJbo24ir1bDLC8Tkvop8xdXwf3ly9p/bznIB6Lzyq95AXt7B
q/2ojmN93uJNrpnFSxhG8Wnf3pzrnSCRNqJ0oPuY7F2lCdAmNF5YjlAYYEhIHKWkkzN8NBNC67Er
i1KZXV4zrI5vwEGAvZFzGrHtMdx/ylsu+jZHhjzl/P2MzTmCBV40FQ8/9cL3ys2ET+vaE0682dWp
R8XPR/ZfaFOw9/jeOsswINbvp4B4NR6W/Xt22702iIyD7zlvtLyzC2zHOSiDlgBxEMUrNrhePMGB
3Qmxm70QObASwObVbZ1h5s4R1RsL0Ccae/Ak7BmpoCBuT3UUPOQHi2ljtVdAl30tiw+YUiVsV8S8
SVh1HYJ7ri585S31qLxcbEQ8MyKOFtbdPTk4wPziTs2uV6HdCDELqkCgr+jnkLHdwJs1pMqpZKiF
GbJyu1T7TaMshLKYow5MRmTKeU/ItBvTyVo8s0IDEN6Pzt3DjgHe2IoyyUYL/yZRTkB5NMaRwa8Z
GGtUkAmceBVznWOwJFtX3hmG53P6LLASBZl/RvbyW8RSpGYJ/svDGQ9ji6acJ9us0qfCMd8gy/oP
fGx2vl7Q6XlGBcUuOssfvko6H/heLUxwna+hwie24I185DHyxW/fC6V/D3s65Y3ng1DzjyB0yq95
QPKQ/9TlUelKuHKFyEvQ4tIjwU0j4eJZ/XJKwHa8Vg7nMLF3DlUejg+J/RWk17ioLLlOBVuGBX6H
yUg470XbN9yLRKWQZWyEdarhGxefsBt1kFqB80jvmc8+md8lxlJcDW4xftbvgsI7Bl8dNqTAJp08
Rb3pjMlPJxWQN98+FDNLRLAe9o2SFiJ3+Py8rptJOffFbVHSeYr+sb/nF8FLXmieB+iGuHo+TlgW
Fkj6I1lbFCm2ZIG4PFc3Y3s4K9RdnC6sGd2KEKREV8YrO/pTYDjcdf8mwTJ2JqKJNq72HUoO4vv/
8XVlnGIKhOPEWqMtYnY/e+0TR744JJ4x3P6UzHlJ+TLqcCRe6PRH96T/NZNWMapl/3tV/0O5+b+L
aGzCEJ2C9eHMt4mtTHNrr3MCaVOXVpVhf0U4O+iCCmcrz5pSIYX4mNBF0b5a3SWQSX5oNrKkgZCh
FbU3GzfzjqGo/1Iznwx/zMu2/ZoB+MmPKn/ii3S1wEQVyNax+53DS+vAMHhOqaQfLOdniLVxSk5D
KmqRpdC5atPFIGRGv3dMb9vnwDJhvEc2+np0+6ZUgYALxZmhX+0br9NhduhfvyS1dYinriY3PuQD
J10OnikFcAJJXiI0Iy3fCiwQgrHgyuReWNHNdFR5drPWCN4K2/JZsPOo737gEQm3mDGv8adKATnL
EHRrR9g6k8J0c3ObytEE/kFssZsy0Usk7hpnIOUzHvFzh50xOdiasMjPaynFxW3VeRiY0Fa5geB9
93m7/g+PdledBZSq6yySCE9duZIfVkCpdTsIoEBw78N9D6CndDTGiLkrm4hWlirgcchAuwulSLAP
dhttzDB7g4hlDKqPUt80DvddjJzp/UN6qjS6o1zEDeXGQgVbdvZc8E1luAD/l8Pf3YnR7wj5Ufx8
+WtrWLNRmjMdnXo3hhV+HFhPoONzuoXfOVqRuCVJNLuUi02CnPVRPjqAbNXTVUaDxzgBXdTWMRn5
zEPuSX9M/hsyrTEizxGC+s+YSF4v0eb5Ok3BVmZqjNHyO7Ht/EWeQSGo63/e94URXsg1pNdNGFxl
6IcD6tPIw44ZdTd+hGvHWGS6cA3isX/5yuHxXTrC3mQg9wyzGClTrysRWNDTZvTfr8TxtcB8BWYE
16tVVzMS0N6mmeHvhX6sogRo+nLhuqpMfCuiNBunswnS/hka/op48GszUimhszIHm08N/MJW8yho
ZISxlBcvek4wAip2dewbBj9ipARJqvUqY6p6azh8XSFtiGP1k261d1bopRt20pyXQsIVmt7OGXxq
UGjrwreZhQJD/ccDCIAyf0254QtCW/cNh6THCQwgTlUB0j8V/ibbtJt5vfX2adOQm3O6ifRBqyar
EBZmt6mUoqlmY0037WQjdF9P4CZghBpJhKrROoexp+gcXTQudZZ9XIgKWgrV+4QfORDwgEBI+veV
jsTDWEW4NNWRANduZPe2FFsG8Pe2QhETq/sx0HsRzsUByLMlOVTNBMYM3IsLDTfi73SgndT+YJos
ecN6ZzaX0upJm06Z4dinoV/TbZbgkfEW7cJX0/H9uQcwZBiDPMK9c5AGvNlaXD4GzZJJ2E75zYVP
I8cZfucStxhrvSBKGvKZR0TU8SYxkIXiTHhm2/tS7VLI98PD+jIuHWQisVDIaZzh7Uzt/VigcIN8
fAnY3Zt5fk8DWhBoQ+FbKFKBgvzxB/Cqejl5f5aS3pxFXPkbz3La//x2h0lOXY4gxfxZuYscK4wV
mCP3zGjtWYnNO4i7NqiyIXqXknPVvgg6efJDkuoCOP9aAxvp64mag0S8avnWXHodLVWoJLnoS1na
YDmv7BPIVU2U4ehSswrdMJO7QtELStiO1BrX0gvAFQkQgl/m3n2kN6NLMuKOfYHODu9qVLI0dkOJ
JYKeYIw0tYVbG768bFC/ybDiZ1qWqhV9AzEXwvOStGo4CC+/1zmEWK/FA4Hs2o3rVnF4mxRN26mU
40LLpeL/5ZABDOjWWWv/e/NaeSa6MiJ2SazIsa+Nx4Ky+9D6GGFuGeE8fK8qJpT6XFWT6sbqedR7
NbxXaCr2a6Y3cMcyXxQ6I8/aIdSqwCknR/oYViCwTco/ehe2VRZtueJxcdzSYRn/xVJAMbqWUzSB
2Ae22ttLON1z5bSaN4silzzlEO9kS8i5QrL/jjsMiY+k2eHTGMb9hpJ+JXH9Liy/jSh0TItrdVSm
w2laDiZC8irFcXVDLhTKFJMur2HYQf/BIVTGtl79BTNzjoWMdntrdfZJ+hCi8kQXMPxznFNM1BI2
1wRuFK9RWoqJne6SKmOfEnrhHJ5WrDfIJoL6aPAI0YVJ7IUi1WoROlR8bb0AukrTS3WXfOXPMzXZ
n+gldLS/uTNPyyQaiojnVfuPydEj2iev0KdXOdNQZpvykAYj7YY4YHaR6dektE2ukNvQstvfkROI
y1X9jfROCN+0qFek9u2VSwwccs6q5vjapsXTiIrDLaSbRClBY//EDGDgeR+qeA5oKt5GP634l9/3
jH7p1jWUeF6Ig/LDbKXBJLo7WsBNR4grbYvgnZsos3LPrDslNgWg2X2EH8DA+d6jlbCZBcNWv6cJ
dBMZcpissL8q9DzIMx+127AOp/Fkj9A90zegesKUbKC7IMpEW8lxp+zfIYQqHAFHYMnE0aRoXvbj
tLbXz8puozDL0HeEUAcz6hvqu1M4bFWnBqfx2ztX7vOX9utiI9BVW6Yr4N5FcUmHZ6Nj+Jkzlb9c
/MN1+NpNbILlnfqXwePJwlTnIs1Tk2yDnX3GVidFdgc2QUdSXJ7KviAnEG3K/vgD8hah+lNPqaVV
0GNsR4VUyXNGZ4QvcI+QmPINiWKQ6eDRELf2qVwHcyfRUKpvWH+jZBLH1R4fnmbFR8okQVQHEriX
Mf14lpCUAv8ySPn7iK6WtQkYyTJRPEvCYbKfZbj2E4P/r+F7S5Pc6Kis8CAADtz0theLxjKVX6g0
EhikmOLyztva5Z+5UnZXmUXrepzQv2Wdsv+yeNqo/OJuvsRozThKwe3sMmDqbOlPHFw9tmXz4l9z
UFNi+d68v6K/0KPId+Oh5RKDntgzZpN+W6o3k433xurBJaiJK0I0KdmzaZZadrEqY+fK6Ka/SzgH
byOfTb66uvuOO75CES//dwvGbtP1740ueH5kSBUmA1SK06SJ9spawVrThDbl4j/ya6qtq4Iol8LM
mifGo/1A6ykZ09P+Ath4v1g1HQ7KLftcmtm2d3Pnie9ouQ93CFpUgj88impWYbVtYU/A1qLPLvnA
0MNox5oCCioPo2udKqNP1wbmyr/MpP6TAu3+VTJRMZslAIU1fOrPf7hPw/y9FtmTQPwPW7j2PyFx
zn6XtSqBEqOZ7scKdVJUX3Grto70pi7oFScLcvR4YQ6ft3/vm4lrrsU10K6xS44+EpdUydgcvjxs
/m0+ysMl+6LUOIod7F/VcYAxn9zVHdVT/9C8F2VksffAjAiAgnt6d6LFAH4+f0HbgPWSrtJKQ57D
CYGbIGerxzXCHAp53LTF5jqQcvhbCppETjfiWIL+fwtVmon+h6v5tpx3qG3/5lqR6olqZ/q+7bzG
vl8aHGjnDpqlHAuxRRaLsZuobPsoidbSr/ZFCNYXUQc38QuJnL8TKwaZYmzmvrRGTv8dAunofcX9
E/qkwim+sf35bSeaqQEb2lD2NCMtOv2yZ4XCAFGZkI5DrLsTxBmFLcJGntOplyliWYtHPibiYboJ
FNfDGbsjRZDQGAsD34RxN0Ms6V4fU46jDJytwvlnRFzA+FYMVsAlB8r0Rj360bAxLulvaWOFX4sy
geU4CzK9fNu48twvctcZJKvqwTmAUGdw+VK7GlK0sWorKTZm2AqiJp8ARlr7H+DRBgZTbk1Y5XiI
o1toCmaiW1Vq5ajl6YH14+MZ4Abk7zcZURZihWSoA+PehbCll0wfn7F00HNg96u1pcIdLll2TScK
CF+dk6HTZRxoZJVd+gK9UAQE42Q+SIBbkSwMAy9nKOroDMDlNJ+Fi9lrVijUndlFUSsGSJkIHRV6
LloepDllG8A2MA8Aprl578hZLAJXxUCYgLvnyy+mXBAK9UEddioV6b/pFCMDAx5m9DWvVVH7xcda
9WjmFuPYzqqcrl7b39tZhz9fsnW82F2MCZMw2FYJ8LBrrDa0I36hIJnXotZtiltZvQYshdHk87Ms
szifrA+cl4MR1SDP/RIOC6Lw0HjJQN/XdPyJDztZT5U+gWSrE9ELbfZchPqXA4P7YkkS93zdjfoY
nlKb5inLGJ9mGUFXzQ5MKoXmOkZa0rRbyQqY9F9AlGcJcJ67aikar3BceGfN2DGICspFza18qDfc
uhY1TYxbWaz0OL2Dv8rVNpdslJ3pch09nI5NR/vE8baxNaoDyV3zdK8JzN9yH4eRZ5Y21/v/3hFH
lX18rsy105g8aU3p4TpvJYY9wrC2YMo6Yv3Lwc1lrP/l9rGl9AveQWf4Nz6/z+PXbK6UmQMLaMG/
HG0XkA8vN2qkCcSCKRO8vXHRAPKBlZaJxvrGnzAVLvRpZil6WkbyN8pyWFUnWwN3iTW1EYOydVE/
WWB39vgMV13hKgv8HO3pizUKFJ5rH20yzTX1FDwlHYM3lWb1zfN+ZF7OCBC+5hjFaitQaE3ywdC3
0pMCTrchIl3LFE5/G27FYYuDAGCqlEJbxPBZcv60mPAc3TTU5ng8iKwn+tJ8xd8ECshHVCyx2CvI
QUWYn+8AkISLPmXW+qVDEfd2CoHRObkempIH4KbsM4FdS2pixynSWlNIsvUiXlfoYBGtCNMGJn6a
dV7EQyuQLCPPTK13fhdeneLFaiiyC8P4t7XD5GGiUYCABLu54X+8ivsdGx9XBgt/7Bqv/9lW0QZ9
8YUdk1vyB+2arayNwDJKg6yq0U7n/M3e+h39i5mZbhZeJFJcIPWs5R7EakHZUox1GBZFzqqmoQBC
rczvJkJ4GFTKgOtkxx5feZMvVUVvkcFL8tNlbeXSFnHQw6sqTnajXdb7qEYPtQlTFjYrfQh7slY/
WTgMLDLinTBnYvUysLyocgOVVAghUkg9ChO9Jbc1vQb0GKUSVIrdWTERXUCw+qa7kN+TgpeS9+XO
KHqlqViOLRHwIxu7CtwMBxnPI9U8AHx3e89HZj35WZdeM2vUu66jQd0MaBEZugfBU1aQEf7YXpmI
wAeDqboz6gzWJ1OkhVKJWwRByzf7YWEduhJ8BXNmffnvRJi94mI7qVBlPNfxUSpQdiKxvY+6YKJ5
YaSU2WuKmBxw3HtvVRRQXYBbGUNqxxCH4vQWnfiDnylJ2ynjKvEX1DlbbIih3vjbv1W/7V8AoYCl
mM9PvH4rMfjTBsDXjInseesdJ6znQ5Dyhk883TO1PDmNx5Tbg6m15oYCmvuC2nA+AOVBrUSQVTQH
WFXbx8iWKp+6lRjZ2rmZ6VkN0nf4MmFs6/N/XCPqUuERNq7m7hwCImLlEkOO0RvSYd4AM1azQaX/
/CMG2xo/qLC9h6Z+BpqtijqSZLipmgYVvYv9JEf+DCf9+oyZDxniHuiatCZO2g2kCa2Wiw+tWcKw
eIYaXGEVH+u4qjlHYorSfdJ98S9KziH9U5M8/QfIOBXq6MxFupfUZZRTed+vnfiIB10U4cM+whCK
DlI5g+FZtWkQ8Ky6DG6TBRq4skfSQEvBww6LTI0SG0z8I/ajUvl2H7osKaI0EY0xkiUNw6aIN706
vIRPIlkjPVtnnjzMSos3xg62F7zmesQryP9y5TJKaW1rcD9qQ1VBAGFVjU2b/3shHDEdqWLB1ET0
VKN8rQX2mHKVuCsmbcqaX7652I5Ma5Job5qE/zTzJiuXYmIB/UkhK9DdCLXbMZwgQezLyuBw81SW
wEV9pJI/4xRc1Do8YMN1NLTLYNnmG6STC5ir9QO0+t2dF3HRFeILX7IEUUUL6h4UWeU1Nn9XGEWZ
+6qg9q8/chuiGpXCNpCLkpUN3ZhtXt4PBkbxD/bVhHPS/tAFEmngRHNxsD+xd81owYHaQ/VaqCju
/cBz/hH1wOVEfYcF/brZkH/p5k23iwKyCYqZ6FrzH9+tnQsbrIEIYw6AV8T/pfKdU9GZwOmAILgK
2afFT8FG4uMHOefRRVbhwhhHKyCFR7Cvv+mQyfCn1jUHms5D6TVNG9yJTmxB9UjQA58FHVNS+2I8
3SAF5wc1i9KfIVhZI2o2iymTv8jmg+o7d4C2csdqJH79rFTOiq6Xvuttl6uGkjMzXwqHKCkAWwCP
DAT9LRperf+T1c0L6pwW8ycR6llgQ0J2I0qfV6eFeLELdsxkDRDiHjX82593y7m/lOWsgOCtTcIP
v3dWk8Eg9DeglCFdDu6HycErLjfFyJIaN8I4QX3HuDXnoODbFwoOfAqf/bQ+TILNlqth854A91/m
hZEhljsrDAFUxq364FR5fFa1rg+jbjgu6Hu5vQ5oK7GdBb194g4rzypOJxh+ihseunROl965TH70
EtGIr2abpPURQA1qjvL/7rjSapIF4Tc2ZWA2cWJuSP3ChridJCpUWsp0vBVEu6wQOpQc+lJms+oa
HnjRf7Q0x9BnFiyJMsPhPYKzFh+gLw+eaYNnr2pBwyeamQP5y3Ac9qFQEQTTPbkK8TjhA4HEKc+C
tDpWuIjM7YOstJP5Gk9kfIki5qX9p2dB1HNh1zlJ6FI2CQ0nUbtdM976k2bTtU6T0doeaMipuxMC
zvpWLOnVaqXTTWB86jZauP95ImacwhMl48n1mBOf806NAzF3yjnpltfM26CV+y0xn9/equVjb4Yv
G2tJ1BrujPokr/EQH2tNg7FE5Qe2DLm8uYr7fss/a3MDVGHRkNq0IDlv01a5o9j1Et+oVvB3IzBi
75viN2Tg7U7dMczVJTmEgsbXvsbIx7/7i1dJbKNhkR9TxXozu1+VRPTv88p6MkBxYp3YEtzGzIxZ
CePWh/fhPjeuewYsZsrx6Est5Z8N9W31bxMzFWO0YsMPW9TgOpabOR2YLVtJ6WMqj0H0px2id0mX
InKbcJZHsUZWY5u/a3GOq9fCLYNnv7Pp5n9gKKEFReTaj50ZNnm/k5fN1B7NmyEWj8848/ELUiQU
L3xMfIaSGVMXP25TP0QOcAIg8zFwL5vSJRq0QrRzxxA7kczO6PI2OAzcDY4RxIXjHcCcsBapYytq
b7K+nAoPt7LipS1NZnnj720BpGW/6lyw1+nn24wt+6xav8XuRLr8qti9TuIlDz30zGctEP28FNkO
TZSUJw8YvkPIfb+GXBeF+nx8RDNYDFjFHQ66gZDeuPX0yFkZ6ObLmtEym4XeayUwuydFAPRXB0e9
VmfofmIMG30C8vLFDnzUhqGUAfU9YM9E4g5pKfsiwTC0OmetdWJcFnYDpSQod1Yfd5stnRwWZRcF
J4nTOULd7ENCSagOoff6wROYrY6vj8++/Mj9a+Fc+5YeB4O8jKZNJGgfvopm6p6Lnl8dmGnG+RuS
2HoZYDVOYp4OceneNnWbm0sYm6bv9HLxL/qDKhTAVXu98Oadts1AwWW6bpYrSqNGwFah8eD4sS9O
whfftSq5FZITsKZTwkRzUPH+I2n7eA1BWevfTbzoDnZQz/pKdDMeOtRN4Li5CIdfNHDiADRGmnn7
0Or6nFE/jXtaZ9zmy+2JTUvy2fUr4FGAnD/MPeksV+UHrkYj7kqvgZqIqOXiL2x2S+aLORSniNDm
IKwTSV1ZJgC8wn3/OP2hBOloEnq0Px8B5bulvMWSSKsVgbozAulZSfk7s2XZ2x1LP49zpUIPfzo7
YTpJjQ6dc4mZ5qUmIkGOWEwESKA37urKWqr6PtOuGPrcJJDH70QYGeeDkvfK8YMJxzGuuy4TYIj5
zZW8W8bKT8oAkdoxRNlUUatHzllmi3tD4a5VzkdLEpwtXf4szNRy9OUOoKNSrSdYZqNb8nvMjIhR
rpE5OkKQMk/9LNkJ/yYaFlmTERzwtota0RF4kB+g7NIg/q3sfLVNGDqJ1mEf24D7I9uO2PUtxzN4
YEB5f3Iro0Ok6q1Pan6zjcR+xAdHJQUTs5eIjCSwEU0MnloC4y6dZF5MmE3+JE1DcUKaSqQzI6JX
maePA9PBT7asVLbFinYq9H1c3apR/ju/ppAXHms5gTrOo6tPedA4WQKNSOpKPiO5cXqSh5Kzi3fI
Y2kll55XcYEmZFTDM5rFcEVWseTIpN3yVL5xmYEBKTqut1X7VQ1gZ/3jviTmec0awvljIliREdHM
mVECFluZTm34Xslr3ewzdgS6gpLdxABS19iA+497cmcRbEqv5lshE2OQzaGGSlxu+NHvURmWdYhf
CKwXndR/cPV9Qo0dWQ9a1nnuKU81Y0vQxlFuiBbyQwFYp27hhfETw+4/ZqtLZHuLxTH2UMoLFvZK
cvsYC9PGPBs4BOicbmppweih6Hgiqe/bamV5r/GLI4LDWXMsYggpHcNi20xn8XekrJb3j3xCD5XT
OFTsI8vDRMXjcx6zgW56QVgDegbP8JQj2NN1u19tdkd4v5/jrlv1CsLb+US7cwx/JltM/eF68PUL
g8psu0TmGC49fgvVPla0dnl/Mj4NCmGypsYbBc1DdNU/8A+PpHfWuEFb8Qox7H9b+kXqsP4ZnBTZ
g3heeBcVxHewsVU9H+nwwwsXJFSjid8Y1BTrVmaImdPCSKB1+L8xRVPV5n+WZtffT27WR0ZMZI0F
wufkR9/OJJutilrgaG4kZVM/knWvgC2cCPboOzrPWFZfQGHxjpWNksYZs2/wBfcDYqx0uusjGbTp
GxuvsARtKIY5ApGbNkXId4Yxki3vXfMr/PH1jYyTfkolZC9LOSeJHsYs4ETieerKZKygwcED6Z7Q
NfI7Wey1/7vL5fOa4BEWzmyFJQU0dQjNwa6oBsVOE/I/UJPMrwu8TWl0uoBlN9dK0zuZ2Xwxm3jF
PTajKewcS81xSVMLLVKSj5V+yFrBgCm+lFSWwcFvV9aJ8Zsqj70Cx+8PI6jXkoDe1jZAlIFOm4z3
3ll0DR1v/vL9j12kmN9rJUhNDsXahrSZluq1/eSSJt+s6PmZF/g2arsjx1taeQhptA7dsynjzuVI
gACJEKZfRTJRDpY9M4rnoUGxncePuNMQYg3oiEFEIVARWFSckXT3t2eRTWimuOWwQYLuXA61yEZu
2O7UhNS5H2upjWVMP7KYGw+x5b9ibC8ENvrMWDikbk+vz4nb+oBSGbKPZ42lVAPB6mNszRsFFCb2
qA3vvWCHCQZtoUKiMeieTVlp5CvDQpmMHdl1Ch8rnid2FR4HOd3JExgyyjpHtciph9dW0sBkOuMR
JFo2rUuokD6sNkCcKCdwkUSRsMDk1vZkQDcVHsh6ob3Wq6YQAcEHpokXM8p6QKL2UxCpnyB3KKsG
h/B/kBf9IcVoDYTkx/dGxh0vSMDENLRoy3xNHhT4QXRbx1prmG2Ji0mNMn03IEe3p9KcLRPYVzkP
P7AdVfhcqbCIRNIv+dWRGhM9wIPVY++QPyKRPTUkWLgo/sEcSIcCM3VeLMf4FmfcyJbln0toKsUD
d7tLh5P1gx+f1R0eDBLLMyFTi3fOOZ+kZ4fI15luVFehGpwKalVBlVS5DDmKyoijqz3ongg2p6bR
Y9DcBfGZfPAo+i3DWknT6YYSRDsSboLY4TpGWCnW2lkuQsVHliLxQwZy2hmIQAp7UcCaBw6y6RzR
/91r8EYUgiovsEerAS6vboMnEAiGMUoVGL/YchEAZ/AHSv5z+2flg3y5EkFBmY9re8nm30YTk9pn
PL0n5slPDdR5T1ZY0i+VZPbfpZyLVUactgZ6aJjhvFp5/DGxJtQq9NkzDrgTce5o60SVSh4PLbTG
d0teHY79oScefyd4bVuZu9IJB/ns805dSaF6d3fBSGGqKDIbx6ROqZcHTttO0H73KARafizSvdoH
XNoWzej4bZ9g7hz2dcoIyv6oCWpXYV/5H3V0gEw096BbH+1cgUeGnUWSBa9vdXu6LMsbdQYuBpcg
tW+8/YYculYst3oXnjqJAP3BR3izqdcWUW6VSQk4fi5/hcBwxlsrhknRYpbmO917GBOqIE84saMk
JLa0Z4qeb1kiq5cPyAwvdWtqiqxJXoxut7C+U2qNLR2Q8S8OpRT4V80tLwLzAlRGgohoCEmbxUXO
pJawT3nzjke3Z57RETNrfIkJhEbVkY3T0TSBwGfX7Jbx8/9psAjb+hEhZgvVMS74id5xPwVnB9hU
vR7xQtEVLrLoQjBMjObYpayw5EQAae3wMwNn7pbgJnd31pp6+xnx5qWOdDKnC+IGyaWgsjZ4Ej70
xH+nLzjcKcoXX31lfwM8mlsE+mapVr8aLN/hlkyGUXHQpyllh1rslQP4StofdQ1MWBBniqOI1GYH
ozc0YjPgZ2cO0pQJj6AR3QTxY1pMhTQdJzhA0w0/Eouf/rQyoiXkVjPeVpquT/RqnBYmR1jnkUnL
kWlRds3YWdqYCSSEYRtKSrOYx1+JAaoUVXofRspUYvIC8NiZElVs8U/L1kOq/iDZeLRFXMaD/Xrc
aqGZzc4w4IROCtw/VPvS+Ujp/5Z6giPHc39WzWjd/pnMzSX6Jyn/+/IrPbuynngxICps00+yReWg
9Ai+Yp7alH1JvmL6nGAqTRGOCNzegTvRQy0CIvolJQEuQLKG8PspMkPCsCTxOfVrZVZx4PV0XtoP
gFvtbNQrM3dW8Ncx9X8gtZbEBjZVY75yNWr9Ftq6rccAKlG1Ep6HY+suf2IZ6V52Sf6j52az8GDG
y1IGLhSL9CyqToo5tkkdpeEo9nzwPHCtEsSZFLLJNUcEO8CVI6GTbzT52WDyfnPaWevJrYzUCHvG
rUJ1iK0SYk5wlJY7+fCredpn495BDjIMn3JCWZR9XFsdkuc/6DJalOsLFnoqt8zUBWpM95moqrV9
kC5crVGEeGBer4XZ9XtTh4nTXIDufcj3TtIp7DvAxYNf7Bge4Dw110lDFawdTgRPcU8BIi77c0bI
lh1sz7w2wI1ifgRk00UPkKSMB8Az/rSVkgQVBhHHhW4dyjrTs7IIABuyUBCj6rGvOrmmCn76jakR
Sar25uHljG0Zk9OhznDqR/rhetC+kMkuRO5yTB4uoShuImCyHUj27xIxknU9WpMsfLQ4EjcUVEiT
PA+CppdlvUjnMuClkY5CKahBLXYWC0zRwV0Y5QBYL79zVXCeD091JH4Bb6jeXXE9x4JyDO9i04Vk
R8OoqCRSL9OGshbG4BY4vHfghB+HGj3qtBVVny4f1QWH1n3iPtT6WmKezm6w4VJEGu6vkptCH5ts
9q3lG6aUmWpa2Kx6dJR7932/Xrs696rhkN4CR+GpEMAMu53EfORmUX7QbBFQcfixnzAtYP/TJYXf
I64Bif9xBlqIV9RyNS0gCYxbbWQoCVPsuCeyr57qUerhOF2fgahtXRSYaZu+4K+BR4t8VqW5lAyX
cCZBxeXHR4g754sWKFE2gQgkg3p37rhZVThYm7f7NxGqSUmX8+sTaxuZoczXcoYB9NbDuNppb8kE
QGXspqdp6Yipy33GohoN8/J58nBn8GRd/xq5zrUlcieaW1tr1BQP+r03NX9Abr9XXE8T9nx4/+7f
r0vcaQhXIC5jGLChQ5wYL5OP9tcXPe6l+z84Zu1NkuIlWba8BoA5x72DnZy6G8ig97ogbJ98/OuA
Mbtx/VmurvDo3LVIvuUl5iFl22M7K48+OqvdmMahif7GiWAa0kZz0wJLdFKxIt1ysFgkjyvkVKrW
Y4jrjwG17LfbCli066GPPZmooCp1ed8XB5InLLXy1p34MTzKi6/R8ot56QGJ49YtIkC1zN93J4Zr
pfengPui+IdVsvt6J22X/dbyaiBqTohxdNyRxyyNoqZ14YPVh1q9BfpD25d520/X04S651sl8P/A
AreOvWXlAIZANAN87K6WLz5soIJgHyKbrEL8k8lYWfnxlA+44edfjTucpVHpdE8Ei+qFp5lMOIMq
O7tOrWqsrU/0d8t6w/q7aziG9Z/A6dIWz8JTq0/ovjIww3kqvct1mX/HzkVjaGgYKJP2gg+cWnp4
l9/Vo0WW9QoseDkV49CF4ErU3h15h7g+9FAjcHG7Spaqv6YEk/4Iwh6HMmRDj0HPsr2ZwMEIurBs
lNhpLfAwDzRFzpzCTGbqE7zkG2d993227ThX2r+trag9wA+Ea0SgYn0Kt+Cg5BQ+oMajDTyTZ8IV
1tuMC0ywfvMDhevIb2wYQT+cbfo35VL3I3vq2AFkZRtkmV9MyFCuZo2B1e8pARcBoaK0Z6RUWiCp
61IJ35FBKPqHe8WxUe3SMuldDunPmFu97dowFxR5+PyOrAE8mtbpiaHaJUlbtGdWhEJ6Nkdime/a
ENQr2B1A3n9cEQSQwTjpSi6tg9TDWRQW8oe7ncyhOamlmz3plF7alFsCwgBkB/Bjm2g3mZ3WSA/u
FYiExjmC3813x6xKs+elbXCjaj/AuePuge6BsRyta+XZWRmbnyQEriWo8h3KeBXe0yISE6G0H2+S
vFBcMzASR2DU6khmfwmNtJRXRpT0TyiF2XF1guEWffs4qs3/RNcJYbUz0M/n7q092au1A8+FGX8q
/KPDN6K6Vmj8c0aKRz2nGSRPdxLm8pIlr09IpwH8O+UrAlH1Av9n4QhEw82b8KTt1wohgC9kxoMp
5gcsngDsPYS4v47InAz/c9mQ3Rhh+usbjjH4aXXQS+HbAHS3w5B+C6uoy+1hW/gedpjEZPMA+eMu
fcss0pLfg4XMdRsG1jS6yfdgSufCeFBc1+1xLDAczlJ3uTGCTywTn0ldWhwsRZO9udBKJIdYW5Wt
rTpZ8t7zgDsvAuI0QM4R9MYsE0DuafS0GBVXUr7IbMeWluxO67PiTdsrMvWGBLs2ElCZL60731rn
Ynb6suKHHJVtfc3HfJRkZKtrP1lLtMOX6kHfbUI57OyedFM51MapLoStCgIiQf+omFh61S1Hh+vY
Y5HhmauWHZpJIVGtsB/dbWw3iXYWRihShwO1PkeoFzsyJ5uKbZ8VyJOM2KxStRcx/QQxsXlcjc9O
pYM4FmAxV5vEIeyNxGJEDZP/9MH1dEVXTWxmbAE9g+FpJzKzLkGMjQ/8FfvKbjDwAZyJXGvDc618
dWt1qIg1rJEAbBj21V/S68m6kxxbc6C/NxlF/bpdMfuxnobYWdw3VHNCfyI0h5TfD9Abs5v/B612
1xGhS0QxG7K5MYl88nhChr0qeBtD03DIki+YvbH0xBDSuCKBJchW+48UU5nHmsrUxLabQv4GApB9
8IGpbaAbkwCkkiE07Q/Lu9CV0lEZlZJO6iBZ72yp3FZAhEsAL/ze70ylZMxZ0gvq5Q3UWAiyxCy9
bLCjMImHkKTd3vbGYEd0wZg0WjOvg8u5oHZElAw2JnvGsmSuZgPSzaDvo0FIvTfUQ3gDnhz6C46i
3r7FzLYTtkDxPWcdPnysTTFT4sL5f6mIhVMQrOtFhKkmtkIbpDdtD/O8zkmgvwBz1pB/R178jntW
y1o6F0kYrvPE6taC/+prK8vmv/CZLCycx+rfcyVbAIY+0J5vE5rfTO5UOY8EfAtkNwuyfkS7nQFJ
qxHNRSt4oiwoEpnW45do3ufXbOnq4x7BEWKSTMYMs1+QZzkLQMlBE87xJrB9yyexnADu2wStGmTg
JvWh3qIkXJ5n0G5Pt6u2OEbFh/lDsCgw6HIcZzyQ9Aavtkg8IMN1l7gF2QKCsoN4giOFboVh+4Mi
Ba583zn4rRPFC4Rrc8BXAvGmEY6yYDSaJxBib3QPoL1SQ8eqys0CXVpZIuJ3qpWx1pbbUI3Pse1T
V7gttaaJspvgzsGdpThn32YWuwPvr9QcXJ63K3UGYJgTBVcKHgVppbTdTl9cPhvrUu8dr/ZsFJ2s
wGU9Nplt4pmAtTupfdozrSzT3uQ8+QKR+gCQl4Xp+EIXxtNvLJzwKscl/vU/GcFXVxQUPzVrcX4M
wDkXII+g/mwP8vuZ15ldFsDRy16jBWHPt/TMMY729LthqfcLO1ZvgzK2foyNbTzfNgZ6VYEZYOKi
LSi1/vLVGK6qZo/BVU2A25hv3OkawxFs84dkN9jAkqSYQs8j+TPpLxMK3hdQSeBuNyIAc0rWwfh/
JQsH6+HqmZqexAtUfacsaguKSmSJUCODrl0JA5Ehe8ZhGrukGbDdYC0w1mpHycVSflYoPvg6qKqX
lrxrt82ZWiverc6oJWi417cz0NpK76jCyMOeHDHEtuQmCBXWzikKfj/yp5bmRb/P52vjzIUYHn9I
xZGqvUTJiRNci7qFS0ZceKloJ/0pLCm38uRmWbc7aFBHga6Vfnkj8jEV/XQH3SvW97pyntvEjXZr
Gp0QqMjkjfVJawxstkUh7je4fPoYGJa9WoeRm1mXH4lzYxfvGW7hieuHufyx6vYNOATyZuy4CU8k
CNN9+VNd3wU+epBYEKU3YhAAJqk8fn9ATn8cQfbhECQbq+DyqUKLEeVXS1j1IVX+hHYsmepjVbsq
+4Hr52b84ZjMjJTr8wUNrMY+vnsm6sSMQRgqFUQd9yDZuNSdzm8GJeN8ewYybMug9UXq42lfxigX
agshAG/Wmn4Hm8Px6rJeNkoPOhZp9NiaLbyFddrGC0VaPAVbnOeJgTDxLLdOWUBgB17KaQEbD8jp
zORoiWEEYetfU57J+FOWUv/VRhKbCyUTPy/UlCdMZ9QV3Y/ebAM96BK8SjsIQ9CFUUS2xB2YXyky
DVEmMiCTCQjbRVCsiUDwrTmnx4m6rH3A6dN5JYL+8ddE8BC8vqaCsNpFA5tPzDYwzH18cosjVQap
7QUS2HL6SO0Rrujm6Kajg2ZjNvWBpLKaUyY3zrHr75WVcUHKv7mliwMYgjqxDGCJqvfhg25gBiRd
1qu7I1Rtg6dAqvm08NZEtspwMEn/waKVv+saC7vAbTvce9xFMqx/xpeMh6v+1ttJCXsAIOnnj6k6
WEwSCZ5vCEGC8rjb8Dtok+p14Ns+VYUQdn539/vokBDKfxF7vEsFDWvgWTAXPyrmw9c0wOvfz1jo
hVJs1W4e0wAm47yZCtWGgIZtwtSUcBpH+nSuNHHt6kXesXj29fcJu1QTTgulw2nRFoWyayFpBmXi
BzjLr9r2B/G9b2NlK6ZkqfcDuPHIgTlJD8Tj/X1tY9nQcJbjMz58kBKZH5scR+/x6nulwoaywZeL
aQgXgP+PlIQLuJfvYCeI+QEx6I5gx1z9mfvMYC5WS2XqW0bu8MkJUPhQGVU1jmEA846ZPrHPDZh4
kC8FriMcqwcjx5UlrbTCHF8yAKXzN62T/7Vcgav95LoTQ8yd5ENb+K+RkVjE7d8d4OfmwiiPusIl
zeJCzf+DPusfDvSSxR0F8scH7NKOQXKePeQ/OS6Yw/z2z0doFg1xn5skApw0NnqwWISno7fRBXSo
WxA+PCvQmVM4UETuGNFRMpoAqjY1rvNmoCJXVmPXL3bpqh0cFiAw+ZZhU6jUGaVxmSOhTaLR/4jm
hg8wGADLbX49oKBof1+CJenb6pWi1wc6Az+97tO0jrjBFScJ+Keglh4LkLS+Y/ECyGDgCwODLyE1
1u8ep9hGaBiSunbzyq+P7DmyyLfgPMx4Yp2W/j5KYojEb7sECEOkt1O0Rwp0R8n7K6LpN7G8Gcat
5rCJBSALEz9L4wKClmBT8/knltSFtQ1wnGwtJiRpmEAWNB0/La0Ormk7O6BcbZ6opY2gFI88CkMu
p1Oh06FwkZhkOsgRIPPqtVk6orhozSb3x3NQkOTMDB2qiSWq9ROBqqr/71oaAm9+aQFL3B40JCYz
MrI/QlPPiBJnVO8kImvS3VW87PFq5Hn9TsPpsYiVWmqQu0ekZowRkmeVG+fc3v3WpYznjiLLkPpw
K2t5HxnjdmUa85BUXOzHT3eP0487KVyyGS5fhQUqngGGLmsBEROzR176djP2js+WnTEJFYeo9ODM
39PJVLCpubhtSZiHgAs44CbVCh3kKizedqiY/4ncVwJcG7ykaPUGMmBCbzoqsI0AkG2L4+qrtslY
OBj1kbdgLGlWpSf9f+g3QM4YyWYaQUKVBQJgLzuY72TDS4xGLK9TOSV3+7yYy/RzCbUCl8ijtJ2E
8VS6IKeMcE6XTVcq8lG+/rwwuwMuz9Zruqe7lHtxkllQ3ZHSSJ3xuAwZSc/DUjnI2vxj4icDTXZ2
W5Ne5D2IQEYBJbckjHlajCYBOWYTIL/E+pnc9P06jzUnNmCQzP5XW78VEs0A1UvECIXtpLAun97+
wZHR3jTMmwnxjk6fJwScD9u9lgJk+jde71NLAJXY2hyPwrKyfOlzXaTSdqKoqNICIeqAxf8h835e
JpNG3Fe0K9vRtPK2M7r0DwSWXc307M2gOx+7lEcrk+nq2qi22+PTKVLSzf9rVmxj8ppho+YhwMaM
sla0RpAdlbYp6ilsBAJhNUBS+JLIwDPWP6E0ljLawVmnUQFm/SaGglNSTPPQ68MTZqNab1Fmlpnw
SMJFgLH5BY1u1XL+9q+e1tr13hyJhWyZ/vCuHQQJrZgrYf5/NOocopKA5RzKN6mYiQ/zfWrScXd/
6zg/AcQ2nEm1PKhcK3cwah0owF8UGcJHN8YTCH6a9RsemaGa7dFshzy8UdTDBvmlEveEsCZLsMXR
2TgGOEMihXRdFuLCqUTKDz75bnjiejx34EHc9usffQvvDmdHE/RYdcTtgJ05khFUnWtjWGcDoV0S
KoA68WuDP1EQ4PwLnjZdoGYnU2jlDuDjxvchrb/3a4S5SmyUFFJzv97NSgPdkLsmFq8hRXxyWZXk
KrYKHp6xFXEArTFXxtA8S9z1sFYQYTZjffQ5ClSxG28+vrokE70zjOkH9QO3TPk0GzWDT0/v3XNO
rtAksFJACzAT3mNFwWFz1pmvX36i3/QgvoMdRpb6dDA4XuIEWwQ/CTQUR9n56Rpg9lXngHA4l7sR
a8R1xbTHkA4G4b2+4CdM0UVRow0T7HDOtrAbVXBmJA8R1gNV6IeHiLZJmISlLYItNIbL/T2xafO1
JmYxAlHrcFJU0kZsoO9aFhckOS2eJOw5q7yptNkdX9HXEPuIy8ZwX2AOJkkTAYKiP/X3+UaRIx2L
n2TI5fO9JbA4aPawPBZn/sQdc6JqHZ0vbMi7s1eKYHNre2TzMa9QSPRyXSyMt9UohLD/j7fqLnEg
e8jtpxResVs6yHOqRGeOYBk3Onow37KUCJuxufI5y/BJosCi54ICfi2vqdiUobPybNuaqfdEzDLm
InRchzFg96NORzX6gmjgOZTculA30u84KUrdjDXq9gyCowrxyUiun9qqOKYNxy/zOOeONyfe3qhP
0+cOJdTCfXqbX2xPY535BzUiibmTOj/kD0SIem6qIU7MiP1pqiwAFkQgFUHQEiJcMsoKdnAStVtV
z+hFUf9xY9HrDlWrIgA8+sF1kcYvUV/bjyrbnMFBUIYTIWEnfmylqcnEO2GjmPLJ579SbSMVpIVs
KSSS+rAbkn94B9yAnx1sN2gomUlrRZq07qr3ZOEPxpbdplbs7ZUpeHaitPKadDnVClBTyF5uTcU1
hXy8NFOV7zUNHAvhGUxByq79qhHxJdwzPCybdjoPwXLPd+A77GPxA/5/+JPCBJNshHKjpz6f5VE5
igDmE4JxPQ9AiR41SMwuuJD0rblvbUGVStSvokpLVmyfO/zTOmXIl+dOPEOVr0w0ZO2Jq34cg4J2
++RE6mX2suj8W2tuKU6639tBTiKSXNFEgrZ893LlMDf1UZEVgnBfkV7R6qKHgy9LQ8yKwhvfZdor
N88gavTcQAlObfK36zpqs+U3Ccf9B10gOPjfwD56bfELCWYndFKaClIRczUwYfany7QTBgV3B4aJ
6S+Y25XafEhYznlE/XJ2V7GJtOUFdQgsxgj/Z2SKzaO1evC3jaxUzKDA74GJ01cHR9rOdrGcpgNV
67GBOA/qizB3lGHA5TXgY/AJdPS8tAhhH5FbfxNZLYKhAuncjn1Zi0A3E5ZaIgR2BWI75AvFnNSB
bOOaJUtnp6Ulne1ACh+o724ikHFuaDSQ2uN57KXX4wbfcwRDVLRrOKBWhnFrkojlFKnlz27VY6T+
gY3WqmnKUXUCZAtIZv83K894GJBOOFAKpwDkkpIQhFXMUq+PPjb2uz/xfDKa27kluYdRJyLef4uS
zkyG+5HHDlNJ/3rF3LLF9jDSld2Em0x1vuVMbqB8eXlrkISbJMYWoKMNNzhXMdxcXyHd1Xkr5vv5
0IvvCyqPq4hlxEIU8aNhsdo0E2dz5sv8GWuPEjfzE09gF2YZ/wlsOUtLiYyDF8Lpa9asIFu3IQGq
ZYS+JBXz/NCDIHOVpm5MBENpBLoW/Yjwe8ILqt/gRf5+4CL08aWbm3mWJj5rNCahZsxryPHx9fos
MNeuuerUh8MagaZz5xI6q+s8PtoBSUYdB9+R7Esi5W1qOUxmap9j00sO9PMz3E52ejhH5wn0fix5
y/DarJ2JEYT2FssoevZQq/6TOtx8wd5viEDcX8MkY1qfiwH/g3OIBn5nYUn3hwG3nwIOC9wPeDHR
BYHQ9yp3pZ0Q65zJ+9T1W+1pbmpA4BDG7Y0jHY22MZvyC7XLTuT+8kEVlV6R3zgIJDS4uXonD5Wu
vUXwbxVUCODDzAznoNUn1K9dD3AxSaasySL2t9FlSx46FRUqqppQKViHJ8KznjycrJMXtrToS6Xg
mSYN7k9RfsMXu+Zyii9U7ZoNC3vneGCF/62BosemnN06tkiAS9qdNbYuD+/uAH9osft0j+VNDOQQ
mpmbXqV/jeotU1gIR4oRdDFdcgcX/c95HHpW3wH+z/jAfQdt1EsTa+UdTQsh2OhpY4bXsBE4/FHZ
fNnzkmKCNOxkqA0I0OE6XOqGRdT/PHnXtgnUUNMRCkPXguakk9jK+r4O7KRVuFp9q9pNEOHEJqt4
PFsabjQjJ4nGI91oWgYok5JwLr6Ldo73exhXLtbs8CCQ7Rkg5Q/RowQH19oMN0UFY26zmIZUcyyw
Q5TsoJHObA+N4emNk4axCqR2bud2nc3UZZoejRAYLN28M1c+Ku1mrvg0yJSXSp8rAaphy4WO7/Gl
NZOa/DGsLha6RkI1mzgTr8ZPzmG67e7+0aEHMsH1OP4dDrkeZEZxSFVINq5d10u7efqt2L0gk5u6
tYl9EDWu9AlYRZNLklJwcD2d7hx3fsXRoNcbZ8ksmrqQzpMfAVuIsqRmVPaEollNxIKALCHxc9cI
9znGts1q+H0+h7dTxO/u5XDRnB7KoGltgciKLcjgU2YEShTNb+jUkrvDVyC/gB9PrA8r0Gm6Qfx1
7sLFbDWQG5Xc1fnpUcwGuUTkYOaUsw+k+E5SEECdQXJpXClLxxjXIq9LSa/gwKeaJ1/dKR5RZuAi
VTMaDxtarswpDFC0YjsOLz8R5tbcmkirXriOYm9YJ5Jd0DSxOWAtSk7M7dQBTS33IBrX3pC+0NNI
MU7O1GvwchQ/fG2uIlksPsWaAnUJEEYOkLUWSZwHwQw33/HGJZmuJar8t2fyFCryFyVIeqPlOHqs
KuHNuDneHz2mG21V7yHWzewqfrxXvjLpv2c2ZlHf6PphLI3fr5dMaaSCJD3vHsirSt+XbMTH+wtl
gENJ2SFHfYAPbA4QRdCgyu2Mg+MeVcT/K6Vt2CX4WeRs6Gsmk3EyvaZJNBgvGTbrfpC21mWCZ4Ju
ufzba8azr0NtPu7f9nfZdcPpVeVLOF+ET9cX70t6ao7nnoNIDtoNGM3E/XgGPXBsNcGcYHCEMjNV
iAF0rNTtayEbyJ+P+jAPR5u9/3o/AhiKgZX3igNxlNyyFi4N6nFwVaU5kqk++k2hXl0Rm5BQ50L6
z22CaIzzAbHkZDJS0HmZJrGSVSvI9Aw4mGelnUK9RlyAEy5PdEM+wcsMfzsjBb0QlL18we+GXj1M
UKf0/2vs5ikjw+Ayzp99CKye2G7kvPh6Qv+4poIW5T8RqTdenGF5dy8RR+NX9DQYNCpZkKCmbt4E
Ds9sDnooMkkwJT0+RSpn6EL2He13W0wGI2ZJdIDI/gm6P452IwevwUHdBu1nACxCwr+btA5kUW/8
DjzlSg22p/0Gg55HCfFpbWMA5eat6obyTCqdSqHXSnbuG6ER7VmpAgZaXSrdmMcSMiGnBga+RKEo
kWAiCjP4X2zEgnHPn1SBfhFQ5xzqtmsIi+XqcFZMDYqD//pREy+hzcpuyIjxXAdqAbMNZyJIhv8A
4PJbKP0lFCkaIoCf52EE9YPj0eKE/D0YBLCbIWIACaSCacCFoFJP7r1KRS3YQU64PuNnOd/n3uiR
a2mpIBAcefgYtLOUdrFkKrDfkg2xpADhg5Yd0smsiGpmukFbBaa35Q58ArZl/3ga3Olj6DQBxAw0
JwFoAmMUehpYEPIZBoMfpvnV5K/DnKcUPE+gNkffdmnOpifijSLBqo0KKn3bN0SuAJGVaV7CvtEe
/4JcTgBGLzEmYZvKk31HVw5sRqYvxd008LGxtARc7CuTfeNMjCMA+oqpMh5C8QTi8W1V0tOqizK9
uju5tVVaQgVJsuXt9qXvP1J0RVKu/i29Zy361nu6Y3piXqqDfl0kRJpERN9VejvvMJ4QeDEXqAGt
BZ9XKXUoZzb1NjJ50MtND3i3brGtd8BtdaaEeQP3JUKSr8gmvV/V9Y1JyQsSjO3IBxgp74MSeXPC
hFgm++fPhOmA/FyfZF1GSK/rA8kR9k1+poyOH0NXJcccipkHgYL00Pn7zEHatcxVyVdV1EAxGD+S
BRDfsAuf2XB5I9hnhRTXi5FTniJGrZ3mcHd0ds/xnJFXwRUhwsaA4kVAGTx2vQJ/ad7ZEq9C0J+y
/f5eW8dQVK8NHVZT6jBnrwaYu8WsKJNsON2mpZTbjiNxnTVxvRQTqoFW1xgd3jueGCZ0LwcntpEr
9un5udyFiQ4A0V1Xy2BpWeVVyRxVTMoV1E8bNEPPhrUKj1a0wQF6xz7pHX79qYe1bJI9/Ht01Goa
VuI2pMOs9SPZ5fooNWobe/05l2EWnqYbiTLxL47TZdq1Q5IFCDkQJxBxGCOCViSt7G4MQAq6AVHF
0TGmtVN5INh+V/jEcTV04k9yAFfgzMGPTBKd8zCy7aL+14AvPJtD3sRz8W1Mf1tXaeDVZahAvEzJ
PJTC94TVIr3jTS5bJV25AknkZmxXaUS7fCYtOTiidhyWnTLWlNbyIhm/AlII+S+Xpm6F6GFZUmQt
VQW+BkIb/IMc/0NCVrjsH31K5orUDbX29SvKDobsQ7YKNtmkRhLhgbQI3gSPXZ1SKZWEzgK6/rMP
tb2MB8GhQFIqI9Sl/hHwc1l2YbbTrOhNOy6d7y06ZsaiYpD22WGbrI2516Zsw8qNb7ANrITX9cpo
/kJ5WsW53/vgBJ5TzdUG8mcLVytn3p4cePJiRu9aCfcPaeflR3/U07BKQCyyG4N8km6sSeu7WRp1
ZIBdNVcDcghTa+m175beC8dfIRxNgjxnzvG7Tyi+ODOhfG0ZpXs/OagE4dRI+aFHzbUvFTV2tTKT
MS+zx+CEQnojSSUcjKqWyVEXq5VbTkifATpmSzrZwTG25oQaOs8BE1XzCqY6AS6p1gnwSTgTDXtN
MA1VI3Vyu1vn/h87N7xRdVm7qPxT6rOUO04zuMhkOb/hs0VLu7S04pwhbaT5ZHN3gMG/p7WkvRL4
20IRv5XNUfAQ5nrIUZOlNSVXWJbRpPABJ7NCrVex7h8jhCq4bPMGc/FwKgQ7Auz64JtzUNiDDPX0
IJmjkWMY+XHth84C+k1jliZQcKJqzI4iFn5lxZ7AKNMd5wF40yeeAp6fbeCjy8bbcAI3r2ZEOiOV
ql9QGUeowOTBOKOasOPaF4eYvyFZ71PJRCtTVp2emHldbWMNKnnE4qpiWH5zuy36Nb4qjOOb5zo5
nr/dElNR/2tZO9KtPp0G12q3Z238rYHCxzEd8EefX0cOW2lJYNggnlF5bAnZVja512HXJp8rMmAi
yCfQuf4B/pf5diJ2id3UlhPExXPsK1hh8lIrYk/K8nY0aZ4nJzF/tsduC/EOG58SKFxrldT+utIU
oTSjJ7GhI3qQNMKJVzufsjeeUV+Q92QvD49q7sud0Lb4ObU12kQYdul2Le6QZDO3RTh6cVow1umx
18CK8ysHRdSv3v6rJ1O9Pfkd2Y71D4qUjGH/aYhRTEtSmWDOe5vAFql6jywYpNg442JEt/eOdMUU
oMkwqcXGJV0/eWvpeSFC7w0klfinVnkslJmqLvY89Y4KJg3MyCjTJDKK3gbZEJbj4emLtog4o2w1
0hBbIbgCsoVuQQXCA8bFN8xzyiv2k7O/1TkBGP70UK22T4v9C8VlyIguCgvbz7bHDyQQ78xr2Aii
7h4wHknba18yoDpcOXoKqvl7DxAe5y85ng0FTPOQon3JiEBl1fsLEdc9vBmD79jWIeX7NExTkEJA
g9P9UBlViTdwibeiVYMdKlGh41DbP9O8d9HdZn7BkB6ZRnWgvtsf71P2lQe/TURQtVRWLbVrJwR9
453Cd0GPYv/pwOzzEpB8eVb2rRr2GIj/hzexfO2bUBmx6IwZ0Zk+r63Lr5iSKA/VOQFgZJA+L7XS
h3c3CptOjWxB3rhguPNQi3GMV9ZnCueKVuUNSW/+LnFLpyRpl1zXRPgzpqOuhsQyzk4E6erlsAB2
pQoK0qcBkCmnrL8+uH3yca6wsBMR+QquMmoSWC1F/KTWaO8CAE4KhdfT6N77GrUceTLD4NBc/m28
JOcw3bdrv1wE63DEzBLVGCDtAbWRyGU7fWU8jD5L4VRoDOCQbbI3gsIBo39ojmZX5y6N7yA/FPss
ZK452Kv56W3q7H1QuKFgvwo6EnYZJS80jXGv2wt26vGLdGJFlVnDytcoi50mxnhrpZuhDsQf9v+k
inZZsKBDVBYyhgBKI/qfQ8SXhogFDNogTHFO7tkQ3yjqppv98AM2nWhQ8aY4V59UmkNNiidgoUop
VUP7KQY9+sfTt4kP2QbxjTg9sM2uNqP1qYcbaS5yew2t7m9HmwF1tRxMK2wbuogbngq+aa0irpuZ
EwUoMAlWOqo42inVkuHf0RNmvmLWTyYZ1QUyVek+WdAaCj5rVvb67zCnd2pamQ/W8dJh6eFhHQNf
cwFZGjuOZV1XqNc/EjQy19colMgGJwlhBx89kj3KKyCjvuK7I4BjioAw33ahea7CcoOtniw0Gzko
VgHPRrIY8D/63Wyae7BdPkhBkXg/OqYV53C/FoZ5Bo9yHjehT1Ws4Atdm1C36tyPLq2ZuoUcVrIt
HTf35pa6Ho2SkainmAfxwQ/5UPFsV5CJRlBA8faFxoR6sP4vCTolXk4oLcVU6smvswDhAccLZ96s
LSgnGDBj8EE3LrvhcyTr+HvSjWqGadsAFY9+V1E7dvQDqJaLBhUDJckcRTvSM1+YzqA38kFqf2OJ
/aT5j6mYrcJqr9Rm3jEJoKwsoNki0TUADgkof+Hfm+ZLIT6EXUi54+j0SScNOzGSBuC8HchD4BhW
5U1Sc1IbJxFsmxk74aXCz0H2LSbYqg2X9eQMSCynRDBIx0gQ//TM3ffSSeM/DS8AQwN79IpC6bgv
H9og1FFXGw+d1rfyowOOX8zN8kO+EQ4jlVot0S6XqzdpqYE4ngn6d+4nTIBJXo6Rte2ET7JeNU2w
5MV+lCQAqhuB7zQEheJT1Ogvz02TBxAK8tQfcs9J4uhAm9CHdatKFAIL0tl7te3gtBpG74RHimDe
GjyKOHmMCJpdNPn19sClR2eCgzKtuIKj4F3OLAgZoJB3Cf344VqxeUhjxs12Y+yAsOfWQXMs/Npm
+l6lhtH+ayT6wMCBtoXf7NTu7kzVjTgcuJTKYSVoe51aQh0lCcOodv7rU6e5Vuw9OVDotD3iHTBN
VS65On3jGmKu1nQ/540PLYy2EnVNY7GYcs/B0JEDtOjXKl1a5LWpwp2ehQTF89gwEt9uzWZJQlUI
TiKr66HvAOT9F+VAJKApg8FiCwx+AHtPAy5O/rT3lDQAFHPXDVcnW9F/pk0QStLPFH96RDekV0/x
hB8XRqXh6Y7I99+lMj6oQpJhq+8GwivZS8mZKgWcjdbLtyejL+Goi9z6m3kbVtE6KCyspbb9foqs
+VVysxUpLEYTHm/Ejfh39Pb0uj2f90LPeMBj5QNfTN6MThubwZmWyA9NSV/mGVuGOCwum2nnRlCv
YAFwltHF0J3G4UxYfGFVbdSZc1fZIOme4+ulomRBp3v3/YzLlS30sgoAixxxPjl5cYR8lReb3pI1
Qv19atmU5SHFs6FeVZnieH5YROQMlJmxyPsU83r/QQplPwgVa1a0Rx0gxYHaWwp01EeTRMMa5EM0
g4frJukferiEyys3tPZ04eDG+MfQ8z77pYQP49FPG4e2CkeFacQoKXoLqRFq+E/nU8ct72F0kv8U
c3ITwZBDAqyRMPLjLmO3rKeyxUQR9J7xrnxzAeDmUbaK+cuQSlkqz4BH/e3z0U2vG4zpQRvfnplF
fYKjWQ+gLIfnqPR8YAk1foWN3c1rgyKp13bHvmW9gchz/atjPRFJ7CLCPJIiALVHT9Odzzue3oSJ
VdoYdhOtezDuAPkR3OWl1iLAWUZrqGIiMRJWcxdthwC48h3BJXGZgCcpI6rDXIeIv7yOU16WlEEm
DVoGF00SjQI5g/e4qOmUGbj/LekUD0gv79qLISyQtWRSlfzqZG7NkPdGV7A1E9R/aGqs1AvO6qUU
w3aliYvg9Rmp6U4mDGoo0LqYcIdouBhVNWjf5WSQs/QXEmjCGuaeXX2wxQhkP1Fkuu7XByF6VZ1d
oWaXgqlY9N5sPZNcHZe3KD1onfgFUaXM6je7wCrD8eDXTVz4Xrne3f/wbVtzMn5SfX6RH3wxUpmG
awg/Jcz/ffWPmLE/njSwMGrF6zsC+Eik4HKl5v/vGiyRC9wgVtO2LKEXoaXabwEhTDptoRNCj4xr
zxVI77Wc5Xg3AGFEhO16T8pXuJzGT/9yeaQU2YZiU7juq3KXHw7J1St49r7ok3o7uy0ghvMjkSrO
1B9WEaQ/IfkR0R6coPgfQ2+QU1Zg5WCsvneIDd4m/fwhnu88yVSJ59biwbGh4gZLD9LLLHSdpL76
fP9dq9jKaHyqKLN1xx6Y4nckcwspkiDoNZNzf3C/Tzw16wxJxRqTdhhDmUwIaKXY6lsj7TLYXefp
c64s7UazhkSBwNrEy1i7HBOQ5E8/SeyRQLca39O3BQqK4DKD30GuRzoe5YSmyABQByS/h9yZ4S8e
W/xMKPsAyBOsewnWf9zuVLsEbvzq7ynxSaLUgzs3TVM4mb/U2prqWrKR74e/kN37xBhnTGtkiC9R
pwsgScaYdo2UoC8drzpTSqbQbnGr/Ff2i8WtYj23QKglaNnjUhzeXl2yKSmdTwq64ub5TIwctaoy
5ZXM9RfTUqTbF3FlidlEYTL3wxcIeF3dqytZxh8pHgBJUNEoCoT5c1uAsL0CP7nSFfwLguwRo+xv
ut/RM/c0hOoqzHKw3olcb7CGyrRcKZ/Mpd7GqZCm4E+jtcH30xhylIQT0KUSQSJVSD5KTmaWP0kL
3OjOesO1MIWXvzs7zH+a6Xws5nNoKLywDcK37HzvKorX8VYD1c8d/6tq3Min3XVj17F/0HjsUcuo
gOnNheaf++0TKa35F+iIWKjuOnWPOc6hIr005tePiTLdgTWm97K+1r9n9myIvXepIIK6kjomGYk+
neBK76HOpYh5XUZYf3ULoCnsZWlibPEXdDS2tCeIODm25M0URWr2tj5ECyBvQdfSa9VG0+6zu1q/
5d+WkiIblICb6icMHHEzDs1pL4P5NuNgnDpfzOmUN65VL2XOrhKpfh2qJV6ruhJe2ovk+64PmqA1
s2g80QmcRo650K0VKzcpCqRmlgiytIA2hlARBmROz8TUSDtTAs4Q/I5uVObRw90iKnU/xeTCe0SV
xnjAVSGbPuB5SMoK6p9v7v7EQEa4YhzFsuMDHPIYqx3xnO28CLosZH5FdGb9UCABVJ+jUX3lRpy4
7X+VdkgpL7LXqhkfEp/k3Yy3bDQ1nGeqfGJ/agKbX6BK0LpjxkSchsZXGxKet1pGr+U8sELWAZgK
FO5+iaLIUDssDec96RcFSIb19J0zmw/zSwdqsovrsPFyVo1bE4LBS5uqnxewF0Isf/9sxrHLf8HP
HSNJQ3mtemCofyd7lMsx3lfEtnZsvne9flKbuINvWpze9TPWOg3cbZQKPZj94MkRz3E0i1d0g8Pi
uy6hC+6auWviANG1Tkp3UwqDVmlCItl3Sutv1qtLunPSncIt8iedAxaVexU/OX/EHlbQ2JFYO2Kx
NiiZXl1VpELdlDqx+BOWNqS1iKtxNZ7xkw/FahCoSQpbeoGtABP0njH6ZyMs54JgDII9Dhipv9lP
nsI2VAalI1EkNfaWUlN1iGwIOJE3CpXms5JuCP+1BR6x1jUWFIOE6cJEbjavPsmqaobKrS6eLkUT
pmV/QGBb15mLF8XydnmiOuJ5/YEjlvH1z+6/iY4oBkZ/fLIIO/xNNK4+VHPdtcdLf9iHvdNXKulB
eaD9e3D/sSQy3kxAGeiIi4mpY2lobg1MaGag4IESvnz0nJ21eayRq1ZAxF/qeFkY07HFT8i+/JY6
r158tyI9yum73+qOYmpmnmVMmNI18bY7IXYV1gtgedWIeYIYS6M7RO6H4AY65L+n9S7nCe9y+CJe
ar+3MQFrComeJ3u+IvswXCDBgeEmouYRXFpB0jgyO7n80XH1KXTpMheJZR3lSiyaLuiqZh8AzbqU
bQNk+Ijo7abIZ05iOV8idc/0cb3EeQ4UmH6cmVmM76s/JPJxZ07LEsoigHrr+IMEDO8VP0Ag4ojl
XB3jTqZe57SjbwK3ZoYJ10KBRCX16wHf2nB/g4yPhErocWFeuwi/xOTGXHBEHTeCZqUeHAVt8Unj
5UO4zXCO40R0a/z9VIgOxzbthuwHgIiqQ38ipDiYL0OebBs/+0K0LoXXHTp3d9g5oCSLnymkk0TJ
JN+qHtf4FpeKdmB5fHU1Vg06vt1uFuKIsAY/Q7nsKbKQM6wIy999ZRVBS+EjPWWKB3brdyKd2qZe
QaGlcal7i60ldv3WEnoG7b8tKPYUfUip0UhW6JrSa+LaZ8T66/h0b9/Wy3JrBK1GQebB2ULLWT4O
NgAmdkFYwUvkNu7Qz7deM4xB5k/DreEqsF42YGDNrQNpMa4D/gAycZhjS4SKNjbBsfH23N3KAbUZ
77oUE001tLXLcJiqX/wkQIQVz47WRdLl3jXEtKnB+4T5YNbawUK/ymJ2/J8VyN+QSPbjifwZGHCc
N22GBfyPKcmQI6tibrRNfh8P+uiwFq8hFjwIKajcuO3kcmT9J7OXNRdrvdZtCwrTkDbk3Mro16aP
MppM+apAn2o+h/dCvPCdd8o8wVwH1A6736C8gu6TM/j52dm2VTqswPP7D/936ixic2IPAUBVdGP1
LMFqHQ+HSzrItcB+JitRJ84ZgEWJUdakHqWjPYmvnqispOz4AB4VlRXAKgn8wB6ToAjynOpE7LNY
CfK5LmwVt2iH0RLUIzFnakk9Adma40ORcK80EJcHcPiXlzfSuEqmSMkFRadeSSc19c5NJNqDbame
ISnWe11mpeusZzhIpukC/ApWCAv9q6neQ9S8OhpOihhyCVyfowPjmBbZleTidx6el9ChtZxl4qph
eqoKMJxZ6myl6LuKpivXHu1ZSBXhblbffmXsheWH6qVHD2hCzygFnWmrq99AwswxSijh/pDIdqEq
IPEUcgzgF+vcXOgZEGGX4D/HX5VL4dwVfJChsk13+NUFcjNrDSUqVnkA1TJHqc7sJ3W93De/tKxl
N39JIoHFQUyYi/23mlH2hN6JuLwU7HqVMHZpcdtrTVivQLAGCC3kcHcnNs7XsGmfTlz4QdeznW8x
1KlSgaSazT0LgF1ax8XPOvJdUqACHciWAAMaEA4BI4HskEoUzZiBBnrnOCH4SzVw8V8XTRU+dtFx
RCyCBQlnol+WN1QUfp7ieqpLwurBn4fQr2zDttCW8d8rotMlQ0bwiWviHjV2yIcEZO7kfzfWqj8b
NAVaTnXfIbIOMzk/mtSf96ap4zb700KikaL1NM08TKS4cHd5hyMu9KuOOQYbzGRtyGb53azgfG1k
MFCbKQjN/1RdAkLhrrZTc99K0SveXYXDKMHjX2yvIys9KRr4CtUHkWSt8g/BOBoGeH8BusKac5CF
yC6mZ/0WNTwdwrCCgYERptimfsowCD5v0TmeRWccb5+w+IxhGDK3w3Y5a1TiValK/FLjiEddaNVk
9trwXH4EbT9yHt3qugeCtdtdGMaikGPUbd+EfEuWbXMiXqGVCZibqUd+/RMhjFTMXH593r77Anys
hdacHJnxLEFWAkSYS+ksdhWW/3U3KIfyR5uNkrNHiXRxb8oHzLejQAoIpITkK2Rm3O1mryByo1We
JAtf+xKLxwfUq3Vjeuh/2C0alzCeCkRWGl2IlPHoSkPjnmd8cSvWa+z2v3Oc8T1c12fQuVOMg8X+
g5fFAEj8fAGqR93aIb2iC6+xPlOs1T/oeaiaV1rdKNDWLZAYU8UMff54XTSIbAqSo8JTob1qQ0BI
P8Hj4lADrMoJL+OuAvrKOX/67t5ju4rf/K9p8Z+SMiO9e1m4eIlHlmOg3FjTvDeMC8VLTcZ0xYLn
WVc2UO63MRge2ud0FcWczwakNEnGvgxiYdaIN7mHqP1hFpEgK6jgy7uL54e5pZsJ+wN1jrq1fNHz
JIn717fVfE8/XhE+vD600YqqPH/Ga6S33/9tmQGQDILsNt7TfTI3ARdLdu0t+HHYraidl7pfGrO4
I8DX3PvHB3g8XetgJ6RerJf0AckNRVckdLrOeg8MtzaaQ/jqNRafad8AkNXZyPukKM1SI7S3JwBh
uU2SkYyaQZ/hYBQfc7c0xhQeuJN8ATnoTYQxKoKxb7+H+i3YmYFc1KaUH3M2tKtNzaAls8/RSvmQ
o0t637h+NxmVJ02FWVTsOtBRDn4NQXN26FQDfi6KIGLGzqUI5Ebsf4Cgc7LLPwKB7Dn/IgYsrbhy
0VFtt85M6mYyMAzLC7S+XtPtV7N2B36jdiAz41SnHDeVGyTEHGFDtiFxmVNI27Gxn6JeLLm/MCGb
ttQITOTfD7T+zhEMdivLQ0NEDqtLyxe2bYlzx6YlMlPSWNJTZd18HAA9TSGjzdWoTK1qYg6P+3cw
wTjYHwTfLYvVzDW21kqPqahMpWYZafSvabK1e+j0h75GxPGxFjySyqt0pfR0cR+yha+txD2HGuCw
wLXE8yWxHBEDgmtoff1GfeZ/lIDaPexQcFvo20PfE+EyhSgDxTacnqZ7mYfeC/0fcIR97Ot+mR1W
dbl1/Ta+S0S+FPYmRmRo13YOqXDf3eQkb7oMa2MHite3uhXNSoQuBhFVjPpb/sLGIPdZfRYXIBxB
OZVuqqwkIW9dJjMo3taMXpg4lH6+Us4IherrWTYk9fGPIugoHPvxA1pGVyD3DoY+hFKu4obQbWRX
dq3Z26iBxoUEWyvd9bLfOqsyifp4xP0oXDtpSy14qPG0OBNK2V76/+6SJutk+PhqyTIkcdL9pZ+t
hGFJLMYHiM+RlKJEG31X8M3WSEjGXfteRfzsoGO4VYeF1wK8x9ruzhlJeu1UfqEk0wXcjASakIIL
vKt4YM6bPE6MuyncXOyCFOweO/4Y3kYaXOTy2rbHuDWQu8JTyyC+n73SczU/xv+hTldOu/y4jTsV
nQ4K7uajEosHlKe4XIsRVJnFnHTvSwoqw6VSdOW//lWSiSetBno6HQF+P3qVumrci+DVucLwMDN2
knrqRTplm9AeGFAw3aMHNOTck1BNmJi3tDRdpdlAJ0B6QLwCRm7ZGPvV7KTxRBBvzlREmgAxcYBZ
IBXwUFeCG9i+Rgc7azud2AIi1r9oQzJRwNkVqzqXER3409Owh8nV0AbUyxGs/CfchcpZNHTxljop
SSDJQ3RhhVW0UNpyKKpmAx7fDierQ1ik+LunrfDPQFHVFYz4jj4VMfD07g6AC74C0C30jSHTEugc
RJimMcfuOJmtUjpGPluQrbwgzkik6NBuO3QoG3NpSkAzdA4mXpH8wu2aE1aDdFf4oPKWpF9QOif2
KrzoGjMlmSZ/ZnBiGJKNzHYm9ODuFlb+ykdMMjwqfzkSdYsyxpTD+w+sejH8Xqk7/MY9rea07Ifn
XT2H/lxSsy47oz4/ddUYxWl/FA2lgPwGhgPBVi0CZM76ZFgJo2WqTR0HU/yhD5nySKtVHci+8UKI
FhZav16wCk9qfEwnNF0H6eTCBfsU460SngyiEaijZfmT8bTGfpigPYfg1HTRZ7LgiiSTznaNPqZ2
OEOtWaP+1b2qQDFPhGWSzZaTOqUSiqfc9xRk7IcWfke5PTdPNzya+oEaUp/zTanyQLwaBTwd6iWv
tkXQL4LDNXBqNVmQHHjjuv1VfNADTRuJSOgk1reJJDMi1UR7wl1opFOtWxq3q9LalVctt6ft9meL
irBF4eBaxeCDJPx8y+ITy7CiqFEfwxyqZ3Rp6sLggcXiTAOV/wSm9nGl52OWeanvve4Mgu95U3Tc
0gFJ3tx2CGNrjNpG8M9rElNsGAgCYZBEItB8Quqm6UB6XnhjqT6ne+2OSYG9CptN9Hq3F2ASgkqI
8HJI7g3uU/sr25rzXAssDNoNeGn0wCmaobwV7cRPx4rfjjwb/uy2S/WnhVBx3fI7naJbdXlKAXdN
ZL5VZVz0pvIQky2REii78t5Qr3dXniuKvCJjcVwfEN3tNv7bO5SxjrnW2zQ0nEPeswLUUAM12Zhr
q9rWYfo9i7uQsCiZ7/KKlwB4/AGGNaPy7dybZaiVsRPz5gDFPLepjYHIYmRkA8RK1NuSUSfLEf+6
C9UoHb9FobqdknHcHMuoweP5PHa5xaXDpE3skD7zVOyH4Z5bGIZVudLstoLyCSiNGHWnc45s6v6O
eBqyP926FJVbKp9vm1Fg/Ufm8HFybZiixNalxPmR82dp9GLWNnxYpaiL3AeD+Ks8L0elKa9bLIz1
0VEYx9ryw+9UWAqZsg+jIafJnDemoV7NdKqpGRILKjADdoYUqWjloa5xPXPo/b1JykcuOHcvzjuR
ku8af1P8WwxmNPoVnWy0VorzkYRZbYqXCtWFaVwHI48aqKwKxef+fWjJGLtT6NLd12M8NHN4dV3G
QHsbDG2YeOMTADrd98x6F2PGD6ozZ7JhxufacmyNXhfM11E3PajS8gPFKTHXxXpVzqRU0zY/hfGp
qGJ1TEI9FjdO7x5ulqU7WiBd3emZZJHEDoO6SCNZQJLqZR7HtTotq8hYMvlAe8a+0I6/aP+Itt8k
U1RTGHRCfW2WX8cCu1l42/iF2K+bzw1l4YD9ECu7ODsstJ2JAKqBCugrvCTOmMGDpqvrK3Qfrr8M
onf4okj+jDXtSNsi+1OzCslOoWhCu1H19XZtXB036un1zlaPOsjl23gaRZSCTc5KuwsRhLWNlqfz
Lb/Qznn0QsbthbUQs8HiVTqmYQqO62zDHpODHEIIpO1HyOfu7K+P6t84whELLQ60M39RP3XVmU0o
SMkptQiYJ+N0KnJX2Tmfn/c7MPDu09GTCHAgpFpVveUl3gh7pppT0An959NOb3sYsh8aWG4hQMZv
jgzj8CU6hZPSz0Ef/twp5Guk9YakwgwZVSdVkR0M7lvvO/+X4+glM3d+Bk/ELXFG8kWVTm/jylx5
hlRAjvEOCS99xs/pmBEsrpopBMYhSSAAQq4jG5R6+d3JCKXhVMOd9LQT9YoWglmLy3jBA8Bb5Ygn
OJG1mJZjbqzU1j/nsSa3ZeXFG8utkeQ52ASJmJF2fqhgeLnnhOYt56OqicC2kHaNRU6B+ovpSIK2
bKI99ek7Z9Ekty0Y1La2e0pAqkmSrWggJK+mTRD5Fp8N7HlSbp7F5BJMP9SnenPUDrabBYErcSJA
uqyHo0aS29wXUg0IEdkR85yXDwr3cN/h2pz852j1OArXJI8MlohEgDKq18jolcbHEenIddtixeAg
W8KEJIWV6Ivm1VGndhuvN/BVPddZNtDjr/4oUTsdFRv0nl8F8lSiZ616NOw6eWItOcGpfzEBFLaJ
Yl8Tx3jf9j3XfQ0AuaQjEnvOXgeyWjswnJsaPLoPHglTKs0FSw7DvFsNQNUp08jiiZb2lSlHPkat
IOAQeb9+2+qejDIdAOIEJo7z9w4NL2zN/n/yWKl0BECrVCNoJVeb9Sec2epdJFIi+I48ZlUVLSu6
BjA6YSLGzGJI9w500BTfP0jIXBCI6RqmV+0VyZol9JHFtht5eaNzTYeKLlWoxum+PvRakCve1PkA
Ux0SDDTv3zRg4/t1COj0wDRi/zPTfhcxqnJ8IpbhrlswvpjI89JolF6PHAu4FERK36TIVZtBD8YG
M39OD3/4CYXOjAQsdao1jTuZvHd0NJJFudh4RQi6rWo1EOQTDHSvHoXZkl0HWQ+bS1uTIiB/8ceB
/XXFe4Z+KzCLacEVg6/L90GT8phEa7C4c/ostHgN1w2oFxVFryICmloy9l5tdXNZDcZDsu1rEJBZ
7t1Cy7sY6caPegcu8Iu+PqL0h+tcQT8T4FwGFnK3V6GaljGMp99zxl3x+tZ3iWd4vagEfieRKBgD
IM86W8TYHgkDEpNuHpCaC5mWFCj7P9w9jsX/G+OoAL9q/DkdBI30JDlufbRHop/YfX04Ry2oRw9T
jZv05zScqbF9JCEWOOea9YICNYoWwXz+vyEcyQcvtDP+/ZVWKLAgzX7HQTW8vADU91mWuS3Qj97z
76HO8fzzwGjOrtV2LiHK/lL6n6SOVGfdtusf4lnKuJfCTRA9+ap5Uu4RSc03qfXU4uYL5sFoSmj8
MnfilhwplGfdsJBfR62OywqNkDTesrKEZC0LrSaBx65sOQWmJwRuGApDYA+eiWMeinVSVIK96HcO
7ARYwXIQsXxK87bHOtbZKqi+O+UnTzF/3g7BA3ibzy2TDnSMnk85l8EzRoK+0UosPMMT6o//lL90
RQYYnHIGRjsht8EVLe5Q7DD4c2MEW72BPk4PaHiLpvu29F5u0Y9O81vdLW0lIB2d6KvUIvp+XXdp
QFENe0n8SzAOPBmrhym+admPwx1v5WXNyr3+Ogqk1o4zBrgmf9WZwPYqe8yVxvcDFftVhQniMM+o
+AzkhetuGFVWeTTp7lor1tQ4LCcR4I/uQwaBsAeHYorNXzdQF726rQUZqyY8VkSyVkiraV+e6KjJ
JR5w2haU/Xd5LJVYZgIQTZT8kK2s2kU0tBCrFHHLLFC9hBWymmu1Pq+vEEkLcUAEMDAY2K0Kbh3Q
2c6qOdayfBacXdtEloQp9TTHya7XII7ga2gxKbqD3tEUIwp7RKta/0/o58cberKDQJSq1eVstQGH
EPCjO+fGaRahXpf4KbYBgtBdDuD3VFw7v2U7niAKTbhACq+L/0mGXDoXtCvDqLhbpaOkNUDD3tOy
AqnyW75TjFoGaE/ZSNwVEMmorsNxU8Jc7eWh45wXDvyiljxE2U6GS4Ca6huJ1Ex7IGi1H7hIr846
XGSUapGnfvAtNButSlnomNgK6Sjezv2Id4uycp88pbIsJBerrCu+xDTskZiuVkdRoflXnK5UFYEf
sdljRelVe6o78h71yZNipo2I1WeQKRITOxSbXeE7eU+OccCTFg8lsdxifYk1bBDWRDpdvaJ1s1xm
4/FhvTLyXWESyIfkp35EbNWuQ4bxQpJGchnZkXpFoqjDS6/7Fwz1Q0D4fOvG/tutN5HnHAnICUJI
U7JjF1FYB1lsCsXcTBGyWetJayNF8/yzZMQrF3QnSc9IiG1HuYkplUSJMbudtN2eymeXZsJDmm5G
lzQqp6k42mAz9ko7sdiw5LUhHpMnpxGBW2q0WZTKg8AJ58oTkGPWidpj7Mwz63FeHbxhLhIGAwGk
8PKPkZQQlsIYNEohYzuObusPIV2D6nI6uYTDAtwKF6fiNIMnJXDC1M0/7ITIDWwY8g5o6XEs1ONv
ERBrUYecEb67YmXr2tKz8ov9y+6ZV6jlJNfxTSvUXBxuZA0e7YNewVBk7TBctdH2z7uwHN64YMMF
MyUiJ5F03p8gBsS7hp1scDxIMGck2BCn0TjZBwB1+lPi4xJTpUW+3bnefhWj15nXM5O5hxPTbcGF
v0P7p8bLhrtICWYN1E9Gd5DyG6vuXjpVGJ/nnEBAlKHmyRqF7itquNIRTT/eaLcY7UKNPRwi0WJS
hmqDj+ybNFdpQ1BkisWL0I9CnLSAbDnQFgpOv2DYeG39/x8ozLQ0il8DdCjVE2hxx5a0S+C+Fj2/
mTSRSvjPpdRS2YX+WT2Ho3cmoYe5fsidjByga8/hemg6CmKZCuE/lywALA41marJ1iAzV1ECHcni
yf0bH8HfB7GHei9E0Gz7GOj5RSFiwSEI1+K9nCHYW60Ph2y/vPvl2B0gqMcRg/WXapvElKdG/YJT
dk+07IYfYjFNvXkIwxudUf6XreLBgGtPDcB0MdTInYYx6ny58We/AMYhhooE5VT46CDRV7YFmiyN
Pp6c0y/4/sj9NFo6Q+MzoD0AivvRBAUdS6ux56bUoaCsj2ATJW2QXx8e/ITDJ1oX6KC0Cj0uwPdE
fLbPoI3kdRFj0xBQ2c7iWIW4qG4JokXJ3tvP9geeFjzS+OmviRllO7MZdCl3+Qbvu/TwWcL+M0uO
FSTR3iCXh7DKIVeFmPfMREqfxDAt/sHK/E5NgCBceQLiG9rkZSxwCBsZWnAYfp+MJ5fWFbwc2LBQ
pIgTQSJjeny3Gj3jwWVOKqnsJPkg84mYpedDujAYszECSLLiHBbMho2GWi3wIJtWCNWdheaplpCx
tULPqIMWQ7QQrg1nuUu6MCkWMiiqRy80nnT8YirbrhVV1avkkQmodxRvQW9Ap1J/qav89yKmqP14
U34GEDvJ7mbnIf7o60tvv/7SHJKAA+pHQat1OQbpDbtVAUepS68cYaTyDziYJUAYY9t9yy2fl6ln
XsDRsm7lSlHesES1wlVhsv/yaK9InRF05b1pP07kTl50IzN3SY9TSGWIeVvW0c5jciUTQY17R7CO
nP86uINKWPakjfUbU3tFmyYxDfK/02jeyhawu1CtirEeHoeFanooyR9iByotnUXniwNT5XWQi6fR
4JL3QC+C9v24xjR5eHTEOOwsS2U0n4hB/42F/h3+bI7I+QRMXY0kqzMgMrt5XKnnITpWdvbCkwjt
Mkb0z1dSrQSJQ1zZlNKzBFl0cszBM9TzzHuqb5dfVcqtqyYNRb2vbz8WGX1ttVBOpG4bU4gaSBCR
sndsY6uiCWYiehGTN50pjd8VCsbGHdarJ60Wjkvo0f4+bzqVrPXSlEPqMi2vjXfUPVdMagu/oobG
pNzYFniNv4I2imN0veo+gtn3Uw0Or2n7FKqW4nDAsZySipUB2F08hVQtHxw1+I9J/E/XLWORHpBq
noNeEbW/ZFC0U5aoSTtCvJfq/Ls2V4Ral0V0BqtpfuLKos0Z67tMG6ugYjAT7Dg6ezAPW3F08mTA
QAYZ0uk4B6hpAP+x0dYLDkkGHA+Ig3Rdjzj4xEMlajn7t5opfwr9SzK8LibTuhNoI/+0s+H9E0U2
mgxdiclzBB+bCH/8D35L44SgPaD/mw7SWvsekg1uQD7nUYK2ufgX0MlaNxnXTL7EJ8ENTAdlDkJ7
l86nx4/Ac0rGhvXItX2+pryxF6ThZXywmViexFSWmwS9ZWWXxMVWT7D3vRFtz+3C/6oE6sPxUfyS
dAYjcZQ7V5O+mb4TnDwTs4ZOqwZre45507/7yZmZY4ClMZO5dVqkIErD37DC31jTjqI0SPWQo4h2
JTt/AiqRXo2cow4oKzXqbcH84bS61Hdf0N4Unnw0vbuQ7hUTCEQBDzP/EMc00uFigCbySLvyagdR
UrdOfhlkaQjsgq9pKYgPbm+dWXHO6Zsz91X7Gy5WHJJ0+rgj+ctc2MMi/xvbCZJM7soWo4D9TqQd
zwxcX9pBLTfLIGD3YBElOrrBg7jSVS2I9vbOBAoRRICCGK3Fg6UqxfIDJiZljJ/1lCk6APUGUsib
Z5tZykYTu3kZamMvBzUONDPAktxKnbq19mH9pBwZ6fb7cH8lTnDYXz/gvxqq7QV1ZCrFWmTFhq2J
TI1QZoIvvuzVIu4xCR+eOJbhpZWAzDKLQorYpcUGCSygWiyEstVEqGTicmT8i58vpimdy01hoOLa
ZIssUgox8DyVaAI+tQn+Cx0t/gv1NUWqJPthOY8fxGGCuEcX303FJrZog+f2dvL9bnb6fvk6EKVm
YyB5sUvgPrenzmtO/YEZt9ajXklsvR3ZnSredWI8FfCDQ4W1YH01QR0XQ3EZuz5K28q9nCI67Daf
5B4tkVTapMmxY9x+KFfUlcKjNG+eAt2KTE3MRIFxQKQ6U1qs1idiTZFqZF+xNikap7HcBhY/oYN9
z9DR9L+BoQMzhY3ncrSFV+LivCYTgBgzEXroKcwRQ5MHNssZJwQgLmE2NCNnfrTsPzPnir8fwdHn
p6nfafZMsUtdbMfQEJ1e8STu9NmW/UEgrnHS78erje9PGw0gpTpOx3wf2vSjp+6xrywcMxK5UBMp
PLL6wABgJr8wRQMwW1Lb+Bc5nCwYCyDGG+6/FBWqHCc9AdYkeXV/I0Q4sniNlRKxPFjU2dsO9AMz
c84GpEcsJPTSUHMXJpZkcemi7o59TpwAdjKRKd4lo6h+zff8AxEs923b2G+PtTNzm8WPSPiFqppp
QArciZfsPrFg/DNx0JaO7dncelHQR/hffoQ5DvzPlABO15aDt2Y+JYjYoHljLyItgnqG3FUg8lVa
1gwk5VrbQlLJBsivhkvcoghh0xj1bkrqZk85TZrQ9fWn9TsUQUVxMchOKGYbfUCnIDvRnwZkBP0R
cU1ivNkbbjG+ySFiZsXR2oxqkMyJ7hRUFINARXr3w8Caf8iHP0lvTJQno441slxB2UZ+Gj4PmyeD
63K7lLmHX+PxpHJ9HdyXhbWdU6aRP97r0CAeT6ayVklMGptMbqQvLtmsy4eZ1+aLSM6RufJgPLXe
cDXI2lucY0lcl6ynlPzAgcpP3GHgrFvlAIR3pFd3B8zvf0b93BqQubmni+uc2tCLb7DuVopaHV+z
7mBfWlZRsLSRqPAp9buKHvD8A+XyyNPtLuO1kxX3ksrR4YyMLUY0pNysf6XbHijjKAp3cvH82RnG
pur2HuqFE6TecIJyW9DCcxqqqcuZmtgi2UpWYmiNn0+oHA72Uo4Fza6hil7ipZjm8TuJaWo+6yW9
Vp97GKEyFTGJb3D+E/fIuVTMdEoIEt34+oeKfP48qCk5+n4l81gc8Jn+uqMufHu5bGxjUTGCnvVk
ofS4YigtTrjEUgK/FynW9d2rNs+rbz9H4d6gIfaqlXZrd3oiuOc7Q4xdFMbwP0cSnWZHUZvHKWbC
eyG+GefWE6Huy3YmvWKimvlNCuL3b/bCY58AW2GZ0baFOjkMZ80x9a0kLlhzNCXRA9tAbT0oa5Cv
fsGe253uR30Vnu5KlapcT3qG6rTHZx4v/VIxZivzl+HUiQqRo1qY99BNrbnLRyBeH18OeOmmQG2K
+7VrJWUBmC1mL6xpu51qUWJVG7Y/uyy7WVI9VLUz2XaNCwuUqMAylGqLZ6AJB7r58HefvE/FCj4D
543AGXgMD/N1gE1wmwTlzBilHgjhqMwxrt+UUBJ3ECzDPObFRI0S+0bHDX7rO4ZwO+QUucvvpvYP
4X/qqiIigewyFsO0zuG6pFxA12tqnHKYdMEodIdQcSxFW1alIQZS72SNefHHedPY4XmCn/HuS02+
2nzfRMpZ3i+G5VoMcG8bOqq0wD7Wltw1q4B+C+uGDAKikv76zdDRKylaDBNecjr2ZOxUL4q+tcAn
Q4mkqjWMXlA47+9QpBPDJYZVfeoMidIMLdi2sLzCQjHKXrD6TuJEzxbvJrOHCtpQh636sPlsgoFr
2Bmm9UufTqwSLnDKeR3CPhVKD24N+Jp9GIBqhStGCfJ4i2Sr/2InfQh7QiPO5Gez0uii8BeF5c64
ZrmHiH69YF1vPh0rh1r4CJave74raQqjuJs2avbbZ/TSVgHXQyNfsHe9RWT88jIxyC+3JmHSxbL0
IoO3/Eez/3u1slFQCQ8bK392Ys86toBihWfmt/MES+GAHJ36FYmRlxB85Wd76jGJ/5dsIFepUpVR
g6W2PJ1LRWsCM6Gi/X4vEVQv8wyFeRIJHj613TvsakDXhgqXTrWWKtl4fO9WUnO5KkydCb9oGK2E
LPtwWnrs9GECgFPNKwBffnQ01px0lP6MTT7Vpt0l2xJfDFypNdFZvU+Zeg4oMdjoZIVA4m5DN9lB
WVHjpFgH200XSbRFOkZtAFBbyA2ag/cPYi0AphaI1dEz3NA2Dhm9RCvaZtiGmflz82xcgg7F60FH
YKj1JGmXNZ3nPyiFFord5H6XoHyEv6NHEePNy9mHlJDR33/AgCJt5sz0mA0m94j7A4hHoZgEA+Nd
W5Kk4AT67cvDhAzOxCSBWGMe/VGT4i1mlbRIUfTkwgZlREZj43Dz11urnDV7dlrZEY5Xu7I6b4M0
TW9bcDZEM7f+jm0VFAQiWgcRFvK468Mq+qFDuySJ1THvDlzQdHdnTqOAT4dHQWfb8AuKB7mVP0II
pE6MYlHYq0kCuObNBoU3IcDnH3jh724Kayc/Bt+NZUFDWLJvjfdYonmxiDP1pVBaUGG7kQ4u2KIY
56QsY7O/2dMa7xwVDPTwH4ui8w4N8Gmz2uKG/33qBVDKfOghM1Mz0xSz1krCG3zHtnXHe/4T85He
nMtSu+ma4+icmKDo2kl9s2BkjqT4OWC4uUuSnMk5Q2wBtznIHp1QUfk5YgkYeY44NnkPTyQSEQCr
zvl83GT++VniimMYHNKrzWFwX0adLnbO1zJsxVgSJu4k7rxCk2Mnq/2BF5pt69aZK1S3eWHlA7sc
dpyiNeQlKrTUXaW2lV1QvijBusS2I6deJg3/K/gaY7sNVqhOWI6GO97oRCRcuP2Qrw+1jMyCdnPw
vpiLfoXULJh/hALylFsfnHGO9Vo1C73rYPiMplgAySfZfMvuD02aBVhX6GgbRkLnVy7MnNiwvC5W
Po5+IOloGZi/RL2snZ65SYWu/L9VNCmU1t2n8t26lYpxJJPjwBurQAmsE8ZD8SJ446upOI/Rkrct
ccR9k+fqoBnzjpmvYKujTKS8YNq8XbsbKnnscNbfCsxSW5SQJ2s0kaTl7IkTkoFFKqLFKFRkWYVQ
5tlzbMge4Rs2wLfS0AzXmsBFFic8OzDjNI9UwRwpb5AX1e1HVDYiZWt/RbtiVekcbQrBnkmNtymE
mNGSfn0NoIOPlYEDTRYCZm5FAauWqowFagpt34S14y7pgoGRhRMdz6LKsO8mxq6H6FzMYYfziq1u
RYGmExrsgmoSDepBWpcWFwqblXvT/wFyHIkU/h5UfkX0gCM6iEdp8TXua1bI+ioH/PojkgO1yhE4
Z30W40RWDhZO10EvnLvE+WpWTWhjHZ3lnQF/eCQ1bva/LSSoILP1UYqw8DV//7xMs8QLnMzNSXU1
0YV6FPVvVmkJjwoTNyZtVnryXXj4CALPMFw18J0/LQVKA459g16IT20/msFren+omN3BJSCaHoH/
MjBLlIkScZ0sy4d3K/Kg7AlIcRDhVmZuUK2VGbEwsfxsz0F8TT/MOlcb8HmjZfBl5PZ0NLNMKOlr
rhj8591mQIu9Bk+gAZud6pPkJxqKtlQk/grLj5RMTYv5MaBsS07qFv5ANGDmcm37rzppALj0HfWj
DQq2Dach+7juK046ikA9GBpikbkHRQQ7W4jlE120AxSbE7R0pIL/0KXlZYcrnzf9K/o0KcirhcZR
M0UgALtKzomqQhK01QprxAT0F9oaXEX1hXn8SXQrZEgjB3BPUVTr5LYaVZnt/0O3Rv2hlXE4BJmS
rxxKNBM8Ztn2gXMag/rvObaNx0Tuf06wXYxcQOIfiNv/cudMTU2UTxzcucRTqO0KLFusu1PNeneS
uOlz3QPG4O8EKBxtDTus8fNHRh+lwTfgfeE5FJ3rZwna1U08EHNC22INKqRFHQoUqHmQZfRqo12b
JNudQO3w8kfNnGI3Ogvr9ruHF1GImz9/mhpBa7b9ehHtcHRzOHgHfiVaRxBzJlwS/u9jXgq3L94/
Hr5t/CwwIV++eTJh3NFws1EyuyYD6Za/dwB5aRbDSbRbPpcKdrZ3DG25Ug6S2bNX4LXvC3nk8gmT
0vFaW88Lp3CUGCQuGZE+RDKifjB7U1DxstwKR2v0WOOrpKD7dGE+5uw8ueQ4QS+Dh6qxkHNbtxi/
OBcOrCJW4FbrF9iJ7lyAYNBRljyR4UJmpv61h5jdlotxFGb8Kvbbln4dqT8CQz3UwDbfYVoPc/Iq
HeZBMQ1Uzgz+PQ9MxXf/J56gbu1wvyJvgspiec0eTNwnG1rj3353S3IQmHxilgUBp0oxdmpd73cs
tsspYTGQahFFX9QCE+fNIrjDeLlLvTVNvkxgPcy9IAVvyi/PH/Fxd7+ucA7BXt6iIU6JeRwAInf6
bo8iNJJgEmJESCFDx1U2az/6qnaGqEXIJo3s1EtPR64FH6OpiBgMaxP/39kyjrP5cIbQJVlSvLtx
qblstrW3XQahmvJVGHhN41z1BSwz8OtQCcDJIaMuxzQeHkmERW3hTc9ROw2ty1JgRq/bMndTOwKQ
+sockmpgphHARO9GVrMo6sSdsHGiNjQ3flHAEi20gl0njHBmTCtp+hhWYjAbZcGkfvv42KB2EQeD
NOGUh6VSfe0Kc+p58CVmdxUS4HgjKLSdy+2Ca74DaoqMw/4uYAtOCuPgYYN3M5C/q+ODoHi1dNFE
HliPIQYoDxaf+7Os3ROIm6Z89ORHJ5YuBGAaXIyu57yrK4Q12k28gClOPnoHKnQtrItxSZcXDpnV
UV3TgWukG5QIAIRFRPVNe2vT13uoG88fuS+lxIi9N+urVIuaetlruSGrYqTQAHZO5GFvrXZXjP/n
Y8TF6tQ5PhDVdPHb1AOQfloOY1s8yGxFuYTkjyHf/Y4+2CKCcsRuQQKi+rBe31Ig2rro6UbS9YaJ
T/yhJiwpvDve/ShuFMMxYLafSNBiP4E5CuAQyWLGcAis+bJ5E2PAXa3TQiPmPKFgXD9LiBuSN7JG
NZlhwq9ZTmLj8rC8jO5Tejx2WCIMGx8Rilq7yaytB7s/hpNNSDpL2qhKDmIJ8ygUheqcz15nG26W
2qj6YRhxo9kg3tvLv6673F3MqH6HA0Z5KlIKotmUXb5GgB9UlvK9ZQjFYwMUlN+Id3ttGt+oYh2W
WVTgrDn8rbfMBEAOdn+e6gINtV9U8XJNBD/4xiHadj+Oh4CgoG/4s2SQjaFfxEPaht3IY0h+blYo
fFYQ09af91jwUBRAcq6YhxOTK6j46T9gQaZNXuryY5yzZpos0joIpKBSEduraD6Itkp+yE5N5Zpf
yQyqyL8yzFWSFTjN3yZJwEEi5cCcirTSdWpMiMgw0nZ/jzXnsRn9YkWYhJz199b9glepgGbFErsh
m5U9UhSIDX3k6fNyfPZHGQRPVKet+0q1zHa2X5Dm4LiP1jsxTnxFzy0p2FcS1CCtYQmnZBmPQV1V
V62hR4iyOjziv6MNoKwhvdmIGQostPQFToOv4muK9q7AINKHi6QzJEWbgpVSzKz/wuI2dYvxsbe+
ydKLjURl+heFRy9QyJPZ6RZVo4fGd8SuUod3A74Jvit0Ab3buY1TyRlOAHBEFp7Io7el2OuU+0TQ
pWiDqfdQ89QPaqYfDd7Crc22x4nRo1ldna/P4ZgsGAE3umZ72bZc5IvT5/nZAYZPYG03Rpn1cDpT
0rAiDZ3vSyp1fHLLPqunxzayTGYORF8wboMh5gzuPxbOxZSzVd9o1zuQ7oNciLuXDNGfoSOExiGa
A2iG1qAJFXtzNepavX/XW7RqTf/sDPIA2Q0TZk+wsHQ4odGrDn3t3n5Tj+cBptBZ9ZLZJX253UHw
+H1AHiImURUJEJWHi3ztvFK3xThVMiX6qHSiY/qabLxxpIFE8di+LpDK5kx2YHzUge0bT9t9XDaj
MIQ7ojaasu9IvKgGiynHllmdkUC8evNJ3kHjFDUd8TxcmrchvM+4oUd51kIc8zsNjRH3PbhHueGy
KD0g1eINwJkcHFtFMcLSj93wNT7gH0qlLX8tZ6BoVbJxYVzY9QL8o84AoZBNCQlWRxBJSS48/Vv7
DRIcp3jtAIqAWG7L1c6YL1z9/nPWzacwuQZP0AwG1slUzLijFTWF7/5o8hnPvszMqye0t0wmO0i7
hA2x3LNtL6NHv6l7CxALKraYnASo8uG/mFHmjH//fxufetTnze0kOtCaOKQK9Ux8zbsw/I3/Mjt5
YRcD7vbguKxy5j1xpEoUT6zv6KQBJfoa/6TYQG0fWQmCINlqMNj28ZoYcApwcbPOwaQZYL+qatSs
ponTWQdJfSK45at4OquAcH5Wi9MBNctzvXGa+uGJCuvijastYgOO2JM1mwrTd+z9xHbPH5391klD
BgzGGyFsrfA6OKNToWs4YuXbBjsXBbxW/nFOk4LprC9kgu7bTZmQ6QvjM0+0Bp/aTsv89tMTBVZG
fu/DxhYbI1+LELmTli7Yaa4RJiFYRPjOgoDcM2OxUq1TK+Tv3iwsnCL8nvmEXY7UE0bSXtwyGIzt
BMwM0BEiX6uhcSuAqT0+qZ553xa3nbS+YUpxsexXqaUNpKAqQzGDpfnxEvudPTnc1v1wLSu0ij2Y
UdZPfujU0GtC7b/1rd4eHDIX+4sfQ2UMlaMi4kIMw9FGglMjmcBrudtQ0BDoEkRdNTtnk1j5nLbc
kv1FZsEqzu4qPZpyOltA31A152lktroJSVRmOfWIIW0VCKBp/6/UYJRybUpA+1UcMulqJSsa9SZl
jjpxbAYpEEVPYFasqYcnkHat0eMdgFzU4FAj0uWwkyUyeSyB0Nmnmb2XLIg3Nezxu2nqhEh5tVsG
5GVPU35Q3XmVjQKBMiO4sZNXR9VGY0h1j/RC0QDRy898O3lGoG+SNDHfpJrK/MqlNFJIwsrABX8h
9hOe5h3QL6phQh6lNbH3TRI+hEXsUikILDj/RiwJWEFMm5HzIGfK1JrdpXUYH6cfrmuRVZK69XF2
pQXu5okSqpt/sVNp5P8mS7vumN+0zQw+y0ZZM9/Y4Ap/BUPY5vGI2AMun/R/lyXolKtui7uMN9/v
UMYVfUkG4gUyCas0mKXGv+xeKpbqm/iMS3BPbPT8AZchENgX4NdNGfxlEdhcwqTwnCeDh+MYXrYd
HXR1UA6PwYhxVQo3VSamVTnwthsNwVQG1i0HZdQpv+xGG15J1PTxAJ5a/u/AEZMOgLVChCuB9e3D
m1rvRBMXUcUHXMwqExze3HMECMtZpHuVv/41A5h4BUBd7o/gl2TMOFNMVJHz8gdtSpR6WnV8NULI
l4m7noop0pTDuWxvT3TL2XZ3EeWt7yz3UqstT3t/C04Nvu7gF0bhMvqCHZD/QWjma6ccsYOFAkYK
z33TmJFz1CHRVJ7EyG8VIMexQHqfGWpQK+VDUJHvcRJIxTC/fTLGF6TbGoKImvyt88JfEh7sYTHC
iLooqC/RqiCSGvLIw9SWnwO0sUOy/ldCbWF5MvEJvpM3kWnx9DwjvnFqMsNYMe5Ekx4wDuc+eNb9
5s8q4KlHQWxPjXwtEsyZxTsiH2jr7oZLNO5xJHO1sSkEdq5T9AJwMg2CN0o1RW0lTOLAD179EAXr
YQ8GCjBcorkDHEFya6tEznLJaokZtba+PTE0JQsNWgkOFbJMilEYwhgq3SJCu3aRMhxVoC6OJKTJ
5D29lh8RlX+ogNEn081+vKPYBA7CBwwngNmk5rLzY4mdk4sMT54AbXqeg3AoyZDyzDvu0O8thk2t
gLNrwq7nrRnqNSTbr9/LQmiN6IRMw8dSiIiM+CPJzQa07Z4HjvWpsZwESHVxyp1D1WqOHzFJ4seU
xLrq4D6Z/HCPBAloyVujA/5+yyzQI1YPYNjJkQls3b7ecKLSb0TywQ1rPjT7AJnAyotTXMJ1rX04
zrXAxcoroCyxdL19KOHZzFI/RsMkRpJ6G6zV60jQlprmZpymMDjcNT1a+pfAwC2ijfB81RJkOWE6
1wk1N/G8ZiI0rpNuBsEuuqKzZs/noilJVpfRWB4UCVikU8ObYE0eMSJhoYZAC73PRUtvTFz+e3cA
fLeAnyTXVUxhjs/ywTMh5t8OrUMshIqV4bOt2lYQpPamI0mCpgqn/+BMzGgZUQUYVWPtZgXiy/AW
zhWUUrtNYT8xoJe8H+7nitfnW/s38YeVFx84xlWWHSa850MopKECUwAhPwmuXYo9cDaYdga5w/SR
82VR0EQdIeyG9sJP3p+dWFxgJLVNWDHh7LbwhmZZ79tv35RbvSLpi0qmcommF6w3ARq5srYTENU5
J6dOqk4ZAJ8n5CxZ1jJjfLPB4aluoNOGyOYXBjj1p0DxxPXXsg3oomP3Bo9ASMozSsq2iCvx3/wd
TxuARJkh5E0J1JwKpYOKsoZbU/X7IwIYXOb/WYNkft3cmJFkGjIzWL5FGknsuNKDDqfoIgBTdLyt
oRUcsKUKFXEcR5qxTZZEdg5EihsqOpGrKmKsXvh6G0BR7j9MrflOVanPG/YabwPL6VX9VbViH545
uBvsA2ORTxhRTihNehMEfU74okwLXj99WFltF6zNe0IHsl24q+yyNC4hwcZx9t5XRWY5C3P5baGP
HzAzFrB27VXe9TmCbrbXH81Q+Qxj7vgWAIHfkVbFdFjJRYOYJqwaFSIwd98Pfs/WvFRopFNN7o1z
PLCFTb445yQu185dYFr/HsNAxI9nZbMZy8yTcL7DNSm+hSk/hfspeUcoq7EI6zGZxGg6k6XxOnyn
qCZ+YDTfUzlNd+hUD7q4xmFFb0O2nRTmsYZR18XHoAXTAu28LkZYVrQOaepveR6f6rBPvYPNU5ux
HPoZcVz4vxNOelILg+KwjhUCxGNB2qwyGkF0wAi5C7+FxfUqrEBsM25jkJd5/OiDeAKJ8rkqWqC/
G5UO7sbeR7ix77pZUq3oJZrdMvDm2Vb55lVc2RIUC9870BTZyG66LAux9u6XpGIQZQsq62N+KzKQ
fqbb3xTN7X+hNFfLw0XHIyVXxZkrz//pbtKd5lYo47DVrXwX3TmzmBPI46wNPb0Drp+0hP4cjNbb
Lvh1pCpEONa48SByOT+E/hzdA4B2fm5WEWALBFDlU/nP1bn1xk2BoW6+FB7WFEseiEd4jKvR2+sT
9eFkm+e8FxfYSkrorubFJRVUQHKhHFJMJl62pDWU4ai7DX+XrxlvJGkLTDm7VBNqS/G9WxJKGVkK
5aHGCyLakCCZXzK/yGaJF4e7KoRmQ7esPw5/qyXeMoUkrlG3HxgM/p4NC/V6/gGkY+Gna5eb8vc8
VjXEHATHiw2WhGH9M6+kOGg1ocWgZUkbHLyZwHhUIl7kUJqYQTmiyGMLEuwXzzXY3shPcev4ZgWR
ytpCCWjrvDwH1rGBmcdBPQ+oTIsgUfZL15ihYGzMFX2bC66K1OtQLYMzVe3FmLOHP3UbPDStPbXd
3oYpqb1fMqRvJeID/KOYNfm3K0o4Ad1D3uROx11J4OXRxpFao4pQLxjBnC9iQ8Yc83i1p1BW35vV
Oa46999WswZAsKtQZ1vN3qMcagwxFfcIwMv37kxOHw9KeITOMSnbrSP9YI3E3HeXqm/rETn46DtK
in8FynHzFnheZj5kaZC8WzsbWqSQyYwLk8HBqkLF98sR0cGwORkeH90am47QY0YAiMZN94me+pCc
IYSlzpY6aHvadAtHG3uuqti3iy1LyAe3NhB5z7Q5xxY4TQPDrI7SQsRT+BCoUfnAXKrHm1zLqZvO
iCZUj0w/eVOxyIH3vMSLxkaw00H9TkC+uiLsI718hpcdaCLnaeHlOwPcOQm+UO297gsCEK38bUx5
peBbXzncPH7rybdEUyDooFMsEBKOepBF4gA+JFd5FJM4bRrZ8pSCWo/pzJo7qQO5qRCCWeQTlSZ0
FfE4HtJUqlJFjywl9mSDdhIyU+OzoRuUNyNceoXLnxEcnCU3Ir5K6hoKCfMbIW+2aai/9FwWfa0h
LnbUSMhRPhlvbFT5Hv7iurz7KZ9DeCyQJB8IzCkYE8f7GdzZpVpnF+EbB7vcVOxe3+iCbYEyQtil
A+zTHZCpV8yWfBFgobcZkc5/HrYBGI1BcsCcxDBq4az0i2iNsdCunzm7JL01xvtipZw9QExKkUsv
14fK6GnbXmKYaMWV3RMUQMKn49uAbJL2fb0qf6aMxnuPy0LFce0gYQxNobfdwxKLhJuqmpYdyNpn
n3AesiSoFLVKn3GP2oNmR6QcnyAGpNiXSy6Naf4faNuuxawutID9dZ1wYp/L59rdrNGymrstRO9K
XEvOuRILwVZ57ZDOH574DNmUjv5Ig3W2OMJORkdHudvsWORT1gB0JZqn1vIJqfNVfvCb+dua2c5g
6tULDKC4h3TkMdBlRxdmitSZgllaUgdGqyqIfd/7GUHAn1sVcTedFQGywWRg1DWufxY3xR7vm6s4
1n6o1djaletbqSjIpDVJR9OVZBHuvB52QomryAyKbLRL3CETq+tUBeG+p7ZLJbdR8pSLAONJKJDm
bP3HEvX0puZbd1GIQsARnhPyRc40/Zp5LSOqFN8bYmY6fNvDdFrnItVVAXEbvskooVsELl3lUHER
i3kvz7n7VrXTKWN0RH9dEXu+peb23b2Ys/FDmPFb+7x/ztGmTeZx+yg4oWZ4fphTKEMtWOqlEePz
t6rY2xVISPHbQx97gzfmVmZXputZH2GcsZKVAXTGfchaIGyn9hgVqQt+3ZAP9uxvhd9rOILNQzbG
U33K8SyItzO7HIttBJ+1Qe2UVzJlx++vMD3sduweUUEXkGbSVSBxx0QJ6AnZjtQjun3IYZ9tp1K4
3i8zAwCIK9KM9mAMU8Tcm1BdmasSsQv5PGJ2L82BPjlOcA7R2++rbt6SgmRknbQ9onBuqH18RO1V
QoU/iybHtDk+m9nY6o/95xmt7/DQebbkYDzHufs7xYhlybslLpoMrMjoqzCmF+OikCd/1hfWWgl0
bDmYnkVubl9b53iq8zaaHzTSBAUebEZcFVNl/D0mtrspSftAcWJTK7cl/IOuhkGJ3NbZbOonySMK
mNvCQPwwTO/NJ5Vur2xDmUl+UekfX6U5k//wHPnSgcdSoHxaA2VUosbFFUjYGGYGdYNL2qkM2K9H
eMbKSDvxCnjDCbv8xTe/VL/XzPT0wQjtiD3t3DUedy9ufU432cHSAWMvQPdvhp5tDxFIoblOSHts
uVHlIEsdP1ld6TQmOzd08qdFdBt5+RNetNsXML8n4zGMDhyGY2MrOWZ6brZpAisy8gS+CoLXAYIx
t+ohe0eyzyEF/8w4Y1tbjaDEZdNSvD0n5NTlv60+bOA7Nl8WCvynG6PrTKu5eTSUOp5nk5a+PuVG
7rYAMgfO+g64DTyYBcKoz4PNabX33ifkdEdNcu6UmNr60SjBzO5GkI2/kBarwb5svFacoRDAN77W
WEc6wLElY6HReXLtrKIepAcOfet8V3H3FqabRtRyhcFoHDHUewZ4Z+rAiFBydui9Gqq/syngmRu9
D2AmHJnSR/ARGqNWKY0+D3wrrZ4xvid9zxZve76LIuVlalWN9ehnfMKywThQHpHpOgTqtxUz6jhw
1hA6UqRZnb2ESPImLICxvnRkdjzkCtsydFYX90uvSXDd7vLFKk5shhXibyXaruUP/S5tfdho2JNe
DXJu4spUfWDWGUPVf4XUXzjhN1+6sy8bdhisw7HJ6Z2ia4QwNM2rcqy/KrDddfYbMyrD9TY2RuF0
mPqUb7v9oF5lu7w/O7KgGAAN1MkKRWKCKcwWewBlKqMSESnz1H89h0lb4mkrZDwVKHbDSeOIiNBG
ks+R8XObUwhdoI037/0a8OHfKgyuVq9f8h6q2JxrVCqK63A/b+i2A9ZSD6Z6NE8gEUfs/BurzqKT
HBxH3agLgazHuibgjivoTDjepT4iJH22Uq2zxieLVnHZaXuzp7p42aKp+AoUpBjtBMsWZimR1+q6
ZFiXAhYYKA71/b8Qnus4CWaQuhCwhycMq5vtuNRML5Qcfs6GYo2/i+LCf/iaRoR53vvVQP8LEU0W
QHMcuZUCw8FCdngbSDNorlsmYk8td/VmyQ8lVJ+TfRE/BMR1donEt3q/wnp3v326WU0jrcscW3FL
nNDbIE7UouDAT6rPOVBOVBiPzsBcpmuJko+b9Dxi/V23lCUAfODTjpaNQ0U6f96LCMyB9IlYZi8O
3ddXTch/m4Bv5ZDppcP99qF/32dvwTfkTk4lXpFMnXgg3bnfygPTgX46C7NDUo3EeqkVK4G/7VSY
RhbA+HNvSrLO+HaUCYwTivasoyI39yMHbE9KF8t+JbJGvMnOsNq/t/JWQKuoFHenCkXqA6UkX9Ik
f4itP+aUKm4PM+lOMZaVAgawdSGiycZ30mIt0xdK/lcrDuC8AbShy8h5f7nGoegHaChi+O0QpI/A
+vXc3YmW5bd7ITUX17rDn1E7uIbI2o0PnM6vBriO5icNc0mK/Qif+3JpS5/GDrgZ4D0jQShnWFSu
XiZmg9YwMLqKaRwVqjGypddWYdTmTJ2ooAgRosrEPChFUW3qF5fOhqYuLLXhXx52IVvq/Dvdct3K
brKBGjIgguxci+ZukZ0dGWP24I/nm4ZulNWtYk8uZzUJR03dthCBCUyjuKZXXPSrXcYbVT+LqyYz
XSkg4JNeAZcbDMXVXlxzNl1MS53tD+A6UPDRDVkOjtWofph+gxYv8UytRXD8knbcfe9szvWCF32s
FTKLu6bi42Vcgx7U1gyN+g2Yn/nCiKVQAOONq5kHev5OMCRrqNZPwODgRqWrqtaKfUZ4RUYcQxNO
AqJ4MKHeQOhCTBnSVpWBncqiPAQUIUnDym9ljOdi2XgpfdS6OugUY6iJdzJMTyuFbyYf4BGvO8xc
Ysbce1LwXOwSzf3ItWQSEwHXybAPDaJTOxCHwY+OuSuWd1/54x98Jde5YZ2Cuv1ys8TDuEdJ/yyo
NLqeg8oZBlupdW+JKJUAjJbVYNq3pPqlTqG+aZQJ8UISj1byE1bSVF0F313D/UOQIIGiUhc9bnre
XQFAlo0f2SNEKQAWbAEbXk4BgBnp545S3xyShtVwu4eU4rOonQd7NjOdS7HkqF05ivlLYrjmON9y
ryUi31UbMq2RoEHvJl1IWVFojabwd/pc+CcBUdSVoSYYPVbopzLmdlp76mm0IgKkuVJxHhAEuxSS
UVGCfGD7e522Xi19f47W3srUNfv3Au1c0BewLcx1qrRwmlJ2p66Vf6rqfe5bDZJ4zHN+2P0tkXm3
+Ok3JbbMV2ZwdQbvT4ZVsDWq2pbaQM55RzG+QJG2ETW09ZPq8R2RssIZlTy6Y9Cc/70fVMRTuD3Z
3gCfvkZYBhJ0wKoLZHErvGa0ezAyScC3Tn/lVzsF7NurMV636YFIawg8EJY2tcYDbifHsJkIgzaG
iG8SkKzaV0sizuE1Nx1OhplUVbGcGUQOxxtsG06/OLK2Abh/yOhdyWmUYJNBZ+K7a67wW2OPmAXH
0aBzNgTBqx8YstrN3U21AZ0YpoGolck+JA+m8lmM1rbeznICSaR6cVIMb8j4vgfdQbHzpdaLBARu
4pxrXKT86bvWuRwF2YN7Jkhr0ReZ0pRpbV/MODXMtEcjlIEDjzNXQhZyR7IyHN8z6NKLHV4cUO9p
ObWK1UR/g1kwix84zAts9OeOs53pUs8OaEsn64ImyMjRiZ4fTyg+nI9RJMn684GlLRllqlyfMFHH
4qPVgJ1KCsYIGHMwed2ms7MUNBvI4VYgSz1H3uu/MGzXhykssS6vWNR/UcKRiBl5PaugXsDuYmS3
3SFsVB9QjGm6QW9yLxGdwB7ZPOikyF/0F8B/eOtGBazA4eDMgbABtC+LKEYhsA7NLLHeBEk/Ypeh
TvHnoy8ch3cQwPgy0NGAkC7a9PNHqTsOQBxbI3xmjIPC7TwHfE2YKzGzzLGttVNh6bnf5Xhbk/L4
if5UluCi3MAZktGZgs2thIvwMtwWhslZsQaVB5PzVZrE72E9tFOPmxjTWupWjc/O1KeEaw3m5FrX
F/Sr/dBuDm2IBltR1FFOzVKXDd9ZQgfBR6ngmMJE1OPTH/LGudUhU1pAzzFfq56IddOHBP6JlEpR
rqHvisE9UPVg2YUeUnv2yiI5Qq82niizQCYJ1u20GxnqGvjxnnsVA+fO/Rj+FMQ7+EP4FnWVTYVj
8zqttrdFs5Xk+YTe6T7yviqvI0jmT+F0UOvX+4Ccn2gJkBEhT2QmsfQcCuApUc3JTkPQVaObgmwL
jrs+kYyZ1KyWw36BGhc4avufhVBEsn7Szcget1f0RkNT8d9S2gbIvuliyqcKAScCyDqylkmhTqhX
aoYs0gICoaWFUmPSM5ObcuM0vsEV5vOE+e0J8TjKQncrDMCP0ej/z5eEBmcDiYNAkwrHkXxzgOGh
Y2OC1stuZbD2S22GH8OQ/Kxl/7glUYwFPEQ4NYtCjKNVSlkwNdqrKPUjJi2YdyCHxuECbipyh2Ta
v1X6nsIL42CQs5LK0lE44I6ifetpeLF8Yjx3O35o5mKpELZFn3zA6zCcAgwnnDQ35M9GuP3fl2gk
IFaXXG41toIJp28E5iGVbgL8GfXrhfdTxy5PQHbsfAWgJ/d9fJJe2gHvIH+Q8UXrqXZx5hrCKQOZ
jBKw1CY044eqcGWzk+JjEjnX66PhWuUrscJ/olYuVOYnCL6ySIo+nfkXaPgGkH6SLkIp6cviZN6G
m1VwjeIsxbE1kEHSHrm9dgzr26zBswvwpscZ1I13l9kNP+XBNk7U+tWftYxGCiuhDCp0Crxf2I6w
hlf/wd5fuX848txVpw6VVFV8MjBy+h2s5e3mHIxOktD2R5cenTDGkAblWxJinNbvO6B4wxBNmZAI
JGESlfdvG4dQMTFfufzlhblcN9rAib/4J0ck0IiOofrjTXBry6GgH4G3BveKHMAxQinLd3xODNvQ
ylJBwUZ19wpjNQIfDE8qqQzlxBwCiXCFWCioV3e684FxR41JVLDb7bI6+Ph9ypsgvfZ8kwV5B9o3
b8atsZYCUqb/DYemOWe7/hZZAb9ImSp+JXDGH8jilmSxq5hWkDKLWYpd+8Ks+7IsuXDode7YAjFy
5Q91O8gTOc0gzccXNF2fw+SNm7VV8wFDunImHJS9ZEqxRKLTPMfou3WxgWOFO6GALjKSpb5EFIvx
YrpHstE+iuH1t6JjuSOZ4Fm1de1S8YkKNz2cO3lW1DIoXIsk1EFOlba2w+2ckrcD9sdckTjXuS35
mzh2s15rdKl0Cfcn8Y1DznPIVY+WNeJwChs/Q5N/4myCsXOxQzY1TsJHLiCJIh9UiY0t08UrwmRP
bybkZ1+Da0tmmo34v2CVib3fvQpiHQCpMCvZEPrJdkzxGU3qBuMK5bP1K80cY609zmLvZSKYLYf0
Hm0tNJhGWpoldY4tBcThm74piwKaKMluJKdszz7hgP+pLJMNXxAeNyw/moj7c2gEbG2OYCxedf40
R/p4BOvg9VGc1A9BwQmZHbkMDU/aXVduP4gm2I0qFVKtPULHOYppYaUFCT5JPAfXkMa42GjKdil+
PlQE3XrqdeRxEo8EjKzo25jyVzOofjNDvkV5IiNHz4LqiJ3yg749knlKN4PSRzS9iBF87drl+m3d
sgC1/8+O6BVPyImW1cPTgRxTlX8MpaUi6s8hEY4uNxmbfX+2jpz+CYlrjVixCpB/UrX8hliLixL8
IyQBMXKJrPwfUmxtwxrgO8Z36M2D+U0aaA9vp/P8Q66xyRVp/+huVBPRknCdZzCXv00ZBXqpITAb
oD+5iszZPkhNCoYCu/VCywpY4GtRAxH6xDOl8b7tyI9kbQX8OCBe7ec9ts57opTOU/34HIUqKBgn
QwZQpEfUCYn0xMNi3pmHc5LmP509Pc2YVKcBiepKsypiPh1u4ORsk2T+ZhSkOHztBJNDK5b7rP4Q
dLeqb2p5OfiXs2BmVAV9TsRhVFG1HnKDQjF0N2HcYBppMWAedxlmx2s7m9zYxGpIcYI2D5C0Tfac
9vkyXe4EBuBpN/wLcWShiNyC2IExwkvGZHqv/m4HC3iMAL2qf92MGZEtej2VNMarxFvm4+hpYAAT
RpT8UefDUrxpMyL9PI7Dezy1YCMBSfw0enwFyKiDrzybHRznmGIwqMmAuGo+5ewbvwbIzpmosW6S
/plM0ZvUOkZSN7u9zGn6hGpkLMgh9vQHAFbVqERIUDk+RLIjzNwnqiLPe+knRC6PWPXk4MXmcT3k
oraOP2rfXNQ0Jfq8xsx0lMzrdDlmwd/ZmHrI6VvJrXdtAgJiZwAFIRQd2NAggUx8b4b1KR3dG6cY
yYiGz7EDT0qnkexxqANF/tD4FOzkx1rSao4cFyQhU84IfVEht+qsqixPdCW5dzDpf6HDJbVY0ast
NeaBPLivogw+SikcCtPVMt5xWBrRCHik9eFa9lQAkP1s73RlAd30u8/blPFXwa/RozjsLYmc8h47
EdIYNq7SYAOnnCGjrO85/+jOXpcOhHxUcMkJIPwpcH5oF/L9kPWhlAbjHk4X8Pl4dHtDtQRHWELz
y0E8DNvCkLzAs2lmjll8/zPS0nr86+I3KifVbWVc0PXGwLnQ2nQmuisGnt+8EeqgL5QDmcRGfoOe
3WevSZNne4ho3GEdQoyrFhe7UORlSikbma4Bb4Bw3r2Iw1+pMgYuDCpjn5yJcgK5x+PqCuiPl/lA
UyuZLHR8HPvTDO4kgi6Wba2gCIY0ORq1O8sGH0AFRp228v8OIEXUkItm1KrEO9QN+3/mfufdrWMc
5sooLdhhDyPBsWozP/VJcXCta46KLFsQWUBf1usji5Tvaz0LtFYSOG8qvKcCOV0dODrsfh5Max/Z
bNOQjg9nt4zFT+d0hyB/o+E8ZI6WXw+vS+kr7Eghb6jCdt+iyy4tkKRcQxWbcdf6drSTSK5CKKEQ
yLBO9Osu7j3uvhME1c+q5JMYjd39+l/avK/YqEhkIBriS5OnKoPu84PFHXB6JftPeY2rh+6omkUy
2gw1AOfUiNQERgB3dJqclISoAbyy2tt7ti5QHTGeB9V5cYjVRoSSWkacZm7uSx/Ul+4eHgYvjBdC
JqqkG8HU/t4bpD2OSR93mCoB5F2sMLPopZeJoToHrm/+zIL8UHfz1CQRhjGbw/oyyiMPDuLK6UKR
Qwcvvjz0JqPtO+hBgzglmgYu9d/Q1arS+uwxLpTz+tl/NUESa4ALBj8UwxKKzy9GN8eASs1xHdnb
8F1zohX67XEJV+tMtKTDuiQFHoKlu6aDBCd05s4Wx5PePuvlPd/7T/XHT7jVVtigzPAONAbOd4Q1
E73cnDjS51Rb49R565Ijdtfth0cXsOqc45VDW1s6gT7sR5+QBqfvJ526n2A9q1BL6Jp3hbzBlYU4
HsWv4Hi3D99JfXHqjRQvklUW6VAO5zcL8o5MXRHPwLNp6XjYkNkb9xGTqPoaozvc/o3RTZiBDyPm
PN99R+Wttw4LmoS8CaLl7g0XmjKeCavMreRu490XhBaV6CyW2cDlajSMWm18V7nRaKEzvDT4mXv1
ruHJ00tW8Sl7UWD3DRxyqVIGRg9QaF9c6tHtO2GnZnEzWywMFQDi7WrJRmCtgSTgjltdrk25/5g9
BBsp/iq5ZW/11Nf3VF7UMV2Yf0NbScyFNp63cAp/NIzAdmkzFS9g/FqmS6agSCyWgI+cu0hKNmcl
zNu07aetAtWeVkH1vvE7nWz69w4mKSLqVpNyVTNb6N3F1B0z3nRt9R0hVAX274u8fUcxfT9wMGKU
Jnh4os23H/OQqcXdWdSG07qEtZXHseiP/3LYp04bTgDTd78oCr4UHg3FnGJVRscci5/Io8ZWrHv0
B3ucGqnTgkW+024uwYz+GJOsFhg16j5jXBfFUgsogSgrVqhmqKuLgA/2ZDB+je9bZYRWGpmKRjL9
Py7+RzgLt9xDUp+2X/zzcnBAZbA8dBnVRLsIWsBuJGC8uqxjROucw3sAN2MEJvRvmhFO8vNayMOt
s8/VA+z+RKY89lUHKS3MYkmhB192+VlyHwZ0c3wX2F5m7o8SNh4XOEbbsku9PSBUXlFc1sIUjOea
dgaohkjFo0neLQQC+DtacSlRldz07OLFKW/PZjPFVa0JlwQFu/+zm6pmsWtty/2H/9KkODWLO1de
9a2e4OgzILCMq3ItvXh95nhKOjPSPwVhLEuD7C8DmULXEZ4snXK2odu6tcLMcep65QJEr8l7tOBw
LGhFIeoZ/65ytNuOEQ69zJ2iRhi9EYEIvy448ZbzkXWn/CW/tQ/BtmR45SXvuFElW3qlqNv0zq1M
OHJ0MSz2peiEshkB6VhtZPca5s4EK6Xqd7CNJhqsbRJNToz/LRfoupxCB+/b6hSS482DAZ5r4Rf6
mgj+UL6e8kYYDoWZuZ32UAcoiGV5W8nzUZTCO83mY/WKi3g6kkyp4hfS+T4tIj7QVWVTdInHw0/e
8for/WVDBpLoCAyJGWiCXIy6QmPtgyfLE1ZKhkRvUJUDd9iVcAg5opaJboINsenOxJ/CTMoc6Ll6
YQ0hJXlPCc1lgfi2NjxsgcRxEHvK+tox5QuyKcwJKQcQj9OmPJUDD2qQQ3YgPCgdvzIuzOPXT7vD
yfaTKUH7+hjr9ovfjA6js86MKusiIho6wk4XBjgvyUV2ui4GPjS7kFIA4boNxn0J7auRqG0VADrP
Q7CeCtMNZiDFg0efYB8IgRhaSulg5mmptJ4AarAgMG5+TVR2ClzSiu1uzbZPuedhgJIbAjRxEiu2
G+uwNxi6IgNeDt9b9+Qu2TFAa92dgzdCz89lzqgM4ngXsiqW4YLL6oydudS1x4eCG9UhlpV6m/6F
BDbfPGgQPeFeGN2vmue4cdVFvbvhJJb6TwzeLib7dAlbkpZlZKpYQGlJbCeWdawZGmHKDWbtXHs2
OrWX0phdgQhaVu2K9boxbksq6FrugL0BrpEfCGViN0UcHZi1NRIESPW+JQNS07tAKEwITMUcShqr
R0cS4dhvCr9USJRfYossMfRtJ9MUe3x60N8x/NzS9+SzvqlSanpTqE0OUOgBSZJ6J22qa2oABM8+
JI81LulEbRoDmAi6Egc0/LwBTRGom2GK4caI3+YIJeOZx4qkSnr0invCoFrG8VU85cu4uwmxJ8Ak
xm6w69uYmUjeCDcXhQe2/QM3Tid/0LQx8lp5sZo5kYmMPrZumdfqbnzjMuDsaEL/mdNaZCFs2h9D
hlNrxXCgtUgDL11ww9y/c2MMeHpdmOmetlAp3qOrEpjf+ixrF1qLGO1TTiXnsZZenIB7IKNVVIEo
IWooo6lgGDpqLyBMBcsg0TGvaFPLyzl+P0Zl+SMWb/E7HoKzY3+o9JGO9VCtA6iv78ijNb/63JgQ
RTEWKDVKe/H8wGApqB0woZqLjq1eLmGinjV8pe9eSEpwSnwOWJzIez2yLSmzsK46w7fI2dtXz7ci
b28CHjW326h/SodIoDJnba0IJ+Gw2X7m3UXtC26PCq1Kkx3VDmyu6h0pUXtmYQUKkia91n3J+ObO
fIEU6waKqL5MlTApla6LCNZJL8Mr/RVKWvMJlq+v8GkMFCKb/bBj0iGA3lpJy0JiSik7zqMb44n5
V0Bs1mB4gChj3vZqDkqWWMJOB8a3HZYkZfJB8JKFEoN0IiqDOqZtp/Hf1qFwVSnyV0dHcTVV9M8p
Q1D9jNfW5a/UBMDhZQBCqehSC1CIR9zeQ31ke5fY6DnPFNlUN15qXdwgIv3+6T1aOaDD4/do4gBr
smg+pxTGa9msHCk4uV7IIG5VB9N/Az3PwqFzLDwPeQ1Lufa/O07048tunPv5RTXM3zPS2HlgPYUl
539YX9Cb1cdMB4XiHGy/LFtEK/RQtkT6CcsuLK9q2TZE7ZNk/NiJQB2Ik2HuJm3skbQ6N15D+sh4
7hwOMHqhVeWEF12s8S+xIpNUGYKK82gquSPyqXxev00Pbl1FL8bFIENJG2E78OEVqcA9j16Zqdy6
QdsVbBvVpf+hzJwj9RJ9awBuD2rKzXyr5bOblorAMqQ/nP/gDmv1q/2vVnEnVwcwkJW/zID6ND34
mdBuY0P0kx/O84MdsFJLhriKfD7scCm+kUkZWFfizo4OwNWZNzQftRxIp3A0xSmJR5L6e0+5MBZS
30o9cPgzw+KhKuRg5G9TSahhu7yax6ZRUWEbESyLOT55zi0zt7HMHnbpQnfv7IIlLs62jRZpR1sE
Nolm4Ke/VZFj55dIpgxmENS5CgCgMH23CNN+4zVfaoCGG14IKd+/3uE5FBeJ22zYzvYD4CoiXYKA
yRv0QeN3cXXGfYvEfsZy+V7a4/++doO3u45ydOU6wZIvW1RWq0pzJnlG3icNCndffzHjFZWqiJVc
eNRSdAeDmaIh98hGXa2/jUR3GDswOLPrFi3SKwCrxeqocwYvbUlEWLsVJ1BPJaHAgeZNcplCK46h
yKLNz9hxgDL9s9gASsIp5yKINX0d88L8DGsCDcWOjepkrxKEEsBacU46YXH8ikKuSbL4OP/EklwN
NsmCeeZVcIdM72w5n2CmSblTecLRIfvc6eVeEQWbQl+EN7kFsXKlJrTO+eqjdZJHEYn1EPQCnVyI
7NfEzn5oFuEzNSBYK3xGmsRwalMJdg25KQaUdQDsqh1hyHwkcI9bC1Ebi2+BaRSEa8PK+Js7MaRP
Iz0LHGaYv0wZq27yNPzhH/yJpeJZFVWM+/GthD9NKUL9zIVFb197h5NuJmpu2QSDglXJFktU+rsZ
bPWDpuNN57h4lQgyVmJ75QXTaCLav0bpyStORuAz+/tWZTbDGzMZljyM/ZVnt7T6ehPxlJ9Q9bs2
BhwflLE+HZ3nC2nR2OapQcbOsoJNJ54NyIJr/E9onpI3UnOVfGc0kCbGT9Y6qAUpTuuml47xVapd
KoKJ8JoLQdiAv2gCTlNfN+VQFPtzuHMT+jnxi2No+F+qHVjmMk09U9ySIZP2T0WuDezIKHnSv5BW
QdyvMctgoCu5w9I50IsiswuvjEU0OFNV1cltjjjqJ2yR2iiuMeNT7GFhZKNQSbX2D+Y/cRjFrZXO
S3PTxGrVL01L7ZUTEgTEzQyZSCalfw7nBefuKJMJfb6yp+0xMyeA0eqUXzQ7c7Cph+lfQtWlDfEk
K0JzktKkThjFL9lb8tiJt/6CLdQSBnDXt4BDreOLxaDwPj5HbkIzDxNdYrp+mHKcJlahfj86k4Xv
vE7ECwe9RhcdqkJHjWZeAZRF7dd3ufZytVorMtKvRMhNQkySEafcl5LdybJ/b7FiZ+I1q7XsPBUF
t0BY1wglm4VJtr/nYZMzegkPEG4HZVvDM5LgyGzybI+fweEWlW3Ck3Ojj98gGEPc44WJYMHGnuM+
8VshWbzC5jX5Gc8iQ6QS4xBtNBPkzwfU6vrPbb1XToy9ai6FisqkQi1BSXMGuOH1nIsscxWPezHB
uvq+oUfoEDYlpM+HIUV1YCLYehJgpMY7HpuKR9pVP9P6AJmsNBazq0+LVQ6uSbiHkNZDoB1Q200h
HUN7QpwuyrX1MBFjHry15UADQ3jZKofCUonrHZDpxSjm0nkqBqvz1SErsDHcx33JaL+BZuEPMMa1
a/qONsJHRINKN6egdB0faQH8prjbsfFbUxEw8Qvy26MJPkSZGwQqOMqo569kPeR+4+ZmL3fWgs4U
y5iiowDsCTtdsg9yDZqlnRXdiurJ7w6ZkHoire4PEMUCM1fwhZ3WbXPiiqNETOd0OjO6EbsBfNdI
F4uAGqpVpWg48h8hczCf3gMP52fP563b64rM5DXf742syzAgZFRRf4zQK3MqTR/9rxQhDd4LvE42
wkCVcYXLER6MY4ktLsQ5Sjl+5QRlj2kRsERApraYs02bStwKobiTvd7cRL6aKz+8eIJaWWQQgdxW
fkbhq9tVlFqscADnHc06OpvCj8ZH9e0/AOrsRJlqgvtHfebCPstd/GBNovMJPVVNV38HQO8J1TN7
7qXm8oBJZOqjlzfquyX0WzyZttli4TNG29dBz77wko1PW2KEmEf9vgS7S9QiPE8Z+AWyFm+jk6mb
ortQIhO9OvI5DNm8HXZGxkm3nornsS6ScxnErxXLCbYaGeCzRTguwQpnNYebTbVDzA6ghVfbcZqm
7fLUnveLIxQ7336YePUkjM+Qdin54u0MS0AAx9uOjRlzc8wSMdoispHgv8jkACpJMa2yfzZ7XLG3
ZrHQT4eBmdfDNBgsnbzMzek1LFd2z07qDC197GmQD+BQpYm5WbhmljSCf2VMnVLQAVLx1Y8JEgxp
XwvpU6yCbFtiydWAl/sxT5UqqS4E3b3FxN7G1iItdqtnByoszrbeYIaLprCEBuee8/Z74luPeV7T
MMxqCCPW6ne9C2UtWSguiHK4yNH4fd0eNCm5ZjYxBjjvtTm3ag/S7R6RjlsooRR7uatjnNNH1HIL
6lxpHqt0/B5acKQVTAJ8S+aImTElIY5FtOuYYFSx5JHcrkxYgLbFZB2U7Z00WD8bPm0Bxrgaa9yj
BDyhfh63lkyLLZC/vVfNW7XR8iMuiS3jDlACY8DD2gatGl37tXtirW5BbZIhvGqUPDQO52b9QX7m
6C4KZrkMGgkU93D3n61Hz6fCtirMCStM5LjkKMZSUErh+e5gDv+5Kj2avsZtethV9Dqm6XMGyNfF
DCWPNIm3Z4bLPbN0UMogfXQsqjK8LQRRVBBfS0W+xfMSakwqEsWaNUCDdJ+DIzbPOqNRGlSmHpmb
cejKGU4N2mqzGlqeaHZfoKxmBsYdfNQZ+k3XEtTeOro4GbE+OvjSvejQICLdFVPSd9AlD7NRJh/w
689gzzvfLPXQ5SkhEsZ3ZCivMAvdJRmUE/bBsdnVz+6gNclRUrh/XBc5J2dPfwGfQr4gM/om7YAi
gERdop5sybzdvChkgT4aGTCCuymjDazYDqVy8U5PnlE+STElWQulCYJE7mI+shKu9Ta2+mAqG6qd
CsSD//moQlvvdOANA1Kx1D94Ka5B6wNWmbsjC14KuI9hZNRtqb6jVdIyDBHzVos1hGOF+CLKgHhA
E7KHaTdxK/EdXQK6OJpe7Gg2xxfkv5RCtmuVUVpRxZdCRSZyPRRFB5GYBU/hYJ89v7Iy6tLLJ/z7
oLgH0eduVBdc6fDwwUU8aXk+rKibp7s1FXIwBMOf6zVB3IsFVUivadB90ObBMXMs1+OJqLTvZqQO
uYOWYCb/KPpdWUCcLubXwrbzIj7F2xqpmOaEE6RwKnOhpayBNAu3sMl3nZMIQ2ES3dJ9er+6ck/4
9JJgaYYp5l2dV67DR6V1jO+0UK0gKMas1GjOpSRyMsbMIHSYDVJFBqEUtY34M5ajM1wl5uXpY+tg
v/kT7Y6sMl1gJ3ZQMiobjKBIbPaGVkiC/rDe6uFYCCCqUeqFjfcu41ml9THMuM0g8PJrXCUq3grM
HzrPyjraa5vctisH/07v8BByarFmfztVj70ysV7d55cIw0pY92nSeQXWxr5orlHeGQLpdAo8jQ/a
ZvOg2mI+bhBObGOFnhoy+3WhjxHip+qVpciDCGYDZuPpuj5k1Eyp9nRl6tFwL83mhFrdSQwivuYR
GV/bJULmb2sfvoo7fV6vn3owa3SnQITsPDZ14Jr4MZ5qyvvu8eWSB43R1yt/ZfLzgQCXD7BOwkSX
wzX+mP6ba1ATGQvOUWdMn2o/g7JSE3bmyB/FvbIaEtECRocZAn0ZiSzCdLDmOGdHplok7Yfy50tl
B3lKkY+/8BP2AoEGI+E7pLhPMClF0nwviXt6zqT5+zYpnNq7Ff/cNBh8F61GHpxtNfWBwHmR44+g
Pww6Oj3RmAz3EeJUcXuA33uRUirkg/nzaf3XKy9d8UNHHJ8pxz57jNFRjHd/6QT23Pbt9rHwLdVg
NRchNZZuD/htgQN9EuBWPPeTkBRHNxmo0/xesFOb1ne27uBlCNrylsBkodGTHl058pwAl/doNYie
lgbEvKNmh0nkV1d8AqTY+ALMFdkQwAGElMO7ZOgpq9P85YkmQJqVOTBMlNMN4TO9vhLm9wpOJ1Sk
YvPZMbi8A7H7dMpHB33qmSr2UgPmaSgxLzvzHhhb7N/fSDYLhaQBc2FWfnQKMVWrKnWt1S0VPs/l
q5Xic2bjJqqvKuVIIg2XS/x7jD7gkLU1MkbQyd7AeDLPvdB4Qhz56QvSkGy1qYqBR5+sjJu/8Fwt
fC2DnllS4sYpyH2CJHnxL07bjlb5JVXy+1cosV7KzWB2f6WHmeu6GP158KpnCVLktaNHlXu/nTz8
7kBiZUF69j4zYu3FTTEITcUbPvg++fO0QIxZbMUWM0NJql+jzBTRv9+RHajxoFXLnlK1+D/kEX5Q
SHdMZo1NVTRVFiS6UGFnKj/CfsugapPdLG+CWHq2seHY1fyxDxNbIMDlvt7DS9A7fOIdSAcHzWHV
HkAn+61cFSBo7gmwctrmSZcSon6P27Yz+/68n1R00qaav2Vn6tvHVOXXBruiqHgQY+MM6WUT36hx
lxm2DP1YaLdfnGBkbWv5np0xA1iA96B0wTkX78gAe1bF9971AHKCJ1GXD6pnZGwfiLJ+lBqcqYVe
MI13WNdOD7XEBl8I+F5X8In5hJ9lCIvT+uY7/4FANTitC0zuzp2euHGiGXQh0QuiXq0zCNcMlcUC
uMLaVXg6LXDRYziyJXqIjxNrBMfm0fv+k9ByefjZJrNK3ed8cmDXDD5KGU6rnTt8kmEhrBSCd4eF
EsMdyeHWfLG5qNuZYkpJOIa8ZPBD3JQqMcX+tDUlsqFwYtwn8cYTSVQ6n+L9sidWgD+cjEivUYFO
aE6FWzi7ecUOSQ6L1/+LhRl+TnUV9P8BxN3XbVtHPHhGm+GKjD02CFZIouI/tH/knIPKgh+zmW16
qJgXSncHSwnDd4UFXBRt1EpDW6YASlTNAyu9R0u5BI+l1cuKgq4M/vYXCvPsLl2RFU3TgBEfgjPz
9LIKwIWN/3bP5gbXufUDdorz46ZLY5yzh2s6IsnY2nleqDlvcKS9osxBy3QKDFEWOdMqlVO1PXWF
79uQQZ8IzcjJ0KT8gp1r8a2/UfhntPTP7AELtDIPV/ZZOYKoykIZWq77z3f2FtdHlH9PuCjdfoVY
nQwsUsVtQuXyC7FAhEaMo37Jh+1B2v9CCI4ysHnBlbgq1MJpf6py0voxmnvpXZiMOsCQ8+2Me2le
3rfMq5Yb44FHc6k+1SIQvTN+W0HkNS2kXhPrBrmWB3cTML7YgWPUjOFVUutKQtIlPU0E7QvHXKs2
V7IK/q+N53gpVkS/sCJPr559TXFuBJ9652oQo2aqGsxCwQjdH3tzmudG/ApMEel8xbPv4e0aojna
kKmONY8QVZY0LTQwj/Gh5DNq7FJKZ7tNlK7qvj8HRcPN4Y3pWIUQej/wGhHBGA3oiEkF55m5QDbd
/3pjAmZudIup63wSmKVhHGAhmQP3T7uFJlKoF7IDm6DclWZRLse/SDECDgObzYoseAr2fmXlxrGY
4sdKnWxY3wQizvT7J705Sx8ShJqKmzO+tiDY9LscmeO1jYKXvRI6LtMeq6UT8fv+BgV11aR8/SA3
lepWm9KSySvmCeJNxPfyQgOW1imb30rK1jn3AOb/JdeIlAfQgKIMYrzgoE2Y9vPHpNn352c76zG1
AOCW4NBjkAvM0TZdd2KklP4syvc2vEAsYItVKhaGQVTUmtGP4TABpLom3e8rR0UobkSHH3C5Sa8S
KNwlXJRlyrKyXN5c11IQWSk6i72+apILiu91/qel6+7v9kjdfTjIE64fQjdNtjX9tlh2GsJ2HGBa
hSlzGmjvObzdouZyzYrhtxk06ZB4oSTlTe3/FEuObkqRYVybBk4M3j3ZFbaX2hZuw7O2kKX3whrq
WzPgDMMLLyncBxrkdJOc2/NPZ8ZAqpEGEwpo0oXSsGeT9cAuR+mZ/jq272hshyAHzfkroAe2xA9v
q9S5Q3mb+6+kTVLwT/yumey97URWCiJdmNYozo7STB/L43eaBQjKwMHrLRmVYDnAZy4V6uSFEzky
iocIzxGAM8PSwa1aEay6FThIiS+Iaa43emQ5JJLnbSjVT59SaB7GisTXVatPLblzZoExoMD0TZf+
JLcABRip4O6ZUzk2Qw32b0o2sRUNr1/h+H1KAU+/cKiSXJ0/8HQCBm9y4X1g3iYUC9UMBIl/in1N
VSt+jWOH4EWnHMFNaspLhm/0PcSdZsiC7PZ6PX8aErvyp3ug+5kkQKRytbgftGV4yuXlIvhS1DGQ
PTgQvX9tAju9zxMukCqaR5VwH0XQSHxVM/dO67GoBi1/apLjwa2qnZVt1wq+7xn/Z/f47ENgsktt
SNBc410HbUCm2Us9VfGxZvb46oPeotOlecjn7DuffsByGkcvVz4a27U3RyzeH5Ve05vnbCctYnEX
cacU8mVG/COTm7sYXaOjLYFcPzGbf3/JrY5azKoPnQTAHE2WwFT9WsOHVVxwumuFd2nHIjW4PWc/
mDA5XMQl2OMg2l+dyTv1fojX4jFDSQ/z0HtKySPXY3sz9NeGjqCGyBgXMJSa7gOTV5lo1I9Cxwuv
UyVnNK/u5Vg4mzu9hwzsPLPBvnumQx8HxGhL35eqWn/GdN9R2Q2QJgJjKlyMRDtRxnGev5cMG9rz
QvJQsUD21ZFu25Bi/Ozf1dGMzvW+OkEj5hy1x77ZPttwCvWYML9yqkHTXFQfJYQSCHl9lcsauKsw
ZjyRROgONaxbpkkMFkFXT0KzLNUElUZ2w1dNTmaCG7BK8Zmq2rlkwv8wcAM6qpb1bAEy76nnKoGu
rAIyg0D8xKLMIhqNtpGzNxjKdXPO1+GaeBHrbJbvPZXs5irG4B/jf0XDUg45g4hzrnll82DNnBPw
DfHvmFNGVdn0li4xRiwA2crTifFidCTMLcNVpSsOpr91/4k8V8DMbygUvp+jprZsvZjx2vPG8KBD
McW1RNyyzKF7kgvevdvKQ9+BwEEfPy/5U2v5kOGpLSKHObySPobbZ2cEIJSAz1z+/8+IWRdwQ9KV
KkhBzFmjqXHog8CNC2pu3tI1vkDBFRQMdVSszi9u4K8RXcemoSKoXKJwE3Ij0MsmZTYlILMhEere
Ua930Ze8jm4Bt/64AoiHr139PDfgG2Cy6crZ4R0KYhe5H/PGumbA1/m/5ZkzHK3usEadrI1RzhEb
zlXHvzAdi+erNGQ0LKKpnP+XWhqU59DQ1pE4E+F0j7PFdRzENbaKz1hOtbamMmdWluhb2dDcGlCG
Z4Dgk+idsXhgwFdHPCdc4ISGwIa7+dnnjTcKGLVbhOXO1EgcpBILjm2Y1TlFxz2l8UAFvqWeTC4d
xFDqxHQs8oTsxdK9MBUr6BZLumz/mpe5SsPf7ASCZEgNbJq53hewy9NxbmjyK/EU/C0yBZSXWJwr
857MT6ruRHTYaCETOoFCC1eGEN/bHYg16NJD9PBuS8YHWqzwrFq3Yrm4P2W6jXnLsDAveeG0s57/
fRTj2iwuzyFXB4/OCJ1BKLsfulmNaz5/HUPa3KLWHkY2vFjhyktcmDvP4rL6AKBElfLVL5BOVLcb
NCsPPCCJQcZjjVgf0R9bMvAjtCnG7n/5F6/xLtO4ef2mc1rN+dbEoNTxAq6133K3/ISTvMJLpGLv
1WhYQvaDALM4TE7qBhvbvNXQ/pBWVwpD9ZuwHKjgjkgypYInHN9hxgaV1KMmV01+aKhDzAArcgf7
xEx4eY4Y6JIQWI7faQW0X1EZXVPCyS5Fusni5Ypy//QUKZ64DJZhxr4uLYaKcReK567YMDKZ87g0
VJs1TWtOR5z3cBGbhkWbjf26+b+lQooKUGibD8nvBrBxqrjV0dOlCkDBZYx+FE++EVkXhAtSqVqN
9IcsX/TesfC7EHwYnM40Eiu5w0s8+Lw6Niw9rwyjIwAuwSg6Oho7+BexVQoKpeA8YetwPLGzQ2QZ
rWb0J5CB+dDq3UU3uWxQtWQsxcOqPz/wcMZESsqGvT9T0cbM++2NvTXNl7jEvH32LbcGaTwL+MpL
xwMfWUA26k6lxYM4NKD1YNnWLBOwsYDrS4namZsLJLY82KRPl6G7rlAX/HdlL6vGQlUYiFwvjBuX
EKHo2gaj8D32hncmVzWIjbtW0l3RXCne7ek86b2s23bm77/4dOiWXgU0Ioqb6MVY6p9Z1RGTryxH
zHJOoG8ukyONbDeuyuANXBuwoCvg63AHrnvOSECrFNcj7x25dAg4wBKksG1dlWHlSMG/uKeQJoQo
C7RgnoKRCSkLWNI+iRch50349c7U418GZbf7HNAnBssUmd/yyAG/j+Dt00Imz/13XZXWY4j9fov/
fJWQr2IBw8zNwGpavVQAdwj6p4gHYzlImHoxiLo1Yo3p7249hj7G8+KGuEKQA0eOWo7TPJ3jzDCh
5TD9hUkv/LC2NEY1F5fZHqa4fZB8Gr9kX33SReIUMjfr9cy5BslPyGCdqscD4allsxUkwkl+VSoL
aobNDBtvZ4RKZHLfVmNbvIuGmGkaApdETDpLOZn0ecR4+1RJxhTv6jzuhqYa8D4V5hWiD/rMt5ev
plsafPTS0wIoELTP0XeHJ/EZwg/Kww16Rha8FYl2UUsYJKzrjCpDTYTbuR87Euo6t4drFb13y8cY
v4+MuBQDZ41is3VmJ5eyTn4NUP4fvy2aAdPVEopkqrCeszrTABNG6t/qE2AzRo7t5hggL8sC+rns
HwkPoarWxv0p7eLsbmOnt2SoRNyt/Gn586yvgZ7xpfdzVnNz++vQJZCbqlFvvBFjLqmpF3Vj39ux
36O8SVliKWSk2ZQqC4jpUoJvfKxqD+QL9Qu31s5xf39Qb5e0s4Hd0wJiQZPVRyPVBkS+ehewYcyL
amHHod39y0JsSAOq0Xx6XgtoKw5q24O3BaKumix+lMRfBulhGgk/KwkWeoOqGtTXllNCDjk70ZBz
0So6cfunZyUbYSI/JADxW3JF0oInh0BDPsJjTtbhFMugax5EaSA8FdxC8URtxaAgGyneFfxX2XH5
maHW7iGI7bK9bYZP9unXGT+Dj+SX4zO1Ww4OJXIJQxRrwQXvwe5vvZy9id0V6EcSX2W7rdVDzjiH
03FqlTWvr+4lvfJch8W4cYn6reMWZcUy9Z8EecddMlRe7BHGD8VAYqSdUJfcqKDMFD6VlpfKyr5U
t4aEkKBGsu8YDL9QKyFQvNVd1Rq/7tajnsALlG12g3kBIeVjkG/reOAWJJcEXEqLxMJYBbaN+D8P
tc4m1OdjBalSoa9RZweRZdj/3ILrpyPuIzOHgH4RyRy7op4UFPMkqEFGndBYjfgqr/CyjzcdwLqU
v42U63RDKlPojw11ReTl4GAj0jYDCNxFSEjuQuTqGK+aIKFq6CLysceYT1yMz+Galk1Q3dKuzdXc
txIGmfPbTlkrElPS9cX4FIOeoA7h4TORMnNXTye2C9DrSrFYK7ATV5bDLUbZT5yIvXOWhgEsEPCo
TvYMe+66Irm/E/bDMoc+VB7OXNJbL+MPe5IL9JqJOUXTzilVP1FMBPzOSz3AI2CFb6COv5UNVnCz
MX1D20O4sz663KYHr5OV4EjRAvDdlO9aaDdrjmjCl4U0kXxaLFxlm3MRAS1F/pRELfLH7h2Qv2WZ
AO5lnJ1m+HXgVJjJ04pAIEkpeOCmlASH9go7G0fo7S12uw27mnM0ZWQwrrh7x2pHj/L00PPgtyN5
ixOxpKGkKV6nhCooXs2JW1988XmN05vPM/omz/piKxeByLuySaCx7Tuo1RrFp3pnUgESj9e6y+pu
vDyuG5WBZjyNpwjoYbVuvzAatBFuY0Dw3HxFYOFnmLTFQE0/aKqgNoUKzuyGS15QZve7IBmL7fME
oo72iVEXOAtU6N55Xq9Q6jL27yODwztcfhHQWgQDnF9/5b/lgZWYoa87cClcZO5ciZg9PM/pNxTN
igPNi9FqKWRMe0SZpeFRBkHwdeOlRHh7oMJwC/wFUct41Ij7NekUQ5qAguIVve83GSr0T1VstuMa
KR5LN98ABPNJlpdtANejJsSVpH9qFRQqIz9ZakHbM0U0hanX3ABOiML10CJ3rz5/PFXQt6thQYrx
H4foLYQlsXXWn6hPfgz+MmU7cTnYzypHvSw4rjjNE9cdTVMFtx70Nbir2nLMmN1neFIqYMP8Ufq2
QdINSRtD6lZ5RGzZdMmR8nGAZXDRe5Q/NxvsNKQuug6osKfsgl9Fk0R1SV51OYLWMNnKUeg5Oc+k
sDLjmP4DkkgE+USkvPtmU9jEv4JGTuP1dUfMUzWDOjm1t7dqtPo94m4W9xpmESggxDRokwYHIQ+y
6qVG60FA1T3Cx9SZ8e0mkUUTqinKOGEBxHZJ33ijD2ACQC0DQwDNnGDVrHoTABHwDUllC3fLyk8h
DuHvztZ3FiQOSQHi2RD4gQWVNIW9qpvy2JXeMAZZ0H7EuLwSctHYHmXgyUmz3n4gxOURDMv9wqE3
iGC7DSXSccVTyZX0svgkMYxyi+2X7cqrSW3bDDt7Z85VFZAvkdbnRxH+rA9j0ChplQKQ/Wvwbf+E
nfOlzi/7sccivA0nDXpSuFGoon0qdxRe/9Ec+g58sLuKrMvz/VveN8alEO7h3VEfRIhcCpHGIrH1
FYIHNoxZEegoEYAF0vyoKYwkIpFWiw7KraqW9GHvSp9hsiHfcBBm5DBdtIrXxSbMvaRoNSTsfQ+g
PtaHjncF41CnqcfsXkgaZmj/vS1EpsU1pcHxisBW2VIcpVU2VPpy+9fvHwNqrYL70Z3vw094GLuv
yIcd6rbC8YcOlzJ4QOOQkg89BHzIAdBzJFdyOUEU5iGBWLqO+XDQSbmE3YyCDSV7nVk/rQBQzRXq
aWXRwsac6b/k7oy0kcVBiVIpHQ79V9f4ij5XENn/W+j0ijXGmyx/pCS5H2hv0vclqbWczrY5cU3f
jvdUIlf1S1c8610IYzwfNmPKg45LMXFOcdqgb552YPartauLumqIqndq/RROjiBFH+T2Rz+5lHur
j5gtfh9WAYpQZjgRuwM0O9LrfIe1ksmWFAs1TU1u3gMqz7mGgFhKLIrrrSv8Fe7cx2I9R6j0uKag
axnfFPHLBPcvgc00aLxPbrBKRtwzcwNO3H+2ofxEFzjcD6FSSP97BRYIEMbozex14n8iT6nGbsdD
qsGhuPpUGFdnjzJsDxhHA4i6Fc0ke//UWwmEhv8L6llgOc6TUrQUDpWkT+KfVKFJhTMBICax4drO
PYdiVcl+ZsDNecYSW9zHALiG/Dl6S2E9+PWGlA+s3GJlt5YCFfgdvarMJJ4aH9QPpshG4/JCTX3R
MQaOCJwP40CzDOjwc5crjjtgHtXz54KSFt+6SPnYV+3wSe2ldjc9OxCJPuQf86Kn0rb5QIOTe2rm
ZFzQq0Y3b6Ayi+LMnG89lCiDjLGSboBbwvAPHLS6+Wu3BLqg1fD23m6QXWmmofUn9g1nBnJ1vuM6
NCew1G/XzNa4ggU68NMdB4HrfyFOkMyefIxmNy9/jR6CIlFsxs23ihA3CUJPnzZAMaFTMWXK7ATB
8z395X6uVJ4zaaIqv55roF4EPdjOY6aJaPtvbFEPI24tOMHPm3ez5JSvtIJgxU4pM200B3H97buG
Tmhfa3pAEdN+Mn4+fm/IlLCUWYPDIWFsa1DRJWDXe5qdX3+5pzXeMsZB0XifPjBW/2b0PJPTtZYO
gHVrBzC1DrQpN5znhbqrhVx1TYRxzAsbFyNNTbVwT7yGoiN9QdCToA7I5fxK6TIJXHTDzT4RhHr0
Ntw+HRxJ0Tz4JmBWvaDTYVKtc/iXMK++Phr7UB3+Vz/Xwvd/Wa5HPhAIUPEiqyOo2S+qh1eN7ZAZ
q8jVG3z2JprAJfJH8tT8yI2fV1karVRS2toRauZLsYwUAqL8c74vWBGbq9oU7ge4YgAervnrJ9Dw
CAG8F4w2F4gvjqa1C1tOvgMebfkXsu5vLcrXHp+BuRvwZJK1h3zXAZFranrhqooNvZfU8PvAa1Y7
dy+kxWpNN1WNiPdoDqLATJqqlbUcCw/F5VTe6UtzzaB+LWkOZJJmjYNxZ3Oq4lWxNLI94yt1BSyk
M1jgkT2D6W3ssI4JbHUaQSqX1IbBF0z7YFqDsbAcLiKEIwSlIC0hHeaXWnb5H5MQGpDO6pemseyp
h/T6Sh0pDsShyWPWYZgTQD6kcIMabCNsoim0DyAKAjBkZwOP2dSRLsz+wJwfJEkl1aJumAZb8eo8
q0FQLOiv41PUYntV8wEMsU3LcW3KhjBvANr9iNF1QTwU3Vzl7QvLbq7qX+wZaIzusE56T+3gWkjw
gW1MpU97AX+lX3PbYseIKtPEg/eCbRgcD/8+Jsu9a/r7yHsEN98jN/hUctmrzzNUIIhd2cW4glJM
dks/Lyw8LO//osnMBEzlI7XO0Wkzyoo/rwtoJHWNpqt8c8L+/r8zKRCyt0k2ojJqalvY/WTCqg2+
Utju+nNkvYeZtKby6KjRkpneI9w0KCBxw6fBbG/d7KyvEQ7//G+S+jCvKWHmdKyhcqjSPPZUnqi+
k5jyQ5dVdVyg9YVHFjalAmC2/sXs/GQzNi9U8quUi02aISuCzfgjciByWRwpF4JCvc8H89ZEsAMi
6PYrAczyMihajevrUgFp/9+MgESUr0BQkns20AdSS35+9CT0jCaTHNJnArpVKUVbdTbrFcQMytNa
1IcXWuRhRbZs11NfVZpZICQ5xHYlyj0uw08dcgUydYSKzMDLgbyK1aMAyhtUwuu+VzD2qd587kVY
w3irWEWjoUh6mxil64PDfCin45UvOR0TYIbdd2eIrX1AZKr1zvEX6/60xuTqmiBb5b9Fujj1dXLW
D7VdZxGIPUCKmVUEh7ySfkQF97/oe+rrjXpNi5W7EOxt9y/gJdwGCZOmIdW4LAMCS0mDY7RKfL/f
h55rblsImFiOIwyi5LWiAHO1pbsCtcUhiqExR9Gis/VPpFqu42sAZfBoU6p6iBfosyhqJVfixE0l
wnF9y14c8/M7eWtHkPV57GNcGGtiCIWKqhAvTxoYSl9gagooXOExRDhA4+wnWZUBr+GjC8cbfb1h
eldZYMHIf+J4uY2YwgEoEOb+olv534oUhe1TNDEHayUpvFf5MeKOwyWmCPj8zhenDDviLIRSDLfb
FDOodjofcaQWl6O427vp2mWMJPkXfYbcfdIldsMfwbaVq/rDVT5FB4y0fubdpSH4TVOQhOZF7BhF
Gi1BVGXMFFeeoG9skamo/VKPqXA01WZbb1XnReuhv+DQQWpTJToXRmVvLWDqJG66iVntvILbmwZe
4oWu/FHwm2sXFzEzi+Hl+4RG8coVN8+BQ7XiBzlnWuMOQHReK2b+BsLpFYT/qcLILLqoiicGGduv
JepJ0mO3wOoB2HUBBmgwl2VuWexjBU8Ie5SSnF8PPrf1gYYjk0RljmtAx7ho7DQ0Kz3rfRPV5/Pe
jm/MBo8/exOcVE4UlTus99pK6wjP6MIdSSgKLBvkhKdGNz50kB7E0eOnvANT3itIi2cWt24gvJ65
uQUFW/6nLiDdCvgxLdoAsS5pG1fxbBHgEKXO5zGY+/i6x7DYaaI0orSTmk4cfVjPfguE9M3st6lU
rluaOG1ep7dz7ziH2Xpae8fcbXjSXVVvGYrPe4vBY/jWoDcuI52fSB4/O/s+IvcZOs5WRVZzh4T2
vIsIjEOOB5VStvjSsetbmGFUTyor0uv0ZW1juU/GgQAKUUZ+kGk+IA8RkFYXypxuri738QEfBi+s
jpoSbKv1v1P0eaoOlWe6R0YTVo/oDs9O8C7d+1W6wSuPbMDL2masBOn5Ss0uNd57+9Un5s3hO6xG
nT+qex1ui1olB7nyhatgeSkvNx3aaLQtGG7XGovh1MBcyCHFTlLvOaivFA0HA2q63p2qzPfi3K1b
Xm4UFOYpicHbkzXd3IVUGaZiq5o4WBzZY2z8Ns4dLZ3+fDLrMe0aG/TSWrsiGfDP/FMRew/S6kQq
R89vLqE+Lkx/xE6iUdc2Yq5Dld3mSuXbHChDtvJtRir+gxxrut07XyhIOMTHVB8ZZJfRqfrLu+7M
GRXYs0KTG4SUdRwJOPx/4vwEXUNsUFWVYlvCAbkLwu+ugKMBxO8JlRWjPv9wgRaIiRuuVhurb4Dp
DVXUZAPMPCt/5PeDgxDFuXT/umf7z+cCSL2loRizGd1gXkEsmBTyAa9A9LM53Q0Zn3Bn+jbfVX7e
eDDbzoHa6qDwifMRzyFpeqtW3ecdZ2dmncF18aP5p8Mfe8c4Rlr6HCo+teHX8H2YYxEkrkG7OUmu
X5C7IscXAB7jKuGsbdCPqjKCGtDDEwBQrkpIz93F44akrmHR4bLMn9D2bQ0+VA3QKblK4pBgn3nu
Dw9SpDByH4Fr3FeMfKtXWta7/HZTvIe8eufZoDupypZ3MOP0n54rDgpnZBYg8AC9FkUVt+OfAh1Y
0ZMesv8Y/LMOqhBXA+ile1qkr/fltLok1f9CS8naR5216OY56ybt9bU31DFfIIM2oTUQ2xWDZ7SY
630vBB7yHCxw2tbdoMLT1VXFxu148M5SVI4boPa6DzBZcQLzv57wiMdtTrOHzVJTLFhmlrOgiKfG
UHVkJ5n7zccDry0jzQEQO9bbYFGImEFLxjYR/SUfvAv126C92oQZijBTCjq/xj0NvwC6XbYOCh+8
Jlz26u1P4Gxqfgy8uNIqljEffgye2Sp+MMh5iphE+xyqVATZ5VTvUacMgPKgNKLlyY8ZIR7LcZHQ
hx9J6AnE9cyB5Cjk2O7XZnaGHnNiT4jHIlv67BotvwuoVc7lX6k4iuNxp/SDQZy9+TO9ay/e5DAt
8UPONurYhvjTyzkATqky8FvRHmR2fU7D7ymkKa8lSMxnWJNhAx3pOc+griGGUByJVURfe0Jc/9i3
yyN3qan9U7aShFqlt9qghQgYjTpe0uY2403PSpvefPVPu4JCm3EwL6xB5J0oLudgMhptXQok91JV
RRMzAdbKWJTDFEBLHq//5sDMf2N/PZ9YD4guStdhYtuW5Xos55urvni/pBp/blC0JRPjSwPry329
q+TBDaNFDnUpT1XwfBZWdUh9thoASf6ezEWypEtPYOmYS6KZeurBiCUvdCbCbRd/mbZhGJxKEx5P
lph0BxKYQ43KZ0BnWXHSNxxhmC2bm/HlfvEOwM3WUWE5soEPoP7WYibUjfQr2VI7YA6DhuSNOhe/
bA4OFsJ9/xim5s2BugAw5f3ErKLfU4Yc4hgKqBKp2kIqNEO5P0GtDw/XePZJ//7X5eSxDGmx1EDP
DGlrobrX2kai82LHOUMGy2HNjwyYs+L4Ja/NkfxlTiyuAPZSnVX1h0F6yJv65uk9oBhDCBd5cJLJ
P2ZND2VFhCIBMfGhK+o1zO7o94oZ8YSX2htYpTFg+d48pKmqFn0vrk2VR2tP4ECQG0Yyg4f2exhb
kD4LReImFXziAt/qTRJZ0A8PqiKwG3MScHsfzP7vuSp+LrvcyDi11Bz/E9XpfdxrkDi2gfaS8FOh
2Sk43fU6rSUM1P2KtBFKkabxZjHnNjsQjwfZKWCJ3djSpqrPx6wf/xmk+2rC9kfY7H4ewuujX7GY
kHPPZrss4wThkQCoxDU1+40Gub8cZ3h/ncXzO68jcZ+pkb+FkeAcyEHkUeH3+09ZfCgYjq2Qs0Mt
h9TiP7jiDoPqHallw7zNSni4pbGGgEL2Ewyeh85kGInC5VNuvZJVoHZuZEhl/PEPUa7iY64J0orj
8kYc3uZu1iK2ULvIHQrnBA90OLokINcPtQ6y1ugkaxhqXwOmAzoDUm84Q88TEiLiNsy+MDNiZl0+
JDwkcyV2kUnPOrvTr5GdMoz/MGMZ9viY2dCrwc7r05zicHo0tywHXBqHRXTOw8iCv+bzxvYlyJHd
Ype8TTCKJpeag7iONukYNlbYrF0GqKPLDRR2NK24zSjS+eKiZOdEIhy5bYSpKn1sdPLa2qK8qZsQ
mtS/rIGqg1sKiTk0AIvUW1Ryo0+B4xfdHzQugHk3VqcK8UojmsGiOuKTVNsPmINAN3GxIBm8F4tL
U9uny1EsP+lWZaR8kRs+6taeYecWmn4pp4q9WJDwxQSOAWhOTzYNk/+tXBKCMpwzke3S0ZJVrv3V
ee52G0ivzbyxzi8lk9qNFCBDXgob+nrRu9GWeE6ocMjKzXOfoRYwg1iWnGR/Be8ikoElWwJFsTKS
kbrOKZvBUiNAs4XQ5PZPHfC35dzQ7JCNayDwYimB9L10wihDwQwdU5S4njfpcDOcovSEZxXi9n4L
C6qmgQ+vRRXZZcjXoR0BPql6cLvlPbzLUEj31gz1z0O1djQ1oHsTWRwaW09Ax0P7PlZRaJv0Hmk1
Vrjmpm53WYVMLonWtC09m6dZaWAHcowKH+ztq0DbByGhsR1DLF2fEcVNd9+LXdfWeU5+oh0AP11i
lURIBBAkJWmWpIZMTsk5JrlzOKOOKNJQKah9HiRhljUnjotXoLPKQliJFMGa/Kikjyv0tk0JGQmm
rfzSlWl7Hq2l952jdM2nfYudHkCVNRARrg5LCaemreDNItogWYDr4FAOEJRC4YwKKqjHHe6C6LTM
3HeQ6HleTAPYKhNeOFp5xCxUDqXICDBjQlbTUiTto+9XxuE/vGzSqlW+iJYaTR8BEaA8nPEvT7lu
0ZMoHpX5tVmYKVE5YmJotCie0azEAwIbhuAwZw6xIdBF0g5xwc0PxTy+qazuj7BFpvvSySsXJXpW
U1q5/DeNepLs0B9C1olI6xsxVZtMWyiJ+ccHBnDoXRJHgLVbKOdB20k/xoUA45Jb3vVi3RRKyGBt
49hb/PPcY8K7ED3MGjC5kZZq9bgnmaLCbasoZDs8ecUMXWZqeQaK7dPYkqQUfvJMl9iAy8JJCEqU
i9/LFMDqevepGK3HLDiDovTi2kliuNKlSeqPYKoGB3B29E4DX0DD+yqmuxkrtWOIH1w9T2Qrqgm+
w8xApcR3fLenmZE/Y3N7+clhbmmVoZPJl6x/H7i8uv+m5HJvvU3ag7cwzV8UjrTvyGkG6kmSPucF
EUjCjXmwL4Au95wzhcqwzs/IuwYiS0/HwetzYNWxAsGQkYTA92EYmz6GkZV8+jVXtw1HHgxES/LK
9NMgSszWIw4eDicVI4eb2Ek13oMjvwFSVci+xmKMtv8ulw9y22NuP3Qm7TqEQpthkOnRdLVzM62Z
YMJBuXkeX+3eFHJz1OHV06bDV1iW5u9+Njf6XYUzeT3N5FIYyyr9Y0e5gltpwtWt1idqx7UblsI2
KWv1uieFJ4/NRj59uizqdjTH7IIxibGFhMDtsRKKmmkzJkLtTPHqU9fagk4FR3GFTVsPlat0e/Eg
MOt2aCjOEHUDAuspAzVApIxvqdAKJ6YHp383MYKnGuiVrtpoJlbRZ5RwmdmTUppRD7eDsjSCcgDh
nNhYDVbZBhDc8K+/tDs47DEWxr1cXuF0EB2HscDr/xL2AlYC1GSCx5MVDm6nhGZWFodZEf3/FzHm
0/4JGy1gQsUUfao58MWv2kd5FdJKpA5qkfW6fdNDKH0ffkGdVgr7oL8szWzRsLHgnwDuzRD/7QQU
mDOcJWjmx0O/a8NOnlT2LU7Q/zsjGKRbpnNvIlaW6sW4KjYsI/qFC79K3aMNH0MRYBBMnPp2oOqi
8RWpIwVwYfzztbuX4Q78IwMCNkoc+HcemBI1aLq4Aj1mV7txzGxGJaRVGhwGpTc3uGs3ilMcEgFZ
TD5geCLmP88qBSw12bjgnq9uHXinEiouA4kEZlSwRilTJsdJlI1bdOkzWXqbxUwMLou/fSyahXmJ
5GxyeuidYIaBJRMR5PaAsC7pnwKGMsnnU5/BGfcjbsFB0B1MbRMFYayADpuw0TbMMPYceGMbJU/g
pAcWRyJm8BoS9QkzZMaSqZcyhdm61P0uPKHyquLu2ioIH0Ql2oSLI5JcQ5ZnnUYbw9g36h3A4obw
8+X1zk+Bqdbx9vRs8yPAj4s6Scpbkcr0oNVmP6EeFduOfXOEVY/iYyqJ7WvrgL6cVqAwxDqt1AiF
11p1pIvBqhP6yQ0abA0MI1vGL17cEwVclURf0T9dYDu7t6jUdPXQR80itZPc6sHXWMfDwHjL2jzj
6Hm62IzdsBdCgWgmz14AhDUC0Jd7eFj14324xtVFHjp7fJemBcDo46h6eBfgGQaUebUiqsa0u3TT
39kmNNBM2PTyQ+qE+EwftQPnMNXDpBy+WLA3Q5QWzmTkMTAEm9mKBtbgsIlKXvHHw1zSiEbb6lIJ
vvZIjxugJb5aVuVcrZLTknpDUwG3raOE+U5hoa6AVGFtvWs5ogDiEC5Ow8ZQiLTRYJQf+dDan9Ap
b+9cGBhqehB9rDxox8LX2+N2Z9t+VJG9zHw05fgUe5j4/ORZNo73wn8W0Qel6z/qr42u8Zoz4QuX
BHfd4r0SzliiHvlZ6dY7zre7b4v+1pcNorAbtGmB0tWiOkcwz1x16F5PDBma3oKeK+Fw2hXvH1kA
/j+FqMhIDe45p5tJe1wxzRurrm7GWQ2OQKPp/G0acaCnqNV95QdADfRlw5oNtZrfUokoEsqAA64l
JJGfLVqeOcd0Pxxa/uVFQErff2pePFneV60zeFRPaWvptDpW50Mg1EOFeAe/EwOA1XsnTRpH1lRa
A0TpGkAzusSZF1Fl+hFL1ZpcQMW5tPVpsoG0Dgau+E4nGscGXnU17LuVBF3ERc/sVewA3vx+9zhH
xqbQNHemYYC3WutPXWSOIFlRrpbNsj66WA0QAem21ku4M/3O5cp+ifepEZt5nxEdun10uUNxW/g5
EYWCSyx5o8tauRgcLNxsctwZDAxfI27IyhFueF1rNROiZILz6pCQvMc8t7QO0vDxBrLWceL4aghX
GGU7vkagXuJEDTp1+YRxkiyymNZyVOTJZaV/GEOi5SF6hbmZ7MLjOkHl4FEdc0AbhGXlcoJd/2QA
ro0KF/vBphgsMJYwYBgk6S2lbsc0NsvQSzSeV71BLqLQH3G2dtBB+X1RDyQFMNDPOBepWJ8BiNHQ
QY1kPxxwMnPpIPRAmUWvoYioCwZz//1wgk9U/RvgHZfbEruKgPXxEXRDLzaR8PMbHKwquR/Efo0Y
z+QKmbGRZ1cKxcNKAnAp63Ni00e6RoV4wscsKhRf77rqgX6JNt4AOgFAArXIzx/M0w44HPkflg2k
+OOzrbgO7CXWhFX1/PFAUzqRjhIw1BOF5BgaYkV6B8R6TYMYKKVMyaavRyXe3gVZEuO5JyNVi2lq
QUpYUcVUK4Av91rYFpi5KnrxLRsvLDKpBMQcXlSy68xkwXY3UcRS5+88MRHEYseXL9cLynRU+/2U
WjMLhaQpMvBR7cJkFsHCFNWVTfu0KYkaZLYBdnDEKr8ePI2AcBkIcrlY+7ro3k64sCRlLGPdndU9
VL+2K0gMNeD9jakCk24RXEOwPLDmp1enGeePRY02JAVroC7h2A9CqhDZWIxSsm1OXpBIVOdTZkYt
/mHrTtjVO/ufVS3bcrMKvQKedBIlDdEGy2UMRBulbaG9ibl+E4vixTQM3/htxCqYghxL+1qEvS7H
aGyEJhSOTCwvDurE+Ls8F2G5ZRWXa1vk2I9gYqEM85fYMLYdKCte5EMrY+rQ6h0aK/WRg+Q8aEXH
m1oYnF8Cim5JwUKSJizkocMTdPYkKB18EkKJHGDUEUhN4PVsBLKQwe2hgp6hK9k7aUJJBquQdfnu
CJHq+m+hYJfOP0UqjCGMzOlUtce0B/qPo3rr0HkXJVBcLoMScFCyfTZAHQg/j7KWjlNPwAYHTsm/
wiwodtGBhbwNsXbY8wdzvMyB3zSfGeZ30rUeb5t7gVU7xh0GhhZcsBGufmB8PgbSezg6AW6NySo4
8I3KHVQmhzU647GbA0Jjp7XBEJF5jZQWH3lM9ItfR6hPm3dEb4Ty9Z3gvoWvQeyjqTlnCWMldXvW
oU9yjhCIJY0kHtKDGBmi9ffTh9Ef+1uss4icxipdmtCHIR0LwywLnILB0+gfPSjb8yeulawVGKcr
5z/2gGlyiOapVMQGhiSnd2PS+ypFzmkD9nQefc9DSwVBigIP5fSrgn27Aw6LQApn3XA6o3c2tewj
geri4veyiBibAqRRGeu+sKo8tXDS0zWdG6wZYotTO3J35b2TIISV9jAHO+L8Mhn+HxzCdNMcsbzH
jLVSKkSvFEtM+uhTfC4qqOpr8+ebsrZhHvyg/V7ZTGnZ1MxpaiIOH4rrbKUZptDBOueFg8fXDhB8
xqoCrEY459N8UHm3/EbNOVL3ZfjBgB8yVKm3r05FPGmQWx/lTmP7xIFP/3w0iWsFmB/Q2iLhQRA4
NfojHof2rWJ6rTJv3ZRh5SuEj9KBNURtuViCa02hWy9xJvfBsAocEd2p3AK/F2n3SC/EaGLVCo93
ndkadVSDK2OJMNuTXl87et9v7XleA8hmlKE2tR3W2aeV/Q5sXcF2rcb+hEA39lFQZd4IRZGRRz+h
Db0G/4PjLAbu/i7OJ+oCMVdT+Soe8I/vr/Bx32OYFomk1h/p0CSnIQK17OM1s7LhPnvHg+qAQwNO
nBcGVGee84qLepMAFaatLFuCuF2UzSLh/jnDe/UwQUGS8bq+QSrWqKAUTdWQ+MExsWPYvphxZ9d1
FKK4b2DOaS1Yr3i5RiLMVqA3v/kZ9/etd2mrhJPQckF0gepKuIRc7RmBczDKAY7x9HXCxyRBNKjO
JFRt9/fv/eEySC1OmOQ9rJlkzyLms6OgvvrDnXHL7ASGLp6DRd3GM1ZTjS1d8rh+NkSJr6p4K9mF
RrquAaZ2qkyFU8V0vTrX7QoH2V+/bbVQ1ne/uM+vTINKXwWdft4Zk+o95L5ybnBhGh/0laSHgX99
WniMMAbG1+REkTdHEzNQsyXZHiHOaJr+cMRm4RIlYVf4F+n09aJO3+QfgRkAo+CR+i9tfEt0FOYi
s3lY2Mw2FaO+wljO32T/tbdCMYx04FZMfU8obGJOIIExQ6M+0DjF3mahHzDrpw60gZE+PdH7IxO/
wRT+dc9O/wc5hAr665ptYekvd6uywwAyFiORE3Aa6GkwVHMsnr+AUUSVGEKqAwO4AWVzBadyhenu
mR0awruoeXT6CYPlcX/klrq/WRRi+p0rBpfU4vnWDA+QVHLlvxv3fI7IlMrclKizC1LUXeFoAb6o
Pwivi67s2NEp74/0lYH1+amE5rM/yx1i69M9uS8rJh6IFgFmz6e35OCQMWOaGR7TejXHUUiJ+AC5
K1A/5XMBAlufIxaDG+2eW6bUR2B5XYRNn4k9N2Oj+18ofjz9Mf5cJCVWdOefAdRwmC8ZPWpQhUFr
VOf3b0TdK0Ns6sIskPpUs9n/M/0jLStiQ1J4S+Tn4NL+44wYr3TCCwxBevfIiVNaXIqFiXBsBZHt
uQ1zQy1VDGEChuD9WHIkBz8vDSZU9VpTXRNWMhbUP7gz7Wv07TsVeYTqExb6/5tPrRU37SAZlOG3
S0jACOVOUzWaUGeV7i+zgOCa0W6F+Hrt/xyAaXyK/PiQdsOnRxhjhKcV5r+jXfpGUGKCdob7NxfZ
r73mK8Me1YljZpIXpHfujZAPcHB77xleh11gLKpw44S3cX0FFPIIeg7/I+LaSuSdttiKI22+5TNk
tw0J9c3inqihxHtLeUjVci+0S7R+J/WOJtS2NgirtQZXXimKWe8H/Josx3jPl99V8DTE7/g35W/Z
28ekWkh1PM0zBC9Lb97BDewbat9mKycuShuE11Pe2fFmLEO/2QZUzeJiCs7UUjca7W3K1S9cVV3c
xx7jifxB9UKIYiERqafUU3ROAWaU/tZID66W1a6NaGR422k3Dd9LpJC8GB23oVjtdjBWR83bpIGT
bkDwqQS6iQuzz6VOJrQPWcEjZ1XjfY08SUFfHtFiLSXZa7cehqo2Ncj8ulZa4r/eM3DgeGT8JPzI
boalToIOFpldsNNIqN5L1Mxs4FUqt64T4PsOOmZ7EarpAF5DW3/SaDsnHe3S+pHfoneA64yCzwqb
tCOpf1q5SWXb4pnP0J41ZcUunsWAN6Borv3g+EBw/JNdjzDEWhMa5FgeF+ueRFoJ4bf5Ary/1XZq
gzuUiISQ9/yOIBrPxgDM8/5O6byniQBQqZ3MIEWSue6EZZ9B47Vjr8lqtMTkuGLkaKntNL4GmcH9
eF3imQgtOsJDOKYkTW/cPWY3VfKmNAatP2O2u0I6z6hy94Oqrfiiz6E7jenP3RpkzyGSV3mx6e2P
wixprKlP7z3tUCZfCVwlTTkypMu7tJVbZAcdxbTPHr99BBOKGZl/0OMNYQopQQeqOPo3I43No0jS
BHmhsXPPSd8bSP7Q4l6z30QNieZ7yM5Ri1mgbnl/nS9F6B2vZa/qvEVAh0I10tYGmIRDCKkKzfNt
wpdWIH19T0jEqCkGpTlDIt6yncpSErAbEmPK2ak2TQwxxF5JFcqB3SpD5Ny/bDKpRnkZQsUKUw7T
bvFhs2YNBB+fZljXpVVFIvDdlA0MadmNa7nDJwssDHXQc6PMJbQIzxeEM3Pb/X8PVH3rXBy/xn5n
mhNP/RaI3mKk+neVfMDVB/KttB9+hcebQPzKfJAjypn2jhuTa3igqhywBeDEPGTQZvgVPo32pr/s
wI/Hs8ORwPY5XnLahiiLu5TDkxz/zP+AW989OtvjV0MW/LY0i8TcdGZXWgplTTB6w+E//SENVTef
CIyxeWi6ahinAOeoI+aHWoix25fi7SjWznAl5axD4lSBHxNtePrk9AY8iaW1Vjv/srWpvTUbPZhI
vbaP5ElMsDhq/ziB70dnAyNQ7SHncKWWVEkdpa4uX2NVsmldSn400bX3iWzyDY7jgVUPNT2w5T9/
jsN7+MoOjE0xMp7aKOa3jPdDzQyb/aiOlmU7swNkwsM91zaDAwY8EmEVBgFnKnJOt1aAlnRjq4E9
gYWob4Ut26fYDBei1uohdJT/QGWVeLoVKHm6LGmsPDw6KJDmXppaK0r8QCHCANbdehmNEpW/NU5q
pZvh+YnOOfCSM+Qeb9AowRbQWER6eglAE3U0OZ5uQTkIIWLiUYyBlVeyByfktymhRoV8SYn917A9
/fU6qXfJw6sDlRzww/r9d/DO1pc/IcGeE03QmfWYryy7N9wA8wTV48UlA7qTKT9Geg9qLHHoQ9fE
VbF7SQPqfZPoAcrYHBmD4C/XewBDU5j0s6129/gN/EL6WmKgj5d2lWXj93j0Kq52sntQMC9PC0Mm
QnAGrioSxOLdz2gg5aZahyBBZgNueHjiuPtcnooh+cS5tEy2mDpmfqJloB3IuPgK15ypZH2cTIEn
YByxmA2WmjKOV/FmO8WVBfFy+3446UbcUzPXH+5intN1gOAABwykVBPysWZOsOKA1SXi025KyOCF
wzE7dD713s4o6XBQZLJVcVjUMbg1CGLbC9Jl3vRmos8wUDZbQVtKnq+vdGgCCH0JYEs/wlcNkFhY
+Ea7f7Sr3GIfL0pg250t0Z8kXa58fVjbYEcwyjnXaNl2+Vhnuek7IVtgDBNa5UkEjhxcwU4Jk0KX
ZwofDxNpFhAHlYcOftUJ0BrlEvwHq0qUhR/sNRAI7r/Z4vkej5R/6S+IEBaXdgOV3mXZLp0sGqGX
JMvMixE43ONq7K9QtNH+LRyn85T2B+3G27MC1/kuh2A0kimVAC5Jmj7bzp1abc7CC1F3bri7Q0xh
RaI1OaPDk0AVqVS2Z9myTOUnE5UuXSV6LvrjXooKMScjGugAXmxrrd8krGMfwNcfke60nADz9Hta
K1F1GdpTi/YkMmGNnlAEqfdVx+yrQUHURxu9Q2hJwQ3tz5ecvQN1BNs5D8dYYD0FuQBxVZ8chnfK
bI15GKtfw6aPaE2mFNnO9ShlbNKKK9JD0y4E/Q3iIMSzdpamoF6ik+KAxmyUs6BRMkLbTb4+TLCI
HL/8j7/Q1pJ3ze0lVVW8yEmwO4GwlJvubueguv4EtajypZuGNhAAzy8E18PFVDqo+8WHlEah1p4X
yJYqsSFTQUzM/Y3qg22bSgBtl4pkWS7LpsX17wOOIP6B/V9C/hqcELATClrdelWmORtyvYvO9+v6
QJrrpGy17y4N5NEpNnB6WOhIjHLnPb2sd6OcBuuyzuYHao01KCuMACkkO1RbrSpA7homgYF6AUO9
9HEqIGvt4qLofYtIrUEfoRfP4KTdkaFVESugWJ024XCZ2PHtYk0gVhYEgSaqePlj6nLMzfI3PecV
oiSzAj/XOjeOFFxMP9gyOHGT31dYMIgeSQogmlZW8jw0w8rg04UTMkrm7fZpiy8iyGYVgoddVWVL
/wr4VjRlMhAqsPO/lHpLk1b6565xyDOjsb3rcHDq84CYVOBigrwsdDVtKiEkCZcolUXjCmNFFrpj
WsoF4OxQf28HXn92fXjSwae5/NYdYM2qt9pno63jbBzAshmmwGDo9ZUEuLB+xX8QBnTpnDnHh9qA
P79u09hmln+gmy0HIJtTF13OSnonzRrHXMY72XMobBjNdb2CbiKEaoZHlxxgb5PPt7pZ65j/Wlqa
2KShUqWmqmxqpW8UUjIL1uzV0aAQCYcBbMO2rBffeZOCz3+rm9w9tpuMZqxrpZUbJEeEuvmg5sZY
qeilkBvqcuD+xp1o6lhtUq/gf0ZYKe08xb+7oBEVXwF+vEZLNz6ndk6bWZG7u9U405eQbFr285C7
vNsvAX6DbCeVlyT0RzqnJs5L2uyqfjucufN3t75YaMzkpRyazJcIWXDlXUSXvIZJWJoWJryXNnr+
SU5D+7iIAGMs0wsncxR5M94LALRNHdxcO4KAPMdljBncW524NOTqF5rEgw/m+2+9h3Y2TRiXq5FQ
Bhppm2E/GW4IJRANDp9qXQHDLyOLcR2QB0nEGKQCu2PM676bvHUD9wRf+ZEjH+gwSx2l2v2SNqGp
gIoGGSXRKDznQ0Q3axt+ULAzqvUik+Fyi+vXH23/OztdqlGRJSnm3XPraX/7b2S6FO2EWkakvqIL
hSxFb5OvB/ZfwJ74Qzk+KSVBl+YcGpGLIggeXg7Fy7RqmKCO+S4hcddlXi7fGRqpVdbOBsBWAQsX
1Vmmp6j2eTLGpEPGUTNnd8WEosTi+wUR68BYjwP8FXUNhYBXC2GIAgkiAuBjxXuGo6CxDqsKRqOC
kUmUrxoYGBU/JW5gtf8sTgNrfvIOGSQ9tv2HdZjvxNnunv5dYneb0Ty3zWnrHUCLjjGYsDt8SwhD
eYu6NScg3pF0Zo2v3tcMOM956oXgSX3WtTrAJNtFwFlZ55SaeW1CNVS/wv1Ev375vX+Ap05F8a4d
vUPGtXu+fMx5oVRjAEcFxSgoy1jd8P2LHtB00GJqz9JWB7k5M/Bfj4eFbKoFPjLNd+Hp+Xau1D4f
9UFWSqaoj2XyU/3SgEAmPCimkuqblfFsDCiH3RnoSTkyOKJXIlKm2CJb2L+pT8XffxobD3J/XWc/
HnG52P9OhoP36JcEbHpVJ1QvOeww16lQiI5B4qFbyZzT8al2bBZt8or9a7/y6rnve3HfgiQvGFtQ
Eg35n4GX5/uVlUbuwyBMmTo+p/jXWKJqpXVbyZ7WsITLKPL/slzQ0+47S8Vkfy8fLIfAu5R8gMCZ
6ipWGJRrxXRh2HJReyKyQM8GYcL/lqQd9vV9Th53s47V47uLdVp/sYB5q7r/NyMYI6xoApYdbgXs
Seqd41MEN8dqI3IHKvJwhzAvncfJLcG/fyIvCN2RU0VPlPeMHfNYwJHBAoNe9bKY2/11QjD3SKnV
3wVWhivi/awWduimTZ1fTilLmJkK9leY+E7M7ir4EF/Lj4zGi0ZhPWB1/fNsUmnSOeA8d++xIC3J
7H9Ccfu7tpPF6bxsBqJaJxsBtI6m8b33cEL0ri5SX0LcBa+q8R0I7sApvAusH1q0TVqjJ43WI15D
jtXtuiMo2OzEvjflLXfi24EZFDcpqVBm50Dv71l3JvImjpq0JJhcoS9D7TLbjBtCsLpOAnqqWX8Z
braFYF73un0+VXCRLzkzqEhvKKqWmgN/AGA7czf84rFtXs+fzExVGB/65oEH36kJA3mio/ShPsgv
Z8+NmriZemy+M1AhiTHNZHMTA1u4L3hNJNrkNBaAQYrthSzQk5KycC5EhrWL3M6Ros9SGnZtTLoz
SqMzN1Xlh9CTD+YbHaYQU1i4paYmLx9OCRjZiBkjSUpc4ECwGbJC5LMZVR4rukhbwdkjpV8EEdoG
sBipq6W1bxlabL6d+akb7Ruy6kG5t/Da0G5YZUFLIL/hBldVkpx6X0B/DcBMRMBGlpE26oM+6CoP
if7WVJECljmf9tnOYMtOeH8GJoxxzP1joLifjjyD5s+ilh5LMy9WGPRJSgBwYvntCACwD+hTlvcq
9K0+BGwQJbQXeP934wT1eNGBoUHvpgfZm/9zsDnWZfGiGUxxAQy7MBE5b8go/dZLsfFuife2eozh
tsNKzN9pgrrZYQt6hQi+h+cV6VWOapwvQrGvAdAKGZUrfXT6jpZfHPGG6Nd6FkEJ/2TzT1JV6Hm8
gq4Jmx+w+76y8GUc7jqetfxsPlTL9SkLFaBd9ZmV0T4H6V097tAX41US1gadTQkgI0XdWan4RAj2
ZwfBMM/Kn6wbHfe7qoSckeaB0Y5RR0gx1WvinqH+F7ZLg92R9hwdC59KzA7Hn+wrs6p6jorFFK8/
KZgxvnJZmoQh8K7rdBjNkbsmjTBTNTsMxCIvt+6eoJJdUlFOMNmf88c3Z3omSGhqmV8AoHcAmlBF
ricmSoTlR+WSOVnvaj52B75cYTpiHZIdCYMwFN/6ZvQFKK1VyRaz/jy2r8YznQpzelZzL33EjOZj
8mVdNePTb6NPn/8KXZL1Z5FYSKzQsuDYX/Kfx4/t/VifjNEAm384/HDj/0/uP7zjXiV96pVXN5vU
DXNpn+Q1JDTdsP3eYOasPkK8AbvLAAk0HhLSRg5J1zJ54NAHctCEg/d8Fggvuh7QfcN1bDkYC99j
mmyX5SfwU9qFc6ki2TU838YqmCJ8gDNyKpRzAy08ya41CkRQhu2788NlTlAu2MEG5eTQFEJiKX4j
5hVfa6uVKL1pRZ9op9PwDk+Wt0yFAAhh2DZ0m8tRpS3STotO7OGXefs88537bd5h1GTrnsrZ00jQ
0IpBXXv5FKS+0iMMY3z2x5QOqR1DDjQcuqkoqKtmSUxtnk8yEkZJ0Lo2v70kRRqDXn230ZmzXGDF
L0vhYOIJ9cH5FHcvqgq0MYjq+NxnTLuSOB5umPqjDuQ5oK7IioBsnbrqEYgYgQpQ5ZSRCkurcpgN
R5r7CcFtdhpiVzoU257dPwCypM9rOPf+sG9ysKaiFa2D29zT+QX6TgLh6UacOij/hJh1qLw95z+b
dVtUSN8DbRO/sWdr3dKEzVOgarfiX54yH1c7xrAqRgvcilMDSjpktvktc5m+jWR0Yls32RHuhkre
00qJo8mJEVtrv5s5pKBQ+Cn/QY8kmVaf6dCfMLvBXgVh++1xqam8iJPPLkCy+Shf6bzejduoci7a
/Jexyu3Pd2BhGhA0WisnW2KZUrRqRaT0rEz16uKBIxvMsTLrrQTS3nYB9Kx9oC8zdnaTy8ByLcpi
KZWHYF4Q8StIYX9f/eoBWsmr9bFPMe9HxILWItBi4A/wEOQfqmZdqjsJZ3SW/MOC7544b+0RhQNt
I8/iC0I6Y1xtxPw9AQFr42smtGdkWXzutkSx7dbOrL3whOMqNqgNwnGJVosYSiGMxue78QmxaQ5A
AM6Rub/AQHU7ufkABs/DzEiT3PQacXHjWc4u5MNegMOisv0VgsSmVOhCNyeouTiRtoRVB+S+17Ns
v4AGsXfv7+cvM/9my25K0qNEXZe/JnDM6VjF/3/6HYgbvGr0BKUd2Lzirv7QtBunxQO6Hd2YDM/9
Y8MWhmY6PMva3kPkBOI6j69fq76bQvPRPCGvoWfVsg2ciTaqlUYBkt5AvT8x9iZRh7P+u963T66k
6Z3D1ww5nEO/0hvC1MP/k+70tIha06vPgkA9kmDPwTj9dgeULDWihY621LmIRVkOYQAJ2PkbhC4V
18DsOaP8gVr/k7YLYiSlIMYzhp7qiB0qRcjD9bFjJLRX/mfmTG2EhoGxJgXdQAD2C08ODXJMNReG
QWCTa676XHD2B/tSpEE5CuKCh7JHPInnLoga0Jle91Tmjtmtq23RcDACwkSwJkvI9f8zNpsg0LCz
SdLbj80+TDnEekR/NInqbRVwMjWVFVkn1XLmb8lbWCiWU9/GwtX/02NNQYw/5dxCl+lxlXyqhxoy
r3OLlTfj4+FXK7Il3o9NDDad9cLMTKZo5teRhd7ImI2/L3aJmClfTBaO1h2FZPQyVv1+Eh2IaB9g
8ZtOZbhUb4swRJQF+hll6NzGG94Jgcl7AJPOmcY5QBw6xlYVMEkmC2IOC25gJdipTtxu2X5zIu3u
VXpXrg9/5yX0eNFh7MAKTiNUqNhpce3nQLOHXF97PyZveG6PJdQ8v4/SIgE3rIN5MY7L5COyQ1H9
jgK2U05IEt1mgRbg49mVMTBC+qot6AtSoW54AkObuHedNKa+C/K/tDt7bzXn3VffKLNLr/pwdzk9
qvxSV/bQRMIEavpL/MpuNFxj6j+eUGtKC2xb+RRGlzY82b1oKirLJIsRCmHzXfgq+nujFX7CrznI
6fenTwG6+aiKcuBJV2Sc6nVnlKidpTx1c6QsCoYX+Gtl9xLRQSTcV/N3Tow5bqXdrglK0Wtpz5LT
80aSdpnv8GKD4pDlEriPAW4HlvuAVrPOYKTnLsInZ45WA9DnIW2PrqakkRglD6fjdvU2V4pve2ns
MF8DfntnE3g1U7po/9M1SLVCEJGHkhxBbljv8mi2LS6lVghbejhfXvVEh8QIDsQ6B/nRaZE/9t0x
Y9f3rH6K6VztiFJLNTsd5w87YBy7ZifIsbVn9g9qtGJwLoIghoDGGITqDATxt4iijtzGkUct+fKf
ToSgT6mOEHJa6ZVx57Vi+4W4uQPGA+WS7vgVVhgnm41HDwpWIBNfuetzr+VrUF1tkfBMZcpIXyC5
hJgrnPeg5zuah+BE5Nns1tguTp9XIva++AdaJ+qDgpD7JZurSG2SWkAHTUb51jtlIe9JZb6RMy0Y
FGy5Xt/Li8ywlqSw2Q1HxhJxhOCQ06H4S/wITsCImZBrzRmN/0aOONHIcA1LdgKU7RyjVhepUO9T
h2bQuEdzKdZkeJLpGe3pa1xlDBlUF1OO5EDPjuMYR8tJxKjcBHwgxnrv9in96fFCBQi6bp5eApmq
txlUQH/je5HXg4nSgjLjNQ2q5E1ZGGwL3LaYfTOnf5VODYRdN6Oe+bVlg2UV2xu3iE5D0hKUvhRy
8Tsb+Apl7t9X+jmCo2Q1P3ETNXl/lPof0hD30knIdVplIe4On/lE4polDw023HAj6j6ZPHvD8Uma
McLMfHe6PZ1G2Qdvy2tGFLiTqBUYXsSk7vR3ttRxdJSN0Ygtto+9+Pyh6WBdBmXId5YuG3hH7hsg
3mHdXLJvTCSIvunQ3kF6mD5f5y3l5xhyE+4aWzTcfdULBwwHWXEktMqy/inKUKfy9LT00XmH7Z0G
f3ixh/kke1iaGe3zw2klZrkX66pQb1S+Rp+iS7vKAdEB13z4dxCckGnLXSAOS57eNjZ6iT1fXLwz
x3RAxvoiMf/pBDrrMHigYw4r7YnoPCIM9xJR7cOR9/0agvpdwbLOzeHN5ucJJq5mSfJWDU5k8ZYT
pFjr5lgGnzecVDOuVfqGgFO3rhwxcQpjQ5G0ioxQfGI3qTTpQhRQ5m1cbhRS+aFUjE6P5awlNC63
KvEamskz+8hBBCxI+z9lQtI1yd82z3c1WiTG96hLODbnDAqUWXuZXtG8qaZRhNVZLD8/N/TUltnu
YVEZE5gEu81XBI1/G3ow6gip0HREWifJlEA42mWtyPqzA6QWq6ScUwWaz5KNs6BV6kfYbI+5jdaO
nWzGmMkOXaT03n154Zg+JboWgoJfGlz3RP5NlGFRaNAY5APiWgsGGv3x0jg6xrybu7YEgddnOnyi
XSCdbLqsRT0WyZtUDmc8L24SQtnZuese+AwskRIKtDXnmeZ/VyeO+p9zvGYUzWs4E79F7gB4NI4c
nUE/6O5Ws69T3jwyPa8rCjUOuRhp7FmI5ePxAcSPT+PKrebFgfPQ3hlUEX6VdbsqtaU55cHToHM3
ZBl1WoMPTSGammSqaqKveXekxglE5VQajb4Ho/cuChhkQ5EtP7nVmF3nrau852W3YbUV+KhLtAzE
doCp1NLB7L3R5jlCE1hQHF9Y+ehnso+TCD/EO3QHkHKV5zNB5bb3HThYMxfrKJj0rqgtsbCaLIE3
m9HbPLNuXUKkN8ejsm0zBWitDJyTBTKpvo0QpVrR2Hu+kr+F9H9jcdUw1/DNWwvvJpfKE2IS62sC
62fuHt++zNU93duW049ZotsXrieJVxhhESEUl370EWEmoz41LWrUIa4h+nmanz1x1eE1qkolgaUp
Yq8LpFhG/hevfA2EyBvqy2atmO56VK9d+ABff5Sk7KWp0dXucCBqOoHQVLULYeIUjy+g1aOkdZvY
UFC3e5fNBKakiOHQqgfNzE00enrgwCHMfkqckdNAj0EHqshKivr8ah7Kikyo32PCW/TEsfBfKl8+
mwLoaUcgv9fi1bpjGrUQDoEChydj7PZ7WLD8ANfGcJmh5X2ivJPEeMVry5cc6ZpJNFfTKYfpaHaz
cQN2iqpWcWV+m8eQ1PFa8KUl9gsyO+1xQ34MliJYih2y/fWaAz7DAFzH4VCMFxgJinJJQ8t1Y/cL
0nAeNx9vb3RCpJXy7tcXlUNxx8Po7DHVwS1utzDKSMcvBRMhnShFkogA8GWEiCuoIMRI750cqx4t
MRqOstpSUc6doK+LpZrfXDv9Iec4rULGursSFXxVMAOKduoxDaNqOtnHkFMaSHqFOomN+zACITEo
a/3Fydsgqai8RXmijyehQLYKKD2SWeqO9dbA7HR3PPfAuWeG08giNboNFevBrrqF9lvKO+bMm0cp
PFNAK8S9YGmy8KJS/OBZeZXUgLQ4V8pM/uzsGTGSqOeovIP6w1m7z3j16J92ZyLJYudoXf4wZ+kQ
TfE60Q5kzCrV86ppBFYpKCXJqZQ7vRwp9ZKPrtRKyDOhtlNBE9v4H9WuQNHkz6QckXVYbrUW+iFJ
gehQrVRkMqQZ3ksGAapq5p36L7C8wS6dVxGDBOiDQRBNnfg3pqbNluVCQs6yHDfaWrripbbKX+g+
P7FQItZ9Dg7PJmeFjHhhR4RKBB7Xt3EjcGb/Vn/Fy9F4CFt6czlifz3T3u6Q3yllppHj5B7fv92S
SQvEVf1NikVNROzHvkkQGSR2rcVvTQOh97qXlte8+ADZY4zkXmz2cqAZ+CuX8mfe1T5+HSwOlg/j
KrexIyuDi+q4NQtLVDXtIURNb+CHK9xvi10BqHlx/+Uk9FK9bfgP7SqehYouqQPr8/aJfBxZijtR
yHqhuyq+a5zltLC4NdFub4V754ADuG4HnKfeVyZhy3IpY2wj3im+RRu7zEnPzbfJ3xvi7ahuoIgg
KRnmktmUQqvI+Fu0HjZVc4b5HkdCpX+qXzPWyuAbWN9croqVhSP5qeJ7/obIjsgrBjXA31KbYG13
x+kWCLibn5cm5C5apvNanBDOFXotwqejBFJSAH6YdP0r8UXB+1CheHo+mGQEwJtrNkxOk5ys9suL
o0NG3ZByRPmEpYfVOY65eW1bDazjfdyiCsuYhjHTeDgn1WLNYYwrlR/gWXN49ZAwFM+jM3SX847j
NPKb35e43oPQKYaaq9ebVvJc4ZGunALuOmLBifja93RuW9ymfdokKP8bAfO7R0DdSaJFmOKrd0YI
Wdd9Psg2OpOqwtNN+oHgMgdJ8f2n94u/SA5/+z4s/JWNw4+Vwu+9jDzaU0X4fuffUDp6mo3EVrV8
5jU+6mfOS3Xnba+tX56hZFXa/wHpgjdkuninOh5of1KxXiJAPhoJoTqMYJeIVm1hXIIznMQ6TtzH
CpAbYYvevSPVhbrf3K/EG/FrmxRRGt41+89Y7UYGy0R1VDKLxvFBJxgk6j1uXtJhkJJBN8wsaMeu
skHHU/UOs01J7qTpb0i4+/c6o2egz9nH5RbXo8ZZgu7abEOQQ3Ua8P/iovfhXysyJcNIhXtNXc73
YMCqQ9vHX4MmkUcGKtxwNGcxm4POiyM8TPqZ5O5NIRX2wdzpQ2sAADL2Wor/kgjwYnVjTV++ddsz
+v2JGsOxsiYp5wTYbW6eVfR4nzKaRk19W6v4R5PEORLTDFxnewcwFQCPbjmsC24/1TFCvUgEZQ3W
yVVemvCd5/t/6xINnaUYpExmelfEihvdr3NWLbwAjtNrLOGGqnS0KkH+rJw/6JttfF2RAWX6unKW
Pa/M6Y9LbzpnTdkiU0A9PbfHW/gRDmE8U+AC1R10bRx7FBJXy2vxhHK0+8wzsxk7xUY3He+YMofw
/yX901OcjTq5Z3+UCf+Q/I6Ogo4Ijc5GfnGlc8kJ2g4xZb8ezL+p3sFBPFx1SFDKu45U+WTxevBn
jEonOttmkQA04Y+jPwEossFye2xuXt5996rE/KV8pstvI2siWXMk4GkhxC/LgMnBu15KGd/W2plc
+150AVvpQk8TITzW6zUqFXrQgcBhNWtpHoHO01WHtvVS6lWLSIq4k/EvAJHvxwTkT0e7ofxy3Niw
YDrlsJNiOWlLTAu01FHdwhBq76pkPEGLk9OnxRCuvkX8yVA0usBUu2P4VynGYl5Ekvn2QSjr2SsF
mrCDSnCyAetJ13lqGl+SZR8iXqV9mo/AQ2Vm25eZFHMO32YqKh7ZumhLIroFDSTqH66ypMI+9ViW
2sGu7vLa+iO39DFCHPXZv3ur04kd2ENAzS8piP1xV3zHVERvLgtTe6bJRpfWSM7uJZw1N6cQBSO7
YpcHdGwruMRsQjZEe6XlECzAZRJs/PkNP30+QpV6gWGWeQ9DKJfGtSoqJhaQ7smpHtMroHi47M/m
avY0KCLUPPOyfKcp5WeYjPQ16IlOSMau2jxLqi957aQ+VdaFGwati+irB8nTxt0DLTj1iF4NNEjs
9163RQio2Cxw2SAxEOjG9dF0BUr+KVELmmJSnsiJt9QXNXbMJzmDBm2+/2ynF4mE5GnPS+AtPGRE
tqc/G8WICvtqfdjLwk1TqOSwIQ7aLV+s5iIMDRFihpN9TQ0MXmzb5Yz3aPqCOzMgCfAa/YIrrCp3
g0G++d8ZF5X5LGKHNAzrPIOpYF5f3ezad9yArJo+lNol6mf4OBNIRdjZLWkNHJO3tjZfEL8vNexw
7O+rpGwoioqN++ES0djR+0xEpBFPZZIWVCv/6hs0AbyOreB+Pi8eCuCEIiaSocvSZuOKIlMgrbXC
kM0UdIEla8ViJ1emzvRtB2pIkZm9Gvb5fz+jhcUa+XKYP9Kcas94c7I4dYHeGeKitoKv0aYa0DKJ
udgW07oJHsL7AJhwYyBN2MeeODYQLCG56DU0ltthB6uSbEqqXWRO6hy7diicH65YHRZ7mewyw+Qs
tfw475w8p/IdhhMLI3In2hqF21pT9+zvPfZiVB/PRjyqMvt50Vy2G7aT77OTwDA80Xgx04vwHWZx
7Rn3MYSU16xtjel/msiEHy1GfVj2fvFXFMpPOREs4rJlMv+67d/VZuycgBTjmGQpnWSRzlTrwhPh
OHHTdOzXHIikxzOynsl/hIJJkVNaV7lZ6V1rJuoovgjrkjHQjXjgqgOkAr8H3pbeDsZkcEnbae9O
Hji+IcC1e+BNU9Xu1QmLeNxu2Q+sfyawEQOuQdbt70Ll+7VLZkdcc5vm5OBzt9+K0zHynk1iPhVe
J9H4my5jfnEGKrOBdqX8Rrsq12Pulz0qCs6FTLN+d3dunHJT5/clZ7Ks7Zk6UvkO2aX+cx/vplI2
7Tsq0jZ3Q3MKACO/M1dWrp1/wJntlIPDyX41wyypprYCdWPqEvTykYuVoFGxxeO1z7mMy/sMHk3u
GDLi1efMSjo5FJDObGwoKpBZKMHD0apiKnXxjD6GT/5taVBvOcxkiPuDI0z84g+VpAMY8ndAw0BA
LspXnDHLUN7yXyC6sn1dLJqGOsoqoC/3+FhBZv7jMxXBBY76GIN9TtnzS041BxbjuQKg3hFhjrh3
pd01wbcLPivwmBFw5bh6OMG/dY05oRbAvOZsDXwLcZk0MNYxEUFq1rWQ3X2+pKfwFsTLihGZBp3N
QAeXEROo2CIlv8SX168APtX/LOpgZZZn5d69pdTiyOt/xMqXhiM7eCYd9DKBCIAr26SVaFYrZ5FE
DjokFSgu360GxXWOaNLedlcTaumZe0DsMjQIzmavyCR+y+KLGb1phgloaS0S20InAZxV7EVlxxDv
uk7NDe0/EEBpW8K2DqbS0Mh6C0na723OqvmAZXaLIgIlcQSR77h7UBsiipMTZw3iy6aBCACHFsHF
ounAWNsw2Rf19xvddODgjnj5R6fSgm/MojqpGVuLONZ5x8ohM3szYqVw3W03CBetDqwhqgcqXKhr
GbHb310JFPuibXnH+/Kp4+zCIVdC7JYJ9r1QSZFOILqttpc0ILoAOwWFxUnE1VQI8LkgI5/Ud5oJ
IDjyEpgWp29t08kVJOfOakGXz9fdLBt+Hv46hBNgFwTTbGMEMdlvRHUFS3kXQ3Na6sJQpq17FqGW
hcp+SGvWVhJu5P35z9Z73NbZ/RpvTXXVffewSQmtBOMTlx/OgKIcIqgeHnTIQIMJsY2Tu9IWqlKx
73ImDFXPIsNdhz1lbwQP82+RhbzmQNfcph8LqUzGtaHXl9Nivs5MlcImy94oXLFvXWTfy9HW9xdd
4O1VUpNqhJLC07lZz+4zafSXXZv6ycbFFA10WGzzc/yHZLRcq9ZLcDywRLMA7nP+gnwYluWdYpne
1reW5JWu7YdRi69Xq2LsxRcr2LviLoY0iRDClmsE2ZWRah0K0OY3VdJwf57k/6r6LXUPeBba9NIG
iux6gexXuxzJ4+Ol9Zcyj9ze2LhhzKbHThUu7U9oxGZBkLoiCR9nW/oL6ecI09mq64Muw1nggQBq
TE7t3GfRtQno2BJhOkMOGzmniGlZS7IIFG+k/bf1TiMfkrDRj+NRRbWiY++XJTBzPPF9O18p8zDg
HsgQtaiWvXYdN5bhIaclYuBJ4q2w7bMnQdVRxz+In6GPqY0akZmZUJtonWTQbR5CbofDABzxpbuu
QQ/4Iu2qxZBKJNNs+HGcPHKicEtrRry2HzaAtgelb1Z+rj7tU5tNOAul//RzqrFg1utEN/syqWSb
Mcs+oVOUqju+d2YaiecocnXTsPNpAsHdMWLZC25N4VLl2OIRIOQm2FcSgXLzx0WM4SCSqdVGl9xv
fHp/8KzVpy/U04pEgrQrzifF3GDAS+IdI6zM6TCZnkULMdyku0R1ZnnRTYGSD6/3s5KeTVMg14X9
hvJu4Vbis8qchjilak1zFvKhdOq7zfIeEgJOaQuD2/+YLYG+u/XhoGjTcN2mIFEwnzBc9I8B3JEY
G4rr6Al7jze3wCd8ZZ4hAerX84WlvpWOUxRwIRpShdTK1izeCX/+bgQOyZL7vrFtruxJAoV6HDjs
SzW1wGHiwateugm/ikbmhx5GYMB8CRhOBjx+TYZdKwKTgBKeoZu5jgW50I5z/yfVErhuKSbhx5p+
N+lnEQWvnvEOjRQoFIh2wieXx3P72kTmpuoFtfIw8vXqw1xuYOWWKGgx1SbeQ+GP0h7shQ3fL7Gt
Iz/9u0VkTj6MDNlIMPL7J+/TSeZ+58mlPgv2pSQj81AbMojumEJP2c3PTZXNV33TFmggAlor9DK5
nmHvYxVOFnnd0Da9bNqd8mbZ2RX/KgbwAcFd/6MmHN1tl/Efl+Z69fmNtHrEZ2ASY/YkGVo0sp3w
Gpo65Dp8pj3cjtBDHpctmv+LRmy+YlMG1rFDJCFVhC7b0LYM84MhjLaFZjE+MayNHaxcsZbdZMVK
Xc1qbBSGc2zsqwGiDU1iKn2il/AApoY0gZCc3eXnuxv70D7e6jGWrQNbGJCeTXnX8ISGR0mY9RjS
BHcGeFh855mSxSw1yJ5AayHwcevn/rUB5YV8VNnTuUmhmndgh3RyDOK4f1z+CtfrpxPMcsJzxAIW
Mnk28iNfJnE1uZig2nsmGHqEldyl4HNu+OaXMhg3hI/7V5T9Sa+MiIxE2I/44pbP1SlLBA1T2MzE
durzXie7NMpxNagmFvauQJwYI8ioABfXqMJd2RDeNNVkpErhJnZf9btb6V0WXKqjDPasHb5K7WB+
vp9dAgSOvD4axfJseWOyZB3vdrISmp4vDES2Jg1IUPT5FQR/gHGRvkLA5VzzJjqujt6tvSBd9e7s
mzvhhrZonOUkAoQ/U9PdR8IDz5yqIrjToFnLK0i0u+8lfCGiCxTUkxjX1L1oEm5hZj+RfhDnWwVT
pWa3yCxd71h3w0f+5u3fW90JF8k3zVbt78/DhZWH1CT4BwSUqNkTujH2dzeLI5qS49JjzUxXIz47
MNr+gpSSB8AleHvjB5KcuTWGfRg4iQe12cuRR5q8WnEmSuHz7PUe8vWK+qTfl5r7+oDs+0Qmzh3I
Bg1uf+iEAq4SyppDRFzC5pZkvJ9JdpopbhF0X1q67674QKaSK2sqqOq7tkmfqCbEolI3F4GfUDJ5
DfrI/FLQK66VpPArFUSVqtVogPWaRxreybW07q/Mc1cagCAWUGGyEguc1LUyjm8VuwtPq88LQgyL
5D6N00knBXTnHZfO7VsZwvc+cHQ8RHqVIy/dyVVtKjyz6aknLDPaGW+iV1qI57uJNujP6omG4t1W
ZSbBqGjfwgL6thB8kNrx1Rp0SX7lpPk4QRhUx9F4imbfp980Afnyx78MvqWMZxaggMr+HNF7Y3AT
dWUfdaBnmnZrY9dY7xsiW5x14hhWxYmCFSnuzIja0j6T77nyoORlDVRnLfvScdAqbSKRF5PUFbMc
Yua6vi6jZded+t786WY8Heawm2NlASWxiMSx+obtmly5wKc6Yk8GEIdNBdh79Hmqqo/8VGHrnpM0
ZTDAoAg26Znwrq87bQIQd6soWy2kc9BqyUNDsOiRZjVwqjLJZazOIBpjDh6Ki8ltSzDF3o2GucjL
hB/DnPp1G0t19B4vUa1YctTU/TL4EpbVl1TIRo5Pd5cN0WK6C1QDnlnE8SOifiqmlVHwkae5ZbpP
txi0oyjwMI49lbBCu8bxgM2staFRoAgG+u+V+4ihcb3LPIPBYcPcktz3zi6wH4Qv9cCQpOI+W1f4
FGj+rgYBue6TCoVLNLIz8ANaW6gIq4Gm1yE0/6kPgKBcmj9M+XQGvcBFFLskk7VM+3d6XoHr83Kf
/QG/axwytSU4GpBHFVP1ls6szFd+SO0WGExuDrZ43LbnHjhzLbtZcHxUFjmnOibYCfDWVAK+jldr
/M9vU/13YzYFlYQhp8ytEmp+RX1fEWjh83XcZ4hocVfcAafLeUMxH3mlPLUe8wB/xVh8ooSocUCT
ojmCRU9hr5BVDYyJ2CYt1biiwDd+WM6Os1oaWKilsJkTR6U64YWumUqaCRtXd/TqN0DpzF6x7Bb1
U0asx+uO+4xwEJwILi6JH2KRizKxRAMs0yz1tNQijv/Y3PwHZMwYoMiTuH8Xfx9iQqsfoxVdjn9q
Mgoa2CWDW3pGdqY1AWy5xIKb+2iuYmvPRfmd/xchD6FSq0YyDGneiZoXMBiwoAaVFIo2VRxwv98D
lG6PryZPQNt6LF3NqwRVNU7OllLnwk/kHYjeQ9tTFDjmR4bPNcV7pHgHyKhLHl4VX5hB6i7iGLr9
4yzBhzSiXi7gTqAHmkmusQtDZ46xYgxLIIVbXcrB8eYsXtyPoXFg8h90Kl5je3KtyX6x4qyXyvbX
KfzovKwK9Y/cBGtCi8TNyHp/Za+Xc5y7Ew5OZX++VcqFVc+2UdMQvnWHSPJrhNSjhcJW/1shDDYZ
A/SFtigNOF3u9hEhdWN8WOZBdZ9vtbXDrGDeOtix3MSYbGTwZu4y+rYvBI/d1XSFSvaEpaebxFFF
LhhNY7nhJTMnqffZJ+pPe+24V/svklX+VzjtMWfGO8cU+Hy5lugkWpvcOseF7H0CleK0j+0dwKig
MCnIGGBzzv7fs+3p/pxqSSKB7VZ9xddF41e7cy7Vy5QLzvHXT8UCmH1zQFDMgfplICCFojh8GmEO
aeJPcujP8NLiXdk5aLpmNhY2jaTAU03lUzZnhpA+Qlx+oVKMlx+bfDQtKsnb2pYYyF2uW8cKoXv4
db0bK2427x84BBeTLn9HT7CYLrw0Y4TybVwLdokNOCtGo4VvcswXqePdEoHJrDWw4Hh51hIU47Dh
lLC5E5NGoz+2LaNot3yPJk2To+HCVc/w/+2B3aj562oPjwmp6eN3MzbTtHnUemEI1YRMZrD3+s/x
fGql7Gsh6Pkofx7vDrYGHFJv/dZZ8IWkeBGox0T9j7+O0cEgMQSmMFIPGklZIBs4dYOk7xpfoi/O
wJeRjGvQPyZj0h7wwN+JfEsaqzfBoNghGqXBsye6RF9ATRpDEHazq54fzGZjpbBcH3CJISaBMe/F
YQuvKf6l7gFmO/gIr/Tzj8uncER8cFuE2yp2O0mZModdh1DesnsZrcZVVECm+7G0/4eDUsElGp0q
9JqXAu7fVGIY3CNCjmwUntX+y/Sp0AzpGAXc29NmSiJ8uouD9xL4A2r4zYRIqbjxLYPqmZFkVXbm
vNrw2Y0VU91eXMlYtX+2aXhc8G0lU7hueyILPNtooDTkYylu2/PNoM1odL6hEH2md1HYXhT+5vHz
vc74nJoLK3BZatnSvgStXtnQN3uS4Dyc7pjIaalLi+7jLDA90P0Ht08I94IqGQVXUhI1I9HO5x2V
k9RU/RO/7UErZWaej2oEnZhzOjPb4Vx690cSSpdXTDFZzgmgl9dbDobvh1Tmn+IbBDR4yJ851/v7
NqZqDW67BY24f6PLDLhV6a+ogAbw+afnsSL5fQCeQM+9DT3ZAUquAHQ36qUuoSMp7aaExdeR9NRR
pdCY0jYawdK/Ilzt0SQpgtpG3gDkSzhv4K2RO7uFq2X+GjWAwZqJV7ktLv3pjh1A2FgDrqf1Le+z
7p8F60zliHm4BRHsbsSGAqWABHq1qCFF7Rvlx6WvMKi9aJ+WNblX+00XRGViA/TknxxKiF/SqW9p
srjUCVs/eL5niDaFnH0EUgcjVMqD9wtBiZkFkJQklyArR3IMBESXUbig+xxh5kVgrSbmHdU/5aD2
7t82EmWDX+wBhnkZPgoERMY/5AcoS8C4oUYEaHc2ruZ0kiMn5YUkejlpWxHZ2+Gsy4fa+GmoWJmr
rl1s+pFSE4yLDPNleUExMe5/NoHeAilp8hyPss64maFhDmaLGPduwBQU8+Z17D0xgKK53LYPlJ0X
m+RYBj/z+SUS68cXZB8GADY4SYatT3hBb5zrzGV7Mse2R0e+b8zEhMDLCRdCb5QHbMOSAcUqAtbc
kB4136grIXPEQ1i6hsPJjfJV9X0/JT3i0bVq8LU+W1nMwhlDCGJHPxyhDX2F91hOS8uJbGm+jBPC
1Erdm2VBdkRrdxjI3cfH3J7w82Gjaq9s1VGmXLoWWd4WuXeN2Il362+zzd1gfFq0k+05YPIbmpjL
ocurFw+8veRer4Gs3KqYEuVV3ZGLUK5RhgNE07pAy9GZhEKAK+DpAFBC18GOxyhKwEPzUX4JofsD
fKX4bROY0leJbUq8WdhCzFb+WVhuT/GMWgJU6qpLkTg3FI4Szq8XHeH+fYmJGknFTZC9oNWQYLRt
vj5fFjNMer9hfBmqlcg6GAZEnkGVOL0Kfs5Xz4vbgB5zl43tHj9G0p4jn1YEIlp8yTloUp2F62oO
doHGyv4Cfqd5hYQErcpevTpfRBjVCtIVDNEYlf/tfpZTXaK6hOqgRHP2qElekTX6fKSywDDXAqua
OIiUE+oek9fDzqx7lkGVE1VXwE/8SePCAYbfI09UqDuiLq/l0BmufuHOnXiHnZmbEuozv5sYz6TU
OGJR2EfsqcOY5RpHvKNcIhJDs09M/ATe1NwcY+YBOSyHUPWgIelnqKJnjkSBkwNr3ksk2M5r7SpY
rhe9vvolHqKcMAKZ8BdRi9BKNEMirb4jAnXk9Z/hNDkpHliJluAGzzDjeRB2fStIsakM3ybhNYrJ
/D5D5uR+R684Gagahsr5obc12FYyRu9ByLrNb2oPQOegnSvLKyJJKwP6cnBnrmGdpaBGkrEOq+bY
w5cQC4uY4Voavq5IIBforenqz62c/mHZcMWugiCk3OQAgtlfSj+KnPSaCgNCQFlYh51H7IzNLzMS
OVXWVoS0cTY0entJJINscpxIPNrShch6KKrcjAAUUFEnB1DnHY3ztv3C7cJd9sB8fG1B0Oepa++m
rFRJmhhBAZL1aAXPc08H13A7hE5ohykXZdZXRZd6tUVjiCRekZTlpSFU3xP4APOM4uuZeIh+fAnl
7LCnnPo4y52+2bsLcBnjChAr/v25yrMgKEmTJHd02F2C0XajnfIadZ+lb6lvRWQwQMJtfd0w4nRV
Ipg/9USAUqBUWcM/9D8XBXxqRgjIdLMwyjrtJ0j65z/MxYrfeBHEvmogVlgdbpaeYFMfzLg7uMB0
rni+6hR9fsugv0Dli0AML/1M4tv3OLR1XTwzD6UfCUCxnhCeqvm0aNgYVEaqcMk1IhkK5buCpHwQ
vNAufbfztBte2bitFb0TFFAAnah/Ey4/3leccU6UMFgYerRDfUBYQJ2jCgs4acC1l+d2Z3tuJx8j
TzS8gQIziDl0t4eby5TH3uui2wMxoNmrf5FpH4Hk0s+FBKzSpqTIvIVm28ZpoH+PbN7yDser/PDZ
sczcDvv+zSkFxaBGZsk/O+6sIYDMXEy3Z4VKxxVPEV0hRYw1R7Db/linAufl+4uDStRo5HxgRTWH
TwBveEubO0m/h02GipPjILtDyK2Xs+l/V29eB9Neg9RuJk3rRPpaREx6kph1JuosehO+WcHxDK4P
/VfZ2tWhCfEnpcTIprozAyXHabrN/aewz6r8nTwF9YYjqSlB269izuxWM48e4LDc7H0z2iK00/4n
Unlkshr5t6FGw2Sza2ZFtyfqALc4IbjnG9vqBp3lY9yyZ6FVnsHUfFWessTho0ANA26Rg2ar07ep
9cJkiyTnNPZvTEz4n2WDHAQHHAqHixAmK8lbTyMPgXQsMtkFoFYbpRVmV7WkryYAxI7WJAnLOUOy
AHRq23uT+9QHwUl01lAxO/7w9VgCLDNzTAoyI20iOebAV9LXJ45MvAfOJHQsYBg1F8sy4pQe2yjc
+kMCBwNBl+xNsE0U24HXL+OJqqkGxlIOOZXmSvX083jc6DEI5Xmiku7NTT1psZMDkLjfFJba59xD
zUdEct74onGZjszQGMjeK0QT7ZkoA6oRzlAufZRR6wbIpQx3Bn4ti48wOQUg1tOMK1njSSUHWzyZ
CiqtzbDj8kKnZn/+CIRfvo98Rp8KaCfWzho5MqmeWUJUBZ3FLd6NcMxYREoam3VjkmAcnHJedO0+
uGBPVyF2EcgHPt6Q8YEix8ipFs2A45tE+k38SAoe8iiNsXGGdYltwD1FFKxRtdJZTlWcalH5lUit
jO5HY4cqzpQWoXZpwxa3KS+nEakQbGfPeRG8dGHahT2C4m7yZ2qvKk1twiWi2zR1jM/3ENXpl3V4
BVjIVu/SkD1TOr1NrkszfHI+eL7oNOo+wuPCPh1HAkwyr3FF5CEixZCheUsiwamDk9eAo4MaVbNW
uumnEM/x0T1puHwDOMCjSxIbNmRvbnpizxbqbtMNFhP37/j/SYotNahrS6yhMytwmCvGH+U4GxnY
tWAtbKUlcmvGDGHAMqgHHp65Bkz54E+S4ktbezS9qJo0y5mvd2dZCjr8EofJgYoiioR8sUi3YfCD
FqsCfo0eSb+t+7cVJmI4eZLKm6mubZtN/m03CPrUH1VqkbOC6so1p0BIM8v1wA2acarwM4yDcERF
kHGQIpVhTv5g5OrSHBVyaPs4EvKG+2G1f7EFsLchLbMZ/WCiORbezXUy3meShxmEW9EvSW8r2ntT
KHAQ++LOMLH6piaAb3XKRsLRXnC8Tolcn9zp5xQ1PHBS1UKkdedKJyJOAfem1Tpk8ch+Jn/mH4wO
1g9kqzIbr52ibErr5bnZk2d/EPJX6yHIXHcoZpP/BS3GZQBwhfb+hyVRsCjSCImy/SHNckLRJBAj
MO1CQJCOo/ALa0ml7z3hl7g+4FxkPqdilveGpSFu43kTW18/xCG6rOUo2RCwcEIDQJzShi24pl7w
XEQnBeAYTgmlZhy91kzqfpTRUklkzO4pjD8CYtmAebPBBgWohD7aUgMwWtchwwJP35usCwsxpGT2
iFhYpTEk28NiERLu4296lUlk8/a2qmwL66QB8wNeYjXz4rQQg111CeJ7fNJN0gPVLjiMZJDo8PJg
Ihh3HD8a2hh5IaD8gqPrwf7uf2Fk+h55mHiCIXeBsAXkCrIalQQ7FcbxaBRcp6TS18UpXJ8jnfTp
8P8QHgApxuPFcMXFet4KWNDdVYs8Rh2zM02NrbCO3IJwsNJpsa/NIBUjXoAhvZu5deAuUSOD87YL
Tx9qBQnsUFRC65FHphzwictlonYlgUBKpFRpvXmguBMaRzdpfajitcYJgiYkqXavkXeukpkcrQuq
f49YdXVVluYS+SIa51yxkilEb2iw5Jztf54V9PCICysEwM+G8TgfnwVjxumst4eF0enYLXb7Q+Im
9aBA5XaMMt9jzyna6O17tc6jNhpMG0Ur/7rjY8fD4YOCbdoXoxuxyKHhX4SPmiVlPzqfoN+LtJeL
PJ1wWGj5vGOpO17MDgaEbLOA/r7BK89bktyncPdulWupMbdWmNHC9ic8LqXs0UIEF80VUOYXA9Vo
JuqXIm3NmjyqxZ/OlVEEdbQEA+JBLZXRcUcr1p/0+YA7ViuqXfLoZCoCaxoZDDfsfTvJ05dKMJLf
U+4t6ZjD350rsA8ZabCoxF+XqKZxMWr4GjzVHq3Se4ElcKagyJu0C31qXGDRF2DfC8mK9XAy8dru
Y6lZ8f9+9pBPb6mG0/qA2G1KNpGeQ39kj4MnFrFDkTy+K0+FAAtmuKaRyAJ8h0Sx1X2aHWz3HrLj
kgBzPEo6b2SMTU6WTN5M+0SvjbklNLTO2TgPH9ggedXxZpachRtoKxrfwY9VHXzd3gtDvFyjRNuz
wCu3/39sYn1s3vycb0aDo8FBP5/Cwj35SAg27zTy1kF1Ulq1IA/t3Z8nq7PpMSFJbnMOi3oM8ddd
74wOQ0WW2bFP1R2gH1zG7AHzwlV2hOwG0zMNcbuOSm7IvW+JjIOnX4KvXL2FL2lXCJw0fkLO8BzK
/Pmb5+FRgOPrZlKzIi6/ll8xrMNZl2/kpuRc3CnlYYvw08FTjb/dbF4wXscou8//bWUC6YcjlC9B
FtiwgvccZUpWIz9P/wx6ODY0YW+bA6qEG/Z8/VPLWGujpZaipW3rtO3tmqKq58Ql2JZx+NA2DCAp
Y+LtaPGMuM1hfLDo/0PgVegfw9Qw5OoPF0bq06DVt1YxfKWuOtunGeNg7gPC3cNeKloD7BiAm6Iy
RWNaTNEvcRUgdHhXMvitdiXN2s9GzGqjH14YyGWBZpWkrCE5m0hJDq4F3hcjHCzlgQqU2W51atyv
OIAm6NWHA9XUxnx0E0AFvyUppozJNJtrkXyiAHhzimkvZDonOMajcS661XqHsBbunnv23Oo/cGBp
A8t0ms2/bLDVmrPd4Uu7zQPSKw8d+uHbe9hFsVT7vu75VmV4mG83waP0RPNQvjuo4XojXt563pFN
+83hFtpcM7aeFJfbn/vlcxK7RFFIptLS4pJqWz7LSu9jR+HahhVcDZoDI3uGkDoGsKDElK9qezBs
d4b4poInP+nAaflqHFf3o8iQvVBOFOIBncoxjx03tfG95qMMd3+k/s6ZsfNuW4PCW2O54WhB4P1+
Weh0mgXnNryQW9cP5eh3zvg3DU+8co2k4RnXfehF9/M5yvIuSFvXcXT6Cy6Tpanx22idbW/RXFZo
E3xw/iLo4IHOPswjzFz9ZuI+LSlbmUjzdwwUKtaBqaK5EBcrJwtjn/bH+pX23VYqUS7PgQb5IBub
mimOj6x5N2ht7O6EsHsgJ8MTwLjKFpoZe1nsBwQnS803SyXsKygwOVzl0XLHT8SzasCI12+HClLB
iGYp7pOpzCZOm5t2vycvocnqN+lU7uTwf/3n94R4WznUNr9lyLWcstZYgPkpa5nnb9ECQ/hs72H6
NtUoa1+aupNKVy7E5Hjfiko6YIiI3e+x3JoItMrFkQHHVq7XMMWpHEGTs7voDtl8f7qNZ9qO/iSh
DYpTcAiFSTIgZ8xxgKNp9GdEdjN9LqPN8c/tv/o3I3lXFnFhwQLoeX8HzLNg/49QvcBRJh682TWU
Hw1i/0UGL/YBd5lLjy15LrN3XKq65PHkwYcpEkvPHxyzGKmfz7WM+ERz6o4V0ExY9o87QKnt8rVJ
nmdCHZSkxYf5/MXFzZumh1b3pgHVbgb6NUmZT6TctG/B9TEL4gD1s1GuoQFejdxjaqlARfcinQGA
xiOSsHayXVJx5PEdIZDcGK4L4zaPs0jjfzhgJk1Tn22b6jCqUPHgTtUBPbO8kx1uo5Mq6eUIN93/
MNwIyuNyU+n4JggyewNBGlsbd+yDucF1hYMMk9yQNAL8ZVHZvX10rZcCx9WBvS2zgntEWMBC3dqo
9gf10vgT830Bs6n4QeFwjzeVpCJ5hoSeEXspIz00kesRSfLHsPxSQ2fUcsQO6CjtQgxC+DVX8ITc
4tE1Rlx7sStkTAD+h0RS6WFNOudtR9ovBk540VaIFqGF9opPU9xFhTxIL8etN0r7mAI/2gA7wEUM
5c+LMIbnC6B1ICeIUVZLJpSlZaNwKmCV7wgWXvCSSX+e8zY8myC0ogV+qZJvtDlp0qsn6JwvQ063
O7h8119qY8qxWsvaHp3F1eFzSD214UvK8kA9kjS1O/y7dDTyhjmw2js+zOpFveFNjxw4ifJYP3/a
Sb4cdWJxsis65eB7q+4efZ+dD8MNqvdsZrU1lXV/zmTCkPpHSPa9hTdrsB6wO7tx6huJ1sQDyBaJ
2lUW11cH7GBsGhy9aHPNPke69IQoalTIqZTV/O4G1PIht9meVi65VEhAIFIjo50Sr8tM5iqWS54m
lM4rpqztsCV6fN3GMZf8RseeNublqa5T/vOmLziRg1K2XKH9sZvCbAFVYDachld6vVNT3YoDTV18
1i3J1h9u6RWGZLa0iotENWoDbwvxCMZm31go99c0YLwmNcuIfGWp0vaO6JoprPlKuTR51jbePQur
5tFWuPy7ielBLa5G9CttKLJiPTyFtwV0jB8QWNd2Ad+5m/j92Y87VZY54YHQ/2NcmXbudesSqSMY
bnLW4OjkhcA7KfrmmoeZIjD6EjYvtqzUaQDBWbng2eelUubKYUiUjxIz1ZqIX/jO0uaJX2iHawEn
5uD8iDR1Ld7qgMyZz6ilxcGe7pY2I5azOXaY5kxFAQ8aCd5OyTkjaDxXE+sX+D1DTJ6NqATigIYG
pKBUQGYUwY0Dc4OZHQk936K2oZ2npHihBzacnfQ+Gt9fvQqtQg1TCOPlfpLkhCGF0gXWTm8Rr5ML
GjKHZ3kBU3+yBPTbFoZhWckwxqx9IMa9NZalQHvjXstxuXTjsWBJMGaVdl0+UkjbWR2P/iwwKCCV
U/rPUKJlpxPqlcqtoV1H5V54PTGEAIRemkui1/ymanHDzihKlg6bLl5/MTctxnBLz8spcQhkM7WM
n2K75gaAya6ky/RUH9TZqJUvxhEg/xyCM7+jbE4LNpPyt4zlo/sBuPq991ZVwfI5boHjZOtFuG+k
SgUvxulc+76tBYkQTsiXI9UR50A6KSoBTEk0q3GJEvP+GnBWRixaCdaUh4Ur9uWcy6uw4jDIAMeH
hVJjEthmduYeTW3EAzFfMMU2E3vvv2K8p8IcQExno5rN31zzsgXoeyrCXoy5O13y0JGiNr27PvI5
35t3K95DHz3LRJsUkH3A8jAWQ/qeUTYUWuNAyCN+M/tuZqb+BYFxip0w8Pt5uN+0p3gpm8poo1nt
yWSRkxJ551/Dml5aXVZlh/Heqva5qzd5E/mV7K5aGwolqm1R1f1dahki/rTrYw8ao3BSu8xQBQGE
CHALuA0TadimvyCzpNmLvy8kImOaPhA5ZkUOLZZ5r0qD/okP7Tv3jq70PYVZ/xB9NOxyWq/vAP1G
6hQLafufE98xMq2iVf0I2cjW0JBWaYjcIMEK/Qbi05m5AQdfNIoFKJKDK9vfmFC3tdAovuf2Ou6c
PPEVXUUQmhJox5SquvT9vFMpmfWjra990nanyUqNKjPq9jvaR0i1CJ9S3s//SN0Po71M1HsMRFJc
3hQCuAAzGqBYdvn2JJ/AtjjW4G92U1aL7kQypffbOOzjm0m05gKOLnhsVDqxUUcIXd48B4zzFV8K
jsrCgB9lbulHfD6Jm4tQkZ65OdxUSCQbhoG2v7oeM3/dD7qJfQI+At8DF216refJcV9gDG/WHsgt
hxQnP+WxAZqxwFjs1xHAL9Nv9jTAn/ClpqfCI5/6zBbf5SqH5wV9ZN0X3jsU/WgdHpdgouZ6uif6
fQJaTNgpHeJaybv6NQulvYu8V1Ii7Ysj+/pIVjxEUU2nq0vCHYFY5ypeUkJVOTFvEwql2mBrNI4n
FOG5Jln2hR5b6Zg1ESZUXCZXlhC0kMrAqjSt57a8OZ6Bk8NPRJ4bbvnbDhvU2UX1Dcmpp5IFKKSM
UF9U9XYxMjSI/5ULH+AUQy1/nEqnHfpGV+NaHYsRNyETgh5kLeiAxehUkSEaiaLFWQZAJmnwyUu3
zxblZHr2DSWpEKKjp1ZYOsd/W3fcfZmdg1T6R6+FdZowFthcZEoBFBdI4H4fMayysSqPt1OqIB4T
nidyQniuiAROWbEM0ydbFhZLa24GW7JHUPRjxAJeliM/ibAwRL/qipx0x8NcfCJSCXtnqNOQNYHD
JQPIBnUnmLLd5gW/+egmaxlLq6OOoHh9VVrMdNgNFy/Uv1n4RHkVkcznERyYQWvhzUOPDoPGEVnn
E58MMiiE+M1MvmI4Eo2gbr/jzr7Rvu+nnNJeoPEl+bapjxIm6HPp0HA/7ZqgunZ3rLiePQYVhdvf
sZYxD8VgKDBD3l/3GWez6o6yhR7fi8fS/5xOxEiRtlrKCMqMD+C+tQE2XOwSfLGXY2eZeF+iURBY
osNp+6hFYrPOMTexT7g5ijkxzCB+MZQy7zIvVkll7xzJ/t7BkBSGj8Hh625QuXuXlSGU0StdwGq3
4lDMqFFScoeNkQB70xwCKZgmm/X+ThMt5X6VmyCqmFkwVTFEdz1TPectizQHcmlcU8gDsAL5r12G
YI7G76viX2uDUMz1j4TP4DjT6tiYKzFSmMwJak+aHEI1p87GeeXhZQ43nW6Xe3VExwX+K/lOk0Uu
JYH+nCCM7VIyfk2qzHHpSjcP8gVO30wJ5yCe57mSfO1sqsAYAu51vObAjN/op8VT1rOPJb/skYky
XqJNFHq9aRoMfSocIAdPjCCXY5JJgCCGDvVohgeokolwRIj09UN+pH5xXAXe2Cm2betML3/IweP7
MlBwOC9GYmyWsNFWwv3kbbaYC/VkJuLhfeUgHST/Ax3NjgUlDgFtWZnSbhoFZjgXuiCrmrPsZ+W+
dAgYOh8LAY8+SLFRx/j1RTanU5YGS/21QrqlpXr2KUP/xwnPthTmAxZ/tYbYDo84Qy6Oi+x5CVmO
2ylPTwDbCx5E7VRM/+6c8LuVBlLeNh+iG6O1WuHHUVVFRtUQd/zSxs+aX3vPyyd4Ybicvy0JuIUv
jAjkMVIzj/r25R6+VaI+9/K6yc/Qvwuc2QVYDIdKy5K7RbCyKZ00tpxbxVPn+mEl5rUmzM3aBqHc
P8KOBCS3dhekWdX+2oq3TvJUxot5pl5XZXdweBELfLT8IG4DqxXYOXkDvLNkET/aHqVkk09+1/wN
Vz4rMCg48/SAZtnw4h9HDBVi3Dcj5GdYUGFVopC4EkNZQcu5nnYJOuYTZp8/R5fKTxDcDPCeHrLA
wLoxDFsEDvTnV1gw4VUUv5GaY0r0SAgJ0mGQWTZWkv/rGhEx+jJGQev3qHBw/YapJzkKRNRU2fL2
KFGO8ouuYSzhaBoS7kB5m405bWwhT1ckXShmXuO0Id5M+0zu28jS/gIi1YnsSF1/k9KSwD4cZYjK
A/+2NqaiD5zibiIhRDyPGQ002xEWFj33FML0p7TMUEXIjvmoVsuO5kotNvAO/qOFn8poKAaMUmUd
88opK6PdDw1SzeSiffQxpMSsAaF0ThnNWcBKBAOukxBpo3pCucdVAXqiDROComoseRd532Gfgg1H
uO0cDdyBwVQE7Pk2fpgZmS0DUi7QBQoXyxo3U6KtCkOkSmdnCpElLPq2vzK2w6XWv2P5kOgWj1Es
BHZCaD9wj33pysVJhvh1da0et52AuT8m80Hz1aHvfn8sFMcOeQTVvZ2RKdxCYUViT1HI0tTPh/VX
YpP+dldCa7G2lpkxEuWbj8/CKzAkyj1xORpN4w2tNf3etnU5A2s21Cqu5WTlWPqrv4vh4rO4EQ33
91twaVqKdO8DWge3Le4vuPBDwFo5PxhnG2ocSJZf5NWD45nEbCXFkfJFXOQjjN0DCQdpQ4KgCaMp
UlmmSd+6zskbXp6D3TGOGKLwgpkArVp1LpP7+6CDl2eZx2JtnNfpjMW4qmA+cFcKPkMCpWY51LUh
59w4f0+30UlNgXggGNU1dlbkpU+guesqPRyRBzgD5Nh+QYkF7OA9pbzGluNROe9WX49FJG4Li1fJ
L/71hEV5ldvmS8yFSszOvBew34WhT4etayW0WUaGgDqWHQ3tMeYdYkQLYylnM4BS6D+CO1OtB0yN
TU6P88UlYnuOxyyISo2EI8BLz8WywtPSD2WVtqfZhgeaNozaVBnF3Ucx9w08nEeUcvXRd47Hkv7S
hnnqt/clSLyZOYZ5oC901Q1MqogOuWd2r6tz6A2fUSC/NfscYkqV0S+Bbwdd7GlcsP6tXjue3SkO
jsGtiYdrBw+MWfVZ8ZDIwmeX7EKeJtbswaUNe8TZ1pHyQwVtZDz0DbPyOqbgv0kPNx/76XBXmO7m
IrtA0hU8XChs2EAEmIWXwtAQTcJOzv6IGlpPDr3C5M7hban19v2eU2+X5XLEHhhnOwONaYY+MJ4y
69rgPIkU9pKHQn0M8mq5di24eCpSByrGbp9HH31rx6iKehjMN8DDboHeb7gpcsQojtbtUlvibyKx
fvSoTZvPXxi1WEtvxKTTcA9pUM6MFPgCd2U961bBjz9ccQhRkTb61Qnyl9ppWJz9IHBGP9XwHKk7
NEDoGB4VqHOv/3Tsg1O4BfqAKt3UeHE4aIMcW8a0aTpVKSdBBfVuar6M7gNImqId9ql2Kry2tC4B
sQC4RhIT5baas/Q/3E95TNCRu78yIT40i/Us87RptV7FdFBGlYg5koXFFPPYLduePIgCmkRFNhOC
Z7359dM904hBJ00nth9yP/yUOAArrkIWc3fT/qIiynFTQuNPUMG9eDqoz5tTMuDBH6MaKPHGG0yy
7jsvdpGG/ep3CctCrvDYrwiTPNW1mvczKgb4zQRImQ9veGL4tMcb7p5866AXOBs+9CVaRUmkoWWD
OGFQgtd/MkHxmKIgcaMPs4NrL4c2u5UK5cuylsVzOcXMDZNgDJVmqhIs6O1efkxy1YJQt3u5tfsi
I0UHLa881XPAwiiKZSIAKhFI7O+9Ce1BoyJq1CR83nkN42B3/Mwfp0BhNBCwpm5WOtYDoRT7bCGm
GFCK+2g6Wv8BPS778BwBq36N3w4ztWmNkPKkSUSi5HX/2yZxkgx8NHh83wZsLk4eeO3TS4V7or7q
Zb/F543Hp/BmN0ymxakYekRQ4SYq00wKdgRw5Lt43gNAB1BwEQcbxkj8xlOiI2zxWJqC7XZKMX8m
Gy6Sh/+6hP/uKnmVGpiqW5BO6p8hgAixX1H8Xp78K992XwoMDTvLJFao5TzwI0F/jBWyuxxxowlR
oPXdTxumGXe2JRVng/HWx0hyUaWHLaxZYJ/vJ3s/DdmhqlAxG0vPwELEJDG/ZqQc+9nobPVEUJhe
K/4afk/Vb5qGlKLavJd0ySDypDx7Lmzh7gR50YhM5Z6GWpbP3ZOl8a8+hp/nZBTjBVkrIhESoam6
pA+DrNxRQEBFdMmgi6Uztv1Y07++KRVQG2bXaywVgdK2bbSMFDg7F/x74mRxmTmCePpT3D5KX17+
onCbjPXTP7jZGTNppRIyZd5sVmSbhpNVKKRtfgAhmmZYEHL67vzNoYYdI8Pzo+So2Qh2tWucdOb/
9/G95YAZ2btgb1A5Nrq12LDHKLg+YwycwHQDaT3oycmHOCSSXw/p9z1XgMdyqUKhA82voFHqNmhU
9tcifcvWjRNcVrnAbIrLgHPQKIjhiCXUa3CDL/solmCqUvGsnA6KxJXD3zTHr3j9Zqig+Gu0n4Fn
Rko6bYZ+tE2YJaBHi98BqpdaNOWx4MNzwNEnSfMW+LRzTmGGV7KLBtw3q1+IH6vcikaB4h990Oib
erhRirX3aRv8NKbTEYEevf5hLL2nRq8lLdT8OuH9HU6HFCru1dLDdYIYJBdtakkZ/EVRVLi3E+oV
u+OtVBx8jSvdRevge9mZZx2cA9gS0Y/kur3cYSNiJdHKpKR8/cCsCp2TfDDCjm4iMcS6g7f/iLaE
5mUz/v8OM7o/yAFyu/cXpV/avVbXrT5ZeziRDW/4I4nrSllLTCSreTdQ5EV02MA3IzcOgHV4aoAh
X+ExqC4bF2dd+/FB9gTkG9INQIT03MOsvLv2Nja8lIQG9axAt/50Xd4jAfrwQP8cMqwc0g6nsXX9
pmP2ecakwlg6RYQh5zeCG2iwfoHOAIOaYq1Q9JTFrbh8V+X6Z2tG3tn23PLrsmj00RZg5NGvtDQ1
lfBSiyQIcYadfpmN9Tn9IPS+HPGi0HeQyVymqdwm0ARdIDcvTicucH8U4XZLB26xmVXPEb1f6gTt
w+EgquBHs74aBdTrP3VmdSp9VBFVqn/gAlq1VZGwR8WjVBscfjwqdr1h+TVi6FzYLXtocsNZ2dIP
y78629SZME0HmfmJK/BrUvExjPH0dHr3x3L7wzmTO603g0wIYbK5H7gaQZK2EQxa4kvCgck7qi3e
/shmpdh6/d39+9w2YaPkHKKGgV6IFVYJfK2RcAaYcAYBNRGld+U4ymQNJixGXUW+ZabnPIISiZ5d
IB66K2yz0aheafKJ72qRV4T2WbMbiZEVcLbosFNoiUs9WvZDgiWamDUoxadARWJqIBfHHbBzJMbg
WFJcp790wdzLXLX4m7evPS8lUBwWqSxbZI4SpiV2+LxiTnRRCMEn8xBquf+l1U/+vC/pVo3Ao7Tk
hxlZkIF7Agr5B8da8/tobor2Ykb8yJbMJ1I2bWdnmnXPu7jcM1K9pQXZJOVuQMjCEGCl2mY0Ig+C
jrTy5YJHwx6DPmYuDQolusNIwnJHpAQ1ssyzJ1WpQhkuq+J/T1ff+xM61gAOKPwm0/7L/l75BzVb
oRoBzcReE397oEQyBoRkNEJ53tVmXU26Z8RCPSRTcjMvQ5FRTHIwI3ReQXPn9B2SShzgJ23WHQIp
fOTAbyYDkh+CJbwVB+k9CxyLUQvWfi9k1RBDu/pUsRC7EdS9KzZ/Rn6jOVkL75LXx4nnHLo+hP8A
3cvQ0h1rZLohDg8iDMV7URE2B05HBBZJoYqmHaPfi/VwTHdXZatvjIZDeKlEcJHjig2UFBL7k1jv
MC9S39zQsy9EL6rC1Jxi9/fOp5Aj6ISFLly0EHpMan7+wb2HEWH2iW7hia0qGhqaKCxTzpqSPXX7
pRIH2vZMdJuhw/o2dO+iJ6vPWfnvbCkoTiwDLwXbhqF63dnJ3Oyf5Ey2b+WiXZ3J0HzqDkT3Ir3i
+qfBqLa+KkgNqDV+NHv0eMXJ5aQXtP4PHK79DZeAqtKKkpCyVM0eJtHbhqEcYae7g/WHGexIx9E6
xvyUP4UaRKOzYOyGGYLyHlBgq2SPnZn5WNTiTV64FD3WBUjuYR3Bb5spMg/nfUdrtunTlq42TLMX
mmsjKU3MAEw3wRRaf1pyMG8m4KrZE8dVEIkFgzB6KDal9gaBmA8mn/DoJpIx18KUxs4pIWDb4Qca
wnVL6k2sxodjjUtn7o9iUUo21XkFLN/qhqae/IlQo3Xy8XmTG+ERhL2d6rA8KHGfpgY7DfRD3HwM
IxmR+G/1ROXmvsB+sZQLWaDSgoIhwQXSwFOGr9R0HsNhVJv3xO1wLSajftfUXc0YveSo+DUW/7rc
riexmRE4OymDfGHd/pvUm7J4O/+7Mfd3uR6psvyGNK2LRZ6VjGwpImcpU5I8vA+xN3WVvnbrngRs
SJ25U09kf0sQ/fJ0STlC3yQdqHiK3quda9je3CAc8hJPIBBrNmH/W3ufALcLoTt59ozROq+LxEGG
F1kTZSmkvGIAfZ+ZBorpTPCthnbH/l4GAQ+bqjn+mPRNpoIP88Dsek3MkL22OOcmUJZ3PNu81wVy
kcHtB7KNFMghXh2dnMh5g2/TLjT8IwKStlRjHH+npQKtCyXpTs3WNqLgNUXSLckSYuDN+Dj8T1TN
fCk3fY1v91j9JAG3WXc8bu4rXmAX4bQ7/AvXFkUdUJ2NokMe3PfP17lIxSH7dSHWVw3Z4U4CTcyV
MYhhCf6LavUCorkzSoFcSCOqIpuuzREGBZ+fCZnot7VIxaCwlQMQvsXHatLQxoU4QINU+z1vEc1A
dapWqeDfNlTpd2U1lqDrGEsDDRPG2xLI2sfzlXRDPQp1cJ7Uonjf0SU8FMR6SBIvKr+b7KTXkIzc
Qi9Qa65h7kQe1kvpr3USX8Hp/Pfe8w062833ZTNvQBn2Jhcr13lY/pfEDYu7FI8VnBBqwOxuBvjD
0hJJhfGcVp/ZXKFOP1ToUtRh9cW3C4F46Vjdht5vP099NcwTZdiX4Eb8kYLvWuauc6Bg9pE0bjKE
+Nhm2vIiZbwXNDdgp8x+hEfdDR16PPxzTRP9nJOanMVgBRCMo2u6uMfoMsbzh/QOyqeNlpsX2Giw
e0bPxZ5yFDDKm7k5tB1MPMMzhzHIcA/e+eW+jNBa0NgLXip27aR8MeHfoiw0PeOqoPoy1swR15V7
ZatRBPZk8m4zvbRcDLrc/MWd51wgb0OmI1bo8sxZ3zk+ecNYecqRZ2qRzoLUgOAxim2L6jLm2jMj
SK3+lNi7YDUe8Q5+4Wi4iLk/zKCznWwIk6Yb8tdIeFqnOtnJ+sxqFP+JVrFLNQcwi/f7I6Gcxh0d
twpnAoxLNTfYF1aoJwInNCtXlM4gYLMpF+u5uC/2WhJQ3pydE5RnPWgjTWWc9397IYUe5TtpDyv0
9TJ7xKoKkmng8KTTcsd4MfYXE2R0MFmkUP9RI3ZSY3/hh0qTPWyHUPSIxkD91of/ku/bhQ1ZnHPh
OKNAtb2deXk/cxoxVRPhtl7no+iSCECWkzVgAx81sUU8brx7AeSk52ItwUQcRpyIZjol0MACiT2H
h/MirO1TStCjUpLKjw8RiMF+kpTbRN4Xy3xmDIY4NW/A46KYZCqlIOiRWUBC8MB+55ndoVrf+oJp
cBnEWjjwsGPZblRv+6OvfUSjFgY7PTirpRg9MNo8M+aQGMpn1ohzf8DCEIZgATWNpvwu87jWvXpW
ZqMtx+UridTk563/mNUX9hffKfqIqgzjPCEhPpoDWlL+Mi7i/uM0attGpM88A3WLzNUiI+DAOtny
hpk6/3V5tNfRWYV/9x+/sOOEG1xg0QghTwTFXM8osVxcESH7bnHDIRuHjLiU70J8tz6TTxHp8lNv
p/E9qa9pp2eosvYxeywirhvRo/PsYSKcos58QQcdB8d57PKPzSTwxXxyokgcaGddgJGzICLz96Iy
09USFF7xq27nUf9NeYbsceVbiM2mDy8Km672LcX0s9Sdi4zkLbUCubGXEnz/2yDGdNSq2jo427YP
hCFB1OemIrzs/1MVxY5aYcc6RFnR9Cgjwd124JxJxaIHrkEYCqLNw+lh8NXULK1PZ4SA+cB9Exz0
YYYA1+4kDStCfHUxVjdlo4L8744CidSmasm6TuFeXvRyXOyLOpD+Heec/HQtI0/8xxt24PvvAGmT
qwvC6LnjRJnVqg4NbZLElUTZsLSbfMZMIu8RISj2W5eL0qMAdYYTdqFMTGi1/4Cz2/WPMeM8hFnF
Q8SPK07wULsuB/Ci/L6yvpt5Q73qR2B1HxW+7Veuk+WDs6C8+spM3viWCRA+S4vkYXMG94NANWdW
pi9Ca03I30ZQN3fpXlOOzE7RK+c1LavHce9chI9Jqjz2FAmz2TnMZSTrvQRZxVkHPppUf80MirYP
GiMUO4NAgfy6QcEENHRTO8UBNldpQUT2yc5Whsb9WI00nK2R/69YVnGcHIHAaaCi3l6ARW5nZSJ7
TUV/0IHJwl17Jw06dspgBQGl9XfRQRaIfq1AGW8apBZupS6hPwkwFF8jUjUCUgL0Dlqy7CAxRRvz
3QGAoCF+yyVBFXlKjDGFjgi+RKI8MgL1MkhmuL4knhdVkAvBqLT25yNferFFlZheinoYmheMkoYH
ca1bWh/ozV/A50/i4TtvV+bo/5bG2CTxp8axgEda1Cqr9+EGl5XRjk1L0gRofz9XNZ3gedwJLlsh
ZnDxQ2qYwGmIBU0qTDNcE5RA4ECEk8WNok94Cr+sG79GJHdC8P0ZBqhE0yqy89JrBvgoNFOC4qpX
pni4urbjpADDrHRdrFh+VxcO4kk+fIj1jCVk46Bx/J+yJki6paOSAm20LoDvU0NDSzOfZXaPNCvD
i9WML9yeKPsw8181KqNQlxPZB5LQL5Ut9P76qaeAd7Z86esmke/I7PYoo9mfptByVJdgybHVmHvH
yn1rWApYcOEWltC1ef/e0HBvSDxRavw2xcMnHgF+FVaDl9vd3H7UzlIKUvhQTamv3+3jFbXrfk0S
n60fYrWAG+GNtOw2Z1eu438oM13I373niQKRl+JUojwqqGjoOexpLDK7twb2NqanyhYLIO+BwjXu
viEQKKjN4vVh9fgjNK/H1aHfm6MeVRKYTZV5L8DD2T+pic7m5T83eTQuhdKlD5OoIlFloHdigSSB
iwvkgZY3Mj6QmqvI43yokco4PhFn5dUI9iMJ5661ChSm3mlSgL7RSBBR48ZTDQcYXeijwS0DeqhE
rIFUlNGu6AdflNJezfNPW9JTn1SjVwU+zxhHA9GfHIUP3h4znlof5ih7iyP4f1s/Ra7IAXWrbFzR
jkSR1SKJG7rOQxO/sw5JIjtaoA57gdEogr0EhE6KZ0Y9UCyVJFOV95eWs+PamHvWRbQ9QISoFHwj
i4WxyvL7HgCu2in5hqnuy6YmdbZY+ucfknIllnUQk0ZMVdHYw4qu6c4ISjdHr42Z2gQawv8ltZgf
1idLTAboVZe79b9yGIZjdDfHDCeFHMBlDtpqtsYQKZilTW8k4p6mPq3bus8ANiGYX13fO+K3iAbj
y/uVXRyN9/gAs67PfGa4griXxCMWWxFlpM2czT13eent8wRLTi6DfXxdVbacTC5lcfzaUP16Arjb
KjAfVxZcidPAbRRTB9v8eKfrs831c45m7zozwissxSogdeDgGyV+NrNvM3xVkLolG+d9Q834esCZ
jSNO9xwWEPGXHipoZ+lYAnZfCGb+16rCI8wtTATkp9hzAAYtXZ/XayqNHc9CiCaO49y0WB6v4tRd
Rx6el5AWYZs3hvKTYNHdAtywwRl9bxUUKZzrYaLHJRWf85KTuYnOa1/u/0pI3annE7VQV/WMSt2u
0izA43THINPUsV5g3U4j39cjrZO6FKpAFO1hHzMav0EJrZzCGUAg/4EGBzGuYkRD63yw3dDQCDN+
lR+oeBuQC/hXIllYdKlqxcIEaM1iuDpxfhory/2BGFq5uH2GGKSlLa9ePAN2aWpiJwzg2hSeIwHl
GELcjPsmVWB2O254R3nRFavFpH6mhxUofbD/FXbXyyZ8NXliphaE2gKNAgIPqBC0bAF9o8AxdiJ6
pmHShaSxz5PYELKcO69DJpDNeRspsK8DPnFminRoPmBwRe2VscGd/6jAW+P7dEvgkbRaClXXfxPc
hVX/GW8ifpLEUszvLKFPo15rkwRUlRCybyP6Ha0ek3J3g1GfjOn68i3bzyyYa2q8MLiyPLacAmGy
X5cVgLJHQWhC6sIFbVj0kHGm3Jd3z2UXMSc5PrQp75HXG0sJrzZ2Ayfh5NbO609xn8YTZm4OqcO6
ACwqYX2nLTph/cQ5hVhaE4gR3JlRJLPUTSR1xudQ5tEdi47HmIBet6a4eXDM96v3F4Q/hq4+nUcw
hsCaEIdMxpMrwDrZTi+wiu/TuYY6ULBbaT3jSCXlSdEMS7mWNkIh8lUuuvsya0dHMZER97BYouCZ
PQ/CCb887T5suKzuIifwH2jAHJmOEsoM5WoVuz8BtekNsdpERGAlHuErId9msIO46uG1r5tBAkWY
/cv3WajYy4EALp3xGzjMwxL78gJCD364tqAewoAPkMWlUg/+XGkw04tXoSRze2/i9VJWXH4Yyfbr
kBMUgMVkgV2XU5ksIRGiT2xRLy+g84x8CH7Z8qXfbNwuBMUwywQLSn+piHlIXCB6K4bX1AXRrVDm
zUPlgiVhHGoPxQHs7x+na0Gg4FhYkuvFhxeeocpv0XDX3z5VW+9LXnYMfZL6RW/Lewkb3IsyGzDs
z+qVt0xsjzxRN/whZggFmHA3TkrtxTi7P65oPbynW/9Ca7rsaxxJoJzh60dGi+AEA6HH/lexdQwk
BEBv+Lf5mVMY2mX0lCMw/+ftnkkIUsIPl9Cqk1IT5SuQRRd9X951oBG/F4miroH9JA8Wma4PfwhI
2hDoufYZggCwZgpYdBodu+RV9ai/m3mjXSIKXMYufkkdqhY7vw7slDFRSeGG2QPQ7PX8TGxjN6Ls
Vk1ny16Hqgp7GCfuLK50aUE2MPGV6VCw/VgxV01OiZFW66ZOWQCTOnL3h14sc4tlYw+//gHHFMAc
/L6wxb9DfqKmZi8/zHa59IxwCy2bVrOAEhfVa0fpDf2ENsKEF6MdhGgpBCAyPUwQc/xJoh/9wu1b
AFpjDL8T73eLBLWeeTCMrBE97fE/cQNQ/YbKiXN77xGOSxvZLXHKPzqsIVDBUFewlaaP5gkDB7Zq
ieqG+JX3bNRetrcdXt6W3Ut/m3+pWZaJg2Gu58JZgzlDidSiU5skY2mrA0DhltzqTwtU3NOa0TGE
zaPjmcaRPQRp8SPUv1OU5IZvyd/vOIx+uXjAdX8S4rS4u1YjCFZ19alASizxFMSZAeBcOMs0GK8I
++uXbktvp623Wn+LMKGNECwCestEd2w6Xqz4hw8Zmuz9z4Wd97EpJdY7GVOuKxEYGDYtaQ0ZF9Nh
/Rbh7EGPQqnTcb9ozcoHSuM1+y2LVcK/qRF+zsa/WwQO6gGb0PSW3sJZoGdT49TSlUyOhh0rR2S3
5lzbklD43ZDMeEQjw0skmdYO9ul9jWJJ+3VqDvqwPc/ynbhWKoG79+GDZV48qQ/cl1OhytJCETb/
jXaiBm9QLCuTmeR4J+1JCgBkiRWsWcolFWFFH01HArpgjQXxSY/NkAu+aqdb/Hqh0Ur0m6nD1Eyq
CdxJdJl9hX/+mETgUUZORsdtd7vq8YrVqZBhtG13ACPCQA+4mBzZV8I4TL+9jgj/WWf49Q6LZpuN
bFFAIv1G9wFE3kyZE3GKCpl4+8VT1XlO68ryvr8wtJkk+it3Ff9p3EbcxGsQl7CV0OLzIQdH+TfB
9x4G4vODqzydMuksCNcz9HsQz8Vw5F1j/h1x2Iz3tyHCyWAVhPUfq651J4446XCGkqwnhjm+ldfJ
NiLvnnxYedlLbHBKN8AB3Yvbh1OwgJvii27PfcvgwUn/8F5uaz778jiXG+qAdg2Hdbb9CDQ2xlWF
KyZVMS9ayCIgDH8WKiOAUs+MLaexSjm3Kl48u0NSDAMCy4kd8DwCwsErWLklSOVTHrV65auMObEv
WvxUYguqbdIqG99lC3/Hh49sUZCoHqBzW4+LTDJDFIGMma4Ifr9S+DoLnKocX248ioCyWgL+sS2a
CFiy4yDNj4u+L203hFysE0LmqYIe7cNMGF+tSwCsGbNoUwA3Ti9fwUgwD6cnNceZ03cGmxvMGVqv
hYRqatvI5makb7kFRPDuFzn5W7xar07cGaAgThN1GmuBvgaY+eJK8O9CkaoBlGBUEbtziFvsy4Nk
lmZWSPdYcwmRsA/+KQJkc2614zOumKcarV1JniTGUuAtLHxNwGqA3l+uRw0IA4yGQGxW4yY2WAbh
MYsL0SF4Ss2gOse3+QG1nmGB24YLaIZaJIMBc2AaKYxpymuif1ZdRahVKzhFhFPuy4eN14/qBpGk
J4pBCCBhXBg2MqfvwCNDpel9ssmPgDPFyr71prDqd582kIkMYFsFkifgesIiW3N+D4JvNUPiMiDn
QcwgFFhDzpka/daILlLSUaHOxZGd9yZNordBZHY0gnGqs5SB9hD3FshHR9n11glnxSfHLtWMR1oV
zSrkk0Oiq6P85oh+STsKgA3wHcuIsRM5pKfCe4TpvIveQq0rZ+OAAbWReCsXBk1J5eTmjiQ66MEh
a95PphkBDTPIjMTt5itdboOjNaTuBKTGZb/TPdU/L+fS6QN1HJrs53KJPBJBQjo2B6vBbhbr1X7U
UYi+1Y2j0dKnTlCpV6RtcYSbXra6/AOmHxLXPNiVcheh4oyYP9U7/7XMp/PfhwRF2KIOzk5UAUOR
uZW2fwxRVoGHgvapPLfKKJgRMYjpJr05X+nWQGhj3KW/5rR1K+vRSCmRvBroZvH0EdvWX61NBf+S
AhALLyVwpxXAncZUQfindC3zo05KbWKwgzuKrmrHtEw27xl6AvKw9FVsr+kB9hOF57Tr+1k7GmN1
hrjfsqP9B3QGfAWXO5+H7baXXd+n5EsqDzq9LZe0iIk9PXpiR1dGhyLpq+j6WuEOuOZpq6xIccb9
k1F867KPstU6kgnuDSt5T3mTzrXeQdxABFfKwEaAMIDE7kGx0Z/mYYLy9aMeso7H2hYwwy2qMQR4
IzCGd6rkOjal+jKNepcbtIs9Ntd4Yuuwkh/yqiVu6c0BXw8ISjvA61zVCF6IXyTuSXxsisut9YWR
l4VuUZB9PW9fwZ079jIA5r6mY4djqvGu+ek4D31A3AV9dRxNyEnUgWZxcdr0AGfkhOXCe9m6AR6o
9Y/i67wXZJso70SwdJNUuReuxATgXRNnW2HM7G59+PbdPAoVzzPmj8r65P2y2fXdOkG2qPswRr08
Crn+9VW1Kc6phmH7fl170kfbsC02KO2OVjTfzyBvEMdU9y44x3XhSBfzmRoVXzPR1txIM7mNIOBG
E1GpcDswqYREmggBfD3/1w0XERq4fLEzCXCXjkZsQIX11Vh60WJo1w+6pGf3xCARLDcViZUWm0Ku
njn7Pue0eAMpDtJd3MVYK6cVND/0S1wEv5IkM/SUjBvE9Hk638woSw7lho0Wn7Xq8PB7KdC86Kui
QGDp+mLsATPNkqou4pGt95DeQe3tOGq1ikGK17WfFjTkzsMR6HAVtVgVF1iRJkYJgEJNQWTAWxl0
WtNs+18nBbWhezGsKl+SxMGvuYWKy0pRYCwcPiKIr3YGliTy7QuhcIBjxnoQUi3D2vaXNu/YN0IH
5Yq7HktaAiq+9hbCFUQg5ulquHJV6RiwLqSEWE/m0Xc5GCOCp2F5dKu5zhMqJJIZNJ1xMPL364wa
hcFjV9N/cW4/ZusbaGvFq/0f5/Ke6T/qPyNG9li6ksSM70mwPHD1PmNZGLF0aIxoot8o5Ut3oaJ7
YSJ1Ks7Ug5jkvbhLBAaWgiLw8ksaFMrPAO2Di9hH4JUADGA8RCmitYuVDa5dB1rSWRcImjFuMYTa
jszG0gG/7mv5hfsvlroxKLoPUXsN3Es3DFCNWBC+UigqA4MfBulsTs4rs0NgXSluJb6S9IhenwHu
30D1kwY/JD2gcI+tz+yqH6gTkNUdBGzeKeKwUCQQY8B3AtF4VzvA6mfaH5894BhdUqbRPG3PVc6y
HTELQ4MyNmXUMzTX2VmqMdut7+Rko/7Hon/8Z+s2F67ucw2ice0tINi5y1fkDt3P1za8X+17ZY3/
oglIertkzwLMiP/aDqBcWgPkeqRpYq5zbKprVlZFUjx/5KlXErPR8050/WWTWlgPnqolwrW6j/ud
hb9LmsfEKvINYkKp69oH4leB2vpfi6FnZhXXuAwDfbfO7H41h9Utu7NwfnavdpG/hJZtigNm4u7V
lh1Ag52f6wMXUMo/a3I1vTnr8oNFYJ83gaReeP39cmCt+pVw4VISZ+ADyyxl6MURdYFqXFQ2uy3/
kKLEtzwF1AsIBgweddl6fy7eI06CPdC0/818WyTzYqbceWKa7W6ndWeikc+SWg+6Gx9MTXw0z8Nq
7pIdcf+TLgUMsfdiGAtg2v46z25aWZkx7AB/Uriyo6pfK+y5q5OdmyTq/txrYXprpgSHYgWA/NGn
g6AMkTjubUdyBZK6xEUnf1FesLhuuj15jsTlIH2eHxgeCmaU5QLcG78kjWyFqrmKU9133YMvi0Ei
aBl96WuyeitSvNeQrgYzIkbofqe+kAxpBwenyQaxBAr06GESH6+pzMlzCpfYDkZOPQSPiunUvgjL
TTYJqYDHBQ8Rsv5/rWmWxM2LkINWN5wPb+szCin2PBD3Pyq88C6bdbAgYZ9pQRjHYCFtUrx2v3yg
Pdx/dVgZsXk83BS1bCnp2jolD2jYomZKC/Shqsg8mIx8EBAr7iPXK9C8xDPAt5RmNs4uLJGaigOK
At6E2kwSPM7hngPC+B1xA6o+rSSUph/Z8BgJMe1vxhCa5IRaJje+AJt//+++4XYgmZo14Hxd8VSp
fsFkoN1ZjPizazUbYs/XN4p2682V7HE2Z8zEe+argijQZ88gVnv2wFyx0L3lL+ggdT4ZGx/ux3Eo
cg+SvMjoXT803PxLaW4s0Q3alSYlNz+3ZIvksDkecDrm1v++rtmckL4hHDfJ0Ne2UnjBpctU9b+5
byy9Zelqpr+5qyZFHSuZneBTD3eONGA42UEFb+PM/CPG5jXDRYmg9a2mybABRaEgsL8RJks9Q5m5
qoQS1h9+OjHFz2UZm2y1zadzdMtZse24P2eWsNinHU3bYSWE/FTAtbmeifk96C0d2iz9SvEJ1ksv
tdI3H3o0FJl3o4A62PsYMMqbBsndC3vopKckB383x7+BT0QwPDEc6jsLJRuc3t9wjsaDhh7aKcmH
4TzTN9QFe2IeVElSNKMIJcqc5yOE3+ZAB/sqvA9GBEX0GPkjs+qfEo9D+wmQQmZ5oIKdd+Su5qr7
1PtKi21+g4WI8I4DqVhlhc0N/ygJF41/SR+JIJLUd/h3/7IU1mku9JPUsv3CJ3PoDCDRXzJnhoMI
DRQt+EySOUAF5FI7tjYezXW4zFEjPQ24ufIUWAXPx18U9AVIGh2G+e490fylcXU5+mLCl/Cm0Pbk
a+USmSWeqK9CHjaaF9ioLdlBd5ZSDWppe1dTi1SKaAosCppheT0ilpaxCNM/ZqSrzt+QrKZIMDb8
/2Pasxv24G0UqxBo/MWNtJe2GW/zgCN6niW9aTA/x2yJ6KxnJuLd+aOGxycwj5OGK3V72B8PDu30
luTs2tnFo6ZjSfXkUccQE0509qxrZ4syIpLYgP2NrUXJHKc+O8R/tYxT5krC6TmWpKOYmKunmz+a
56+eW4EgrZSKZaLPvic4ANUrsBgLnpp6Puzuk6mp1cm/VSt79wL4eY1It8BlMi/CKITFMu3CoKHW
LqeCVe/z2odK+HeNZCNYhju+RcTEYfNKzBICgDrjaam7q+Sq7WhoQwiV3S8pRGwE2yuUH0eB3NeU
iQbZWOL/zJTAEDwuQTl9usu45EzriRobNqiBcridmpPsQiNEVMa7k92A8k/aPXWzJcqFw2N9eRIT
X1+7kmQljX9E9R8FmurSBQtCNOm+Gr8Ajc+x31fJYDZeZWYNVdLm7PMILsLQrVjQDTALrUv66+PO
vM0wuVlUZLnmezbPzjSfw2WEjeH1Fds6xJDUe4L39bd7UTbui0olOTBYEkbywfrSEGWWDBwrVzQ7
j9BGvjXZNk1aLCsOKoGWNVTffwqskDDPddVBBp+1thkty+3DLk46ifyuthlEIjlISMcE+mFB2rER
b3LuGuJ6rotbNcNvLA7QjPdaiR8Jm4rnIhtlggxCwj8aTZmK0k66NIkDQoDA3i8vVLwp/Y1DIvET
LAu1ZGhLI5YPkl+a94cSbNWpnWebUEIbCYkw0TmktvtKYQ/ZzBs2R/uUe6VgF3agro64TfpyHpIi
FQXHSpnPO26vC0uBQ42ctQrVGsFtaG/lOovgjm2kBNSLircDoImfB0M9mgt4CgmZ6dsvv5gLIDQi
YHIKtRKUm++FClKKP8LJcO8w5SrRcnXd2tAAzqLQhn/UXowHwCY9e7SRqV51N99PTdc14zDB93Ct
ycOgG873HUgbMectmGhhho7I1Astr1+8FbKawFRQ9w2sTMTfljEd0tCZanEknQus2ZB+1YXf5dUM
Wm0aS08UeRbe6EuDt+6scFdQnmRPMaFWJfU4uU48bs8q+1rlE9N+LkZ/JQhx596qH2qFWeZNZnMX
PyE/4e3I+WMmpA/+I4vaFwWTmAvWKEb0HN1EKzDdT4GkYaZ0p4GjO2aofROKbMj9kIFv5byOK157
FmwdFqV4dBizeegoAcQfbjEdsn9WikpxvBQ2uNw/meK8UbLzk2/pQQViPykjcGU6Hn9vQ4vf1wNI
0O/8WrgkCJlqt1paboQ36IUw8qPGB76VoCoXwt2l7TMe9glWqh0Hw/4R2u6fwepHPnkZZoLKYLur
EKVGf4Zp/GiOhw11Q/K71rfc1mKt9u2k3jlCFjTd5qIibKWFawyjItVJ0lzJM5yA3D1KfYr6cBWI
1SLOhF5w4jnKh05V3a8mMEETBvN+AeB+A7ZBFAnHwTDvhX916Y5hOks62B9n+ACzLXDRC6l/q/1s
AD6Yw06VtCuWCEjIaiqyMSjnMRLbXNNFj9+0GkSbI1SXoSQDSHt3TVkoaZbmRWNmFYh89MkbbQPM
VPLROIZd2lTcVejmrbHPp8ZydCNl1RmYgAgpUKGUESJNo0/LEniEBPY3+0NRcfgKsEHmqSVln3Hq
a94hUHCadtZXbVh34njOw77fUdAMiGt1zMhrMf0aSWyJEgi5hL0AETiI+o9rUPr0Y4prwS2Gk28p
8RiZDO2qztQjP8krlk+AMPEFJ+THfLfsEAUE/LsbaYtevliKLCITEzDSUfJ2sVVaT2GcY52Jpa1M
dU5r8CAss50gpI5lTWOwXEiX7irAURZVjoBTyjYPNFWj9Dov20UXKxQjiBiuhYEVOrDn12gB+nOz
kYRwpa1lMI65P3SNG1ACdXYZ6fW4tdmjQvUIF3nHKJ6ujNb68CnVvT39SlMpZ2Uu+hZBvi2NM9s0
07wK3OZGGPCK7TUZgsUh7TNGo3dOYxNe0g4FaSQeoe2TQ0uq9PivQSivYSASLRAfWpmBTudJziiL
yzBclSiaxDSE0lMJehMSRw25YNVtDdd+2DDeqWg0q4ICdb8sxwRYlbt62geneH6nUDsS3QRU5Vru
wU1/8z+nYtq58T7NIG/5mypgPOFKhPkSLQh4hJfRCa9+DZhXBpud6Zm1WPy+NUAei9ZioPgNWDv4
1hB//FV2N2XGV6XrNXhN0xxtpxdFXFUYd/Xqng0OmF1Ww9bEoioMXHtCnAcyrEKwtRJslK+RRdo+
C/e10TaxO8SjUFzNOc9k0Vyyqj57A5ptnDMIZInle4hhbi/7xc7fr6tlDpbjdgpr6SZ2LmOEBpUL
+fCIfKVwUeu1FJSlCXT0oFNH/Ppw7/CGPe8FyY5aRPjtWxfYb9aF2TUepDmLuLBD5shzswGiQshR
979CzCAi102oTFX5mmOzCl9Nyvoh0UaQpFR5dMcql6J77apv4gmDC5OF+rvCW7Enqshoj2LwBgvi
Wi5wZFHdIzLLsBYrxszXZdQxIdlPv5k4uxwYNCVFE1vytzO0uYLNu2X5OiQKqbESNK8eqrHnZLnZ
rHjDlq9QPkxKT/xHqRaFJtzeDUQ3GZ0ivVLeFNEGyE4vhILgs8sDeBWdS5Yvo6Ozpamrl81NL/dC
YST0jlArxJvC4ERXAheyKazCt/iE2mBO8oNzRv2qSL23xtJh8t+aKWvBB229QDXfe7EWqAWNAn/y
Akp3DLzN9qeiVimYksfm+BPsR2NweYon2bS6JLlGGbBtACqOTTMcdwoeWnga7hnqo7FRKH7G3Doj
J9vfJInhAw07DcIzwEZOyFWpZcbJ3XXA3jzvI/tq39kRwC0OQ5UQHZIYv5x01rw+w2UYOCoFcZpo
c1BRrAGhYQFmqM6+sqfuGfnFAUNScdBrQGev6GEUd3ChH4qqJHzPS91H4LPTjXkP8mGiuN/Nrcx3
udoJ93U8+dKgYarhCkcAwUvmzhjPxyUx+QMtsq15TO99GLblMc46yD9yZCxX87pcjO69CcUzJi19
TxGSlS1svEgfnPZBIsr6PaRJc8X1gJk/cpUTIb5BHoVoDabGZnUujic8geFAzF835Au0NnckbERQ
PNVx2K40qrN0DLleetJDTdBxh1OS2JWoyB1PpF1wzUBzV7EvpWR8KkdisssWiknlYlK16IKrm6Bz
kOMYo40QXo6zePeDCql1WsyfM0pE2VHlFVUCzAH7I9JTlyVhm38qXe9ebnyp3z2hAkGliIS4xrgb
oto6h5HqdmlxA9oJYuTVHKOUQyBwIottX7+SSNqN5shRLyIlyw6Qw6/TQ6STmQ+YRyKguLsPO9ky
AS1MSWLlVqVpqQ87u8HscZyQfJPMWKkVYUEjTy55UpBhk0F9AVx8YbQsE17EO5D2E8TdIHfAKckw
LxIHFXHpzIR58AUjvhNiD92ppnD04d3/Qfiq7of3Uy3ym3Z9VcOF/qesSafidOVtNIBi3ix86VeM
c5xbzMLdyoiYXxEJCCrlEc06O4LSulcvX82/SvpYtoFelm0Bb/3ezLaTC0oUk/CmLGnLctnc15Dh
mymq7ZpwnS2GoaVMN9ZCm1aPP+vT2QXnMleuOeBTMNbeuKVxTPF6L0wKn6hw04RAhxcdWteZsG6S
aYT/r6B1y5G8CZxPPQeJ47p+Nndjxgov1+U5hW2Cx+YX4YdJjiJkfD2nr4xWLE1hfbcXGzimXC9N
NZrHuDWusux7vYsAwRBAeRBNygzbVEUEnIBAkr9a3V6os78V7LY4V3wL8UkHygu1QS+PMirdiMcY
35TkLQFh2lctJRcP0gCanYUxkajdM4Zsgg4gzIe5xhyGjgLvWcmSXA55EbhAmMhTolkrF26lgq1p
DYy8k92+wxYRMRGRAmwqmL0rmjMKUHISUsIvhNb25A3pXXtkVDzuxa6U2oaH77fLWL8HGk2dG3Jb
KNq9VA8M43Gp3/V2FZxDHXcxUR4oubWqAtL7nhrsD9LPdzNKGxVEvhpymehtLaZjHT0Xvv1C2865
NSg0RVCeafxTuLuK7rGu9VSEfNIL4Qm/y8aQpber3DoRZ2QRinwxVgKEJds1kINO88H3AgBQlejX
ZQCPiKLwB5spbk5zz3YZCbMvPyzBtf3vGwvDc4H/YXux5+pXTUpKzkmCwJjfyS7dOmjTbQXhFC19
DE7yU/+PGj6ojIdL4aIywmguYiPE7ILGrUYtEPlRW4IUJ6FC8Pb97QfkLllAbnt00sk6yUu2keyw
Fu1RXXB6PQreC5hOqrhFCk75dyeDfMqJchxlgszZ0WB1w/7u53qzKrMXvLnyKIirdgTCjJ6DscNS
xUH9w6tWg69N394ngYKgjrjGF6StMRunBr0ql0HFxsf7XXLdC8jQRk9kq5Aufpb1Y6qMVgwLYa3G
9JnC+pw30/2qac4LIXPQ70YXYN0P32WqO2Net/xdt1+JqXovhKQd9D5seSoZCZNkNrmAbfZg8IdR
F3UCB7qCKsCWl/uRqwhzM/vL5M6ktQpf3eg1l8fxvgZvQ73YtE5QUprEQjmF8/9+veZqI4FnV+7f
67O3dAta1O9Uo1ORGzCzMUaqxjUAqO1mUzZ97M71SGqFrj4mSQWYwGAY45ZkIkKX0U5CS+CTCYCh
TUdoa1gK95hPZJ5i1TfFakyg/KJ5MOZVRvxxuHhaFSyCLNH4dfOA0RRO27FgD/ixGT9rsqltt7km
DhGhnA5jtP+dSB/5fwPNkRRfAT1ZtV1tTXpGxWeyrGGCj2pzhY4uJYVZwwzTbXuXPc15asCgPNvz
1/SgxPkUr76wP250N4pF8gSvfp4WEG8fQsmMcdGLbQkUoGOJtXuAqGd9+8tAbuj57ri6GG8wWiUO
hjEYjbIbtXntd5ys8o8DxSXcWfVG0WaVyJGDTpPvJiqYzyrt+nH29GtoSosFJMF4KxqaSxXE7TAt
f8mfKJ9H/xR3obJi133UMTc1hIH525DIkTNI9eQe5AQ81B3vRbaDG1Rdsx43J0PBFFRybYTZLaIN
1JMLbQDpQBpgjfEY9nKZUtx/hkOGbDDV4qNdQXDTjsncLIEyKi9mr85jjUMMzPj7F2+WXyICRTHo
QmYq4EwK42qOkMhqD+s3Me+cW5+9T0jDLopS2NnC0tlXLj31fbHR0EWKWJTduvg5uGYVydsn3Beu
vBY1T6JmhZuFqP1OJg2WMUjeAVxbxeBw6X8/m2etOd+QhHgo/lTE9z0yGn6/nzXLqhXBJgXuh+Lm
oBkQpVzB9H8cf+lagMUuDYW/VrJzRHeLluipvteViu6Jt9+YgT36qOiPjnlgUomXqbd9YTCdgTC6
gyk2sWq/laKEHhLICevN3z/vqp24hlbWKhKpPvy7uH7ZaZXKD3XH0T+fQHQvanqV9waLpN/PEGQH
yBlhPDGYIhNoniOt9Tn8gw0GeTQB4icpfEtlQTgEIXOrJ+5kBjT8YoSKJ6X0h7qaLVpJZw0CrY5E
tx4rRVdEid4XitvS/vDZTgZGiiU97t1Xq73aKkvCtzofVAeRMMQlqFMm/gm844Y7LBv2vNFyuvxk
cjnAUit79VQfW/QUKNRubJppac1zMwkYMcCuh2ZPpGZgxOYyDNt1V5/5UVxSROWQkwBsr10KDcI6
R8RK4KHt7PVFh/Er2a1Pb9VBfN7rro+DtEIauZ32qgy4SV7kXVaRg/UeCC2GPhTEd1Mgwr5T1TrQ
rapKstuzkGIkKVnrebTUtipv4/mFOq8Ynnc93jEMfKvuCs1q48RZ8MqeGj40Z2KBu2B6/ISW8Bwl
iKbM1mJmPi0c9qZDDsjuaS7lhfdJ2JwytwlkWmXtb3nqUqCZEth7g48ngLXux6BFwEKn4tFKdAQF
xUV7MQgfxOZaErOqKKPyZH2n3hZHoc8gRFVXDULEsXw0pzC7oe4hF4Zd+lNlkfYNYEl2BfsbKOOx
voQstgpg6/jyPcPyGiyeN+hSDj+IM8tXcH1Gw7ojl19EQLjXBCr9HK2QLmi9xXm/K/i4WNf6bQqw
P3dENgG7A7o1h/7j7TJHLFnX+BjGYMVIaw8m/ZG0BOfLyASX9l5J2R7KENF3fTeCz7bz5ztmc44V
lHwcORGA++3zwaSduT0aZxbZFicuwkGETuIUZujXjPrbaG9jIUt40fcHHSLyYEiHXmZMInsuAcE1
F/QYfh2axw0fDpj2SPYdyr0LGGmuzE53FguJk2yxCCbm+eOZ1J71kTeJvsVbwotx94kpfKcLSEoI
y8Wo/GpbK0WRqLazwfLGpRjM6QXCU37b7Bp9zx4i/eotRB5P9MFiVBv9bXeVDxteMyo08mYB6KK3
VP5tclvywPRHJvNR3Mnye1w8Xsu5ZoTj+V+i5szCEHpCtfR0BjL7hvqfAXJssXF+hE0S2tuBQscm
5je4A75iWjnOYIVL0uLehcmm5B9gpWAL5ROkTB106naLCh7kTWySuZc/3CvDbppm+ZN3MGqsMxZD
PQmNQ6QAVfbeS4laCKg254CBJUcIXUOE/6sPLeP1lhTVCK4i3qNv5Ud/QyY2iCls7XX/HtdcapZu
65FAbo/nTyM2iP92TAqLGp2+FLr9n7fWKSfehHbUeQJWuGlsfXWf0jIlAukH8Pz1OX7pvvgye5YB
KUc3FDq3pRySXAZ/UyhMgJg5FONJO2fI9kxtJMZbulqIF5vXyT03oj9jhDIoP3UFzcq2HjwzYH7d
k4RoM8iV9HM3gsiwjijVIZnjNhjpg+7X2DDUzIwszOPtCAZDvcfGBPcQ3qqxH80ePljgWEsthfe8
pT3QS+VfdDFr7gsQGyFF2j/ifhkLJPXws4M8+8yQwGI2WBhO8iy7gNcmowhGRS6OU045CdH69I54
2l937D45Il1SdO/Jsz6e8NJnyv7zH/SyhwzH6NtZvcSqXFHoe9Yg7ssH6U5WKtP8GVNvsuVhHtcx
kzlCJqu+0wM/isEV2QERX3ZSwth1lvqyi3/5PNHbtk6N6w0ToDtzc9txoDCKPhgaxV3RydYOAEU2
Kko6Te9M9lGIVDUfU59ABjDPwWqA5OrJCBTnUMhUPos1Mn04jvOJdUFQ5JFZdKYzRFAPlTFY4Eiw
4Y9CaD+Ec99DEnyAVW4PLwbn/9rXDLnZkk2BLKX0yzcZruHeVtqzfiZvTBuuzRUywmNXhbExVYW3
5NRIulBz8Td32+f77XAwawR/bgEF40mHN4fR/N1lvv4JVDT0rRUVlMFqbrlI/ZvNHZx4PM56/ikY
wROKJqIZijjSkhL+AsPrQukd3vyF+q2zcyjT9JZX5ZmAdXLn1I7ITCY9JUIDHmZzdHtNuTsGtGUx
FVylqVTlV9CjMkX/QKnoJqWoYXmHGDzC8KgYg3PtiZpSE+F1q3VmIlFNucfGc/1AEbqzUmjyPGrB
TUsFa6qG7Md9hEvcmuItHzgi4O3B5kF6JtH79uhMEVnBOBQ/N6IOvaWPAOoYcYx+YOQrL950Q4B3
qkKbuWA6KelpGQgwi7WSvS+npjgTtzhRhUQMH8L2343V/T5PAVPKR2Y3J2OlNA5Io38ZeW0YVBhx
lS/3g3t20cRQJpTyRt0T/O+t+IoQBQ1RteetgcjLmxlqAfkSIulINOhZfyggUChtvaUrJXYMr04d
9n73++V8E4L4Q8jma4XfvcuzBOOZcxZaJ7+PaxtHciz64srkfVE6Hs57m/UTQci7cGxWvjM85NlG
Vp3rYoMU5D98uzWYrn8widNs1jb60pfSbZMSL9Yzkgkr61LYHhDeHjXjDkiPnU+Za61+lRIgqftR
Za5c47WUVkYEele1M7s4g8+3S1K7z7qTRivAQVoSrOH7+dT24O5V2ItD41mZsKbFAB3wy+15QUF8
EkLAfsQMZC4i07IJnkeBje1MGI6khfvOPB7N3pvPPGeFP5w7iBRzRh54ZfMJmTXQWinP0FTxTr5i
d83zkWS1Z/7C2jtVfBwMnZqXyTkXYTqz/nSRcughdSU8DK0fqonxZ4MDA4OSxNLCY2Z/RNytbtCy
bBeathHXTxgCMe9RaxzsTrxQJdVtI4mHDc9+xWuZCTd/80gLUG7r3pOFiCmXle7KMQ2BvQ0VmV4R
Vuh/lAE2C0rlVyegFmKCLcB7IrEj9FJtWeHnEilJEczy1wBVQciJIYUbRI14GadA2YuVaJsRobkp
g9ix7QrmadnOBYbh2PHpR6A87KtrpwKqKnEimpUhAdu0hH2HXLx5T+MKwbJl9CJiMhW1slxPFMlb
hvjsu4TgkuAWGfu+oetPgRHlPaVMkXcF8PAII3azhXGYnzsBEgTAvvJfOvDgfiDmOtYnjcOAsFe7
xPUbvG1kF71ZpKHKi0NTvL0cuZtkYJoCTlQNf077Z3YlrsfXWrwmo1hv+qvrzLODeGUEXC+q1sK9
D4CN+IrgfFSBz2IO1VEMBSP1fuwJk/9usc31M2izMNzyoF5ET6ZXBFb/5oadYI1K6xkJqOCClI7j
cy92nOc8sTyUoYhUJ4uPWbBiJnMAHJ5XbHC00IKSwwJaq39U1Opjn1TbSMyvy/bJuqc+T1p836Kr
l7s4pFuPoj466HdPbh7//XFjAtpOtVC0hXSxX9VuZ7vX/7+hDBvIn1/nnTiv3tpd82PpGjSRIwUy
YoxgdHJ2QUjI87ssEdY5pyg17GfXCsePqpSn1345cAIrP2bs6gVVn9CgLM5tQwnHHl6GHqtuRuEm
FBqWUVYRgpT+pfjbNTbIiiDxP2H/aA6k9MnHY4jzCeCTcXeyGL/k7BWvYZ9B6h6sRpFUzNdzYGpi
sVnsBOmRWacsI2YHbmLjxKl/N00fgB+S+ENawJcAWsqCq7OuRxeOnEjb07WFKF+a93uzDQp6PvRP
HmvkBvLLi2IUvoY7+yYuHJwLGGuaqFlB4hZhOSAttBrxE1vvCHcg6vILAmS4QPH0OtHIOq1oqbpk
Ko7NlxAkXpxxNbKkKwJaspjvHmiRu1htMY6V882f/DpFkn5zb4eVXrNFKOuvXnqaWCw5LfhOX2s6
7zvoWcCW4gwqEvOr6HVosM5Zx9Q2IjHtGnQvNRuJC8jPswjj5jk71h78Ww/tivL5B2uIBvkzA+EH
yB4m8xq69Ygi0nMT//RtXSTkxojDKLAlkPmExoY3KFaOUxmiTqv2isTwWRF2ZQMnL8JTXsXCeNqb
aEU1xReQxLQKiSnxf6yivyJSTnN1t0hFdtTHE18rqiEtDG746cb/lSnvkgZke478eOu6AE9j1vHF
S+rz3U0raINdf5PKL/UiodMH+kFPyLEVmSa6BMTGrV1jPqfztNmlkJOaNPeEnl4rQc39gx8CUgvm
Sv7ap9GDb2MykwHithXBvexYsbiF7bPQpN7vCM0Q2eceCR8MdS5jmndDxe+FfrjeUjUJPUFqsV1T
fZib2B4ee/yAqdETLT4vLhnZcRYGzjFiWIK1bZVfrXGwsIHy2pA7PNg9LyqPtmK8fchAt59ctDUX
3uGd7DEKsPMn23hr1UVoSrAjRDkFaokB5bdgd2hAF7A2NGb4DzBiW1+Amlc3wPuG+PTZDiFU5MLY
BOlOw+tbr6jFqnM1SEtgpllJmFLO7mTs0exIXBI9iDxD3Bjnwj51dCBz6Z7pZiPtjTT4lIvkkCKb
jJK/rhi/9cL6MxKhlb/XaItaaSjApB8T1n2YD4YVeAyuqMsfBUNs1mYu+gIyIqcYZ9pU/8B83eFd
zJ6GJQ2jT/DCad5dAL38t1DJmr3jtu+lnjT3dPI1m99QpMOmp603d9KKcnOK74iMtuin07gfm/Wk
yKSASlaxo4+ya0Px8wCZXPoBWgEA69V2ao8WbWsN62L0kirvphovYy7cBlE/Bi3Ch3E8SZ2eY8oP
gYvXPxFUm7zS7MJkPVxE1YqfZg/eDFwUbHs2T3xl1JcaxrcDmQFqrUvsSZclC2K6IpaoJuBew+34
xwGI/O1O/soGChgCmjJ7buk8eStWFE1+z+Ep5trlHkVjiH7Y5CcFNR6xLOo0mCC+reHgYEVIwrQ6
llhSk4KkqE7e5FRyjsQT9IS+TXIxdjz/OISHovrDoopt/xU59xAJvrg+u7HpPAo/5SUKGztuQ+r0
sINZywIVT0R9MhyaWQXFjuz0hCZA6It/J+eilXpR8+UzqVNAT6TXof2TtXTKwsNfwMs5VE0AcF15
yIpWvQ06rsOa9NFIHc1Wx6AiaJ+8OMUza8ZBhXUjV/8BMQN7oGQJ2UcLwO4863rGytEqUFVr35e2
7tW4swNQul6avo+XEhvcxkcOuazLX2ck85PUQIgu6yKY7oMhlNhiSMPUscBx4TQhSvu4lYdeJmA4
0t0k5muchKUXBziaH8Zkj/cSyCeAENae+EKOuZuVjCOpmjZiaq/s+DgNt8bJ61gild1f4zbzumdz
YN6A2r5ydg+krZqdM5Qx/LtCtWhceK08R9r4vvGQwp52qgXGrwZGe4CTc7eRWvqwiMKzMIA+q6Jl
Z8n9czGe/OechYHUkClhKTTnVx1swRyni74KHcnegEqe3AjTKF9MiN+DI1F+NQzPWFs79KZXaeYC
fkZRA3Ogc1rFzksqIaGQt4/T1NbCLThLcAf89vKiIuXakEmNHocidA1a+BcNwIs6LWc3tDqcTvOS
pWFKzSbjr5xxLbE2LlIqhkGfaZ0/2qiZaOjH6vKACKL6/HZM4vtTlUwz5si+Mhb5Nr+Lq4tQat6f
IFFBGLRCObqqnn5rK8OWM5vs2DfIJ/DoYfFRLJx0/DmPGcH9GT8rMDnazfMx1AVhra9fMb2+bK54
Y6g9GKNE3jOZZgAEpe1xYyEteLJlU4vg28LLqEvQluSTr0he6MtjEDgfmjrgOQcvxcL0CC3kf2+/
/u8C4+DARvt2Is5g8IgknnS1kduw67rTLjyg+GFtrfzk4F3RRGewSxHUr3lUCDHTyN6/36DBjP4a
U621txDM1p9G1ecmfytRTR81mny6IUgIIGj/fbY3RwWsfRL/k8FEktIXPy+2TVVa2v/97jHdd0VZ
+nvhYNT6XlVp4DBa0AtFcTUsDMDU+rgWgwFo+2+iwCu8kVkle+0Q+sN8AUiLCjsGSk0ICq/KR0FO
qvD1EOAlmvmmyfEwf7gm1i0e6rFCcMw0wcUoU9LuMmaA4FH1OTvx1hnDZBjgwIks8DBJwxpJKYb7
17CCiRKSFNZI3YMCzEUpD+evfiTTIM3nTt+SsFpqs01A1wCCwWSZbRknsFaIZA5hlT2HjWoxGz0B
TiynDCQ/SSgZQj6OkBDqD93ZzuwQQfw5Fb/Ce8dtNi5LKWUySnSnRDivcuijgtcQpze5PIHJ+izk
T3akOGCjZAjojMyKxdtChz/aZJJXY2Vuu6xC/d3i2iRjxzGI3t3oqUKTsldYBqy7VTbPJynMBNr9
DErpUYLRyD4ISxcLAPhlWJtcjnxGXyJ4YyoWfdvaSODou29/eRHfZSerCTvyTsieBZ2h9XUwTb53
s9rYdUqh8RlXK7hkywGas8zj4vcrdlDaft5HcvMsGc8rZL+8/qlPoBLNMXbZQuMdaw/LBUGXXFgP
PIp7wDfA7egMSaocT/FexV0ElnP0pMeDOcUok24i/JJo7RAT3LakS3zdt36TZZIpM0xTQrHRyIwW
pjfJNDDrIh39ibnF41TfMvtbezfvrow9Fcg57rFn5WPojBJUXUtSqP2ogw6k6DK6nEUoJnt/CDUz
oTQU0QGcXWQFvr92GUt+kyorOtNUf9LrUtBo8Ab/VZ5RO8Sx6y5CMw8QYYvpy+iCAo4DZZdb+IhU
mmyknSYd3B+Kbo31xCHZ5uFduu9dw+ZZoJ2PcPjEukznYRI//gkqvSxJ6kTlAd8p00oodhQq7CCm
r4HLKMHs8U1PPeXSY2pkTyTh3RJ4S7m2st8KADjLUM49KTPy5+EVJe9eHGFMSL2OESUl2rnrgpUJ
2EesYvxDIzAUoOvwF8RGjOxpFsUup941vY3/ujgkA/s7/GH5eHbc3wXi0/WaEmE+yK5HbW0XdfEn
EZD/UClNF4I3Zy6g0nVOlq743EgCAzyRN4y0xQWxAxXYw1oYRHgRbOQLYT7yn59y6L3DVasp6jIn
JTrLHIZurjrmIHVLA6XMSTnrWNVn4euWzce83jqnFxzvAk1h1923y1Rn1rxXg08lbXryjQOflt1P
yRkaq8C5kV/cn1NdVzHyMm+LmNEVJdaBziRVfkquie/cJp+Z8HxApsx3vpSgNuwcMIjU9pfl5QK/
JRMA3A+lGr3Y6nGFBhevyyeO5ZUMRKCkB/ooKhY81Bmo45T6XFAs9vdyokOYILvHmbZUHrRuePWL
qkxSpAnHPBIREUO5EzqkpXOXJ6KWImXfuNPn8YLfyqGCFqPxk9L8F2eaihWcB5+NYhI37MHOP+sv
ynDmW5MWG98WgkWnPI9Lu5BjIAKLeRTiXY5+QKJdMTKUwpfO/qNY2x2JwcwLLPF0hXPB9oJfVKhb
d3/rcWTxzqViIPitWhvpJdiP7rFmaSu/aholgCT9aWBY6l/8R0DsDyS+hxA/RSAQiNXMdGaayN2d
uxmYMADfDQy4bj3sJ8Mwv70XC+CHWpveElev61Fy1SEIVMYnMm4l6hRInaDwutC9oEhvbSGtAyG/
/Vg9fKeT2cDZx+4VgktmM2uqumAVkuaTyEKmhCGAjGiGF3jxmkYgXMFgH4nyx9oQz1CX23uz5BTa
qdG/RORbj2hEnAO5uL3F45idl9dYNtM7iQRzL7tQB5Mp+11Rom3W6fg6ZVjSBDywfXk/5jxsjC/w
T12lvhkmU6FcHO5rJNvxgs7VAUyENLsR1jH3uQpbPIyjBGfTMmpQmJo8cJK+pI9O9QVizXlYxMoS
Sja8Ld7JiDE1FOJQiqC0oB1wK5FMU2UnRv8mgGR5BwkF3oXzuTxiye0tRwBnapd33/3n/Hg1kNWW
eXSfWBr1CIBL2OR/+Y9u2BPuJ2rOIyJsuUpU1PnPQUjVn0ZH79YvrGp2eaYZjhRZvgIQsuTDtjHk
8VX0JtYUZgjNAITuoyyH1iqaBGa5JdQ5O/jh8MaPn1FuMQ4q0qnZOrDMyKXy/sNRRbiSDQPx3pUq
GspNguXV3weIPbiyNhIXyeggq3pXyB+d/6bX9duk488aVZQbCysuy+LrObjPvOl29Jw+mk05Dn1I
ermDQ4r6iCbfhZ7JARhRjnrlApNqvGSzd/bRdIt3gOV6zJOEwpH9a3BmvQmCH2ToX3tQeTD3Uzsz
nB4Smjm28fo5fjU/KnuAKbw7W/aoiLDwOmgLaH323W6Yxk5Pwir9N2XcDuSplTBl012WjVxy5CKx
6VBXuMKQlHr5ak+z3eIhhIwOE/5ZMPr5xXAD5NynOque6MOAu2/IZLoIXkVqQThxtyFZnbrbn8ji
Ucyl8UaMuK69T/yWHcT16aYhXpql712oap4wDPesGwUi/U8RNdSwCt/ynD37Ivr7k9FFJ8N2XQar
bovq1TZgLA7vLfLE6+7MxNnZ2xjl+B057fgLUB3y1kiMiCZaVCHfh2sxuevk6k+L63ZmIIMUbE60
dVV27aGzM83MH4M318bCmtXvLtNZbgwWB6h2ztq644+SkuURMTxC2Cv2ILxp5/kjOORb5luoVItm
rsSOnYqx0Mm/VnQXRG6WT8IJ51DXzY3TAb94h7iHb0njj001uWBH0RLGahjG1DmrVBdc1jcl9TLf
enZdmuED2vZrB08m4K30wCpr+ZzeBw9Z0j3ZAURHl2zc6NX8ysmykVI3uwFaNgePSetf/uPd2pxQ
O8p3Vy154K1BdZc2gScQEWOCSJGY6ElJkmXNOJ8tm24oU18nNIzCuBpuP5joeIE2fq6rfOVsLF95
j8dNnJ82DtQA4mCtb2I1Pip29jOaTe1JDHUrkWIJOWXf8JT08vw9Y8qtsRkozlFAKXiNLpM8os7y
kZh6lPSEds4KdFrnpHtAoyvnhASqRWi18spHWpsqTrpsehDxqv9IOeZMclMC6iVHe2366wfXx2S8
jYMsI4dSUrJsEaLpuqFc6CeMoFI49/L6vrK0IYCNWLird7+ZVup0D/eEzM3+OAzSxxjMgUKecog7
VBURB/81Tlk7dIZWoqT463b+g1rkT0qi3xw1S37fP7MnljtnqMYT1ob159hScTHWyU77UxvQhdY6
3j8gaMugc57BSanzy2BqdVX8lcLMugwAmo2dRAvnpbJgFz1HlP97K8I4RCpewjz3gfpRpP7oD6pT
QeR/JuzrtMQIHL9SX+IkRUZElliBuo5GAqKm3e9dYo5OxX8+qbhSKigwp2VXlk1PUpnyg+Ox5t6q
cITMsbMTqvRmea1hL9gNbKYpRPertSk6hJJajTzzb/WF7x1cKHqf6MOpDb70PMj9C9JDlDxXTlXw
Zdv8o3iOyw7HUFF+34UpZ73QRsDOJ8rKl/q7UHKtAuQXJpbKg81dH+va8AElpwVw87D/uNRp4GT4
qG12FcAd4sYIBXsvxecvADhkPX1DJaIRWC7rerb6mJ5YORKMv0/6RgHPqXRW9bpGG9OtxYUdQ4nc
tJWl5BBP+7zuM23a0hnV1/kp++LtkoztZQka6LhQ9i4FS0hlBb41dU5Pkh/FipNELVlDdjlvHLSX
OrOnjEA/bxAcWMi9Ew9kVFZ74c1y10hIMXrM6Of1xkAK/pfpZQ2lX5+1KEI4Co9A/vMk1Ny/7V+2
CGoLY5OjTnFvxtiSgTVeDdO23ZkCtLcMpG4oUB9Om8WdA+rur5wWP/N04QJLLEqJR+dylLxv1KX+
EBSy+t1EDTDP1NFKEvhcgoMbBKYY/vLdS4NUVN1Ov9VNJYuOF89VFfoPDTseg/+D+qRPNns/jgBS
D4VyDiDBupwPiPj211yT7UX4WDcsdSqXh3/qSPtyseY9BTDntmi6gPkyYgH2MTbsIVjgxjz6NBTD
t0nQeYmXUGX+p0LjqR0rzV/VVYlr5HIx1cFuheY3tkp19GG4yxYUBdt4bSW6wnAGrujQ0f7WFd6s
/TqcscQ92PmpS9WSvUIW3UEfLMTRi7hyZxSoLgrJMLd1eysKgXP/qtxYESOIoHljhqOBn/Gfus0j
RcmZ2MEjTsFq21UczgFx/8ZtaAjmRdHhsmAPjoBabwKoJAzRrs12D6N19qcFZ4x65s5wg+KPLfDP
10Zt7ZnqBPdViCGu7zR1h0jIWe3CzDzeiWJ0REI5jhWb6kPFXrkQJLbsMTxXjI1ZS+1u8llVb1Gw
v6YRwecRYYTA8igJJoZEwNJp+RfW+mchmHY7XaHda3NNCUvCHvpBtJ/HIu/dEBfgTJIO9iZ8SqrT
8KDWiGV940l91C1NnU6Pe/alSz4D8LWD7ydPugl9de5MfFY8cGQOIO6YEgLYFWecQjVOz0MCHrdF
v3dPUOX201fYsHB0vrYRrAqS/1nGZt7RLiuO4GQhtV4s2Fty5/EXj4CxEbzC4nybCiKa8uJpTxXV
XD++mp7lzVp01vSBVxxGxwhUf2n+uU0lcyDMqxaPSOwUpYvAdqGglejDe8DSs8SfsLQgLyU94Nem
D302KUjZylIIFVPcbn2EHVdTnEtay+0H3dRAh5+tuZ5Q28p/JuuDPZ/lOSl+SEFHSVWDUTMehkln
YHJnQQo0liNunH8T/kBprXKrXyIG/lapBAVbJ1ncT739OAC6ICIhSIXHyytFLzd/AS4z0RnePQBY
ctN0UDXYwuqiAy2TIKHK93e01imURdLYU0kYPXMLWb8GA3krgQG0mmltPEC4Wwby1gADHpAH+wos
UMPOSZPWb0JHzRjBRvf2SLoaSmC7nWTm+C9kEe+Qm+XWo2sbYb0kRERufK7SvbksXpSmlpRwZugX
Mvjm0i3Sr0aq+j1VoVal/5fKFtGLfNx0lxWON6fzKrmeTN97DPmwy/NgCImqlBwUCwKgMthzt81L
NcV66slKP0vJmC0F6hwamBfYRa3sRoNxxihAFxep9v5GaYBkNYjT7uOo6Qo6HdTpp7FsH2Fg511B
VOmmdLI/6+a/rbXU9DDHz8qSF8cJ1fEALIfTfnFhYTL/ctru1gI+gDE0Sm0Px5yPf+SwbxsYdlj1
RQtVR9K76Zr9Z3d+A2L7ZvYLcYoWbsPrTSkITXKPEQRYtRRHM2LQ17ZhRGwOYtU/YSt319YxHnic
MmtuKLVaUQMVrJ02We6MdyoU5bp+UYPRJi3hAiQYIgPHx4vcPS/UMo/09b9SITLmRpbX7mfYJ0/v
lwPWcasUefMsDeISFG7oHV7tURtc+GM5PPIMgKEbqkVssqJF0NdwcuZzovLF/oYqmeYMwHDcXtwZ
gdps0YUFzflo0G9SxP50b5yn7r/ScikVqpIt6JZYVac8Rf8kjiAPMgYZZQ9g79a+ljP2iCjEjVUU
+qtwP0bFtzzV9kYNLhgep/QUjyyYh5h5ZwU/JcHNMNUIk6FV4Qd7caGELBPQot/MR3Z9XnyeCe/e
Xj7jpthZTz4/WjAU23esw8xeZTBxbqxaeZIblrfNGi8jjsPQzvnFfMpTBo4LJ/9l5w0ELXiDZwVJ
kgbM/xchKFAP5bR5o8816XkStoKz92M4kKrGKsicvpYHEc+13YD6v7OilV3+9zv2GjNDjf1c6HZW
8c4+kOjvJu0rSidtCsQJeClGLhMpkPZmz4gaZfY0gjxT3xtwQtmI8VafL3bnldfPe2Ex1wCnLtGJ
gBXGa3dUAPhTFLaPv5RMlPrBerCu5GTpvZpLufliqmwUKYleG2VPcUlIDldWsMij9QUqMyaNt275
b4vh0/34c4vefpcNp0Q7NF6h2W/rzv+Hp4mwp1NehMe+1rOiACrpywhyeQA6TJmH/SdlUuCrZ/K5
Dru4pLAeJQMcpZo9i6RUUJobBRFSouT6lWCfuvK8LK1kEz8Q9VyxMvqEEhJ4AAdjTXUIl4t52+vd
+VDR+QTWv1LJLsbfMmyhlly5Bz1ZBh3lXx97rJuNijk1xBdEZyIHyiVHQYlNP2rdaA57axlYeZD6
0bdvn/uPrDhKH/y80fub02NWh1mP2HguyW4M7ZrFAhqf1WUyjRKC+0bYzWtLpPuWv6cqW7SrVQXB
+eAZwGzixYsBVypMuFtV0Gk14DmdyG3iWwKz6YNEvr+RyaOHzivX/CRl26yHO7f1yoCoGvyH24Jv
hPGOJRwbOnlXCX0yXVli51kBJCW9IfcYHxMADUtd9GEy2PpN8itA32ZRWVFUnUbSfadkLz+Gg6Yu
Nicf7sv2LdAPRS8Ys79nVq1t3xBxgMqrIT9uzjdhV+hCufVfZS6YzEPbFqQDvtoq3Ciy/WSK/xws
zti05J92KcNQrL4DSF7XkjOInTXvvufFsJVK9ArHL5wNR8hjlX1U6gU0/R6qJJYRgmssyJXS8d9c
Oh52ZLstO+PtAMcxKOcWqrcTgnI9tmWdRlifVWGpT3hIEBNKSM7NS2OqY+avEuSgugvMX4gMLWId
IvdmLi8vMoCoAdNmuK+VzdvKT6XIQ4VALlWJ034wNEBueG4YCZQoKSdZAQRsHOG7gz/IhArEuoku
Px04/ixkmhkLxPXb5mwjkuAplU+R5jy7694DEYxI/vjrTjslqngkJjpF6EV9Ay32wIaHety/yRrQ
TbBiD8axhmLqsbXqecPY8lUC5AbZnr5v2QrmiGFhbzdlNMa+9ayPTdjTWQGDf8avAPObxujKX7sJ
r3k1cyBXekcC6zkOaIx7aAoRkpDlucT9CVm61zX1KOz3SUMfObB3IzrNg+ZyjvIgUI9XehW73m3+
GRjM8fLJPbgxSw4nP+1UQUJ5HBynKd0clJZ6qpnh38vtzxGjfSwnrSYn9CnD9J4vg6Y/hKq5Go/v
h31bYosVLFP7o829ht7cWoBJxPyTVBA7VPDKGePLB8lmz3/VUjEhVEg6aft7vDLSP3x6Rn8S8OFj
s03EeGVWBrRTNBe4lAuIkVZNqomBtiyW11GE7BZZuP0jge8NERXAC3kSNZuUxUSSiaN/rTRkRDK/
17Y6h7E10wJxHxm1cMtHt0GX1kymhp04EVDYiLZkLzsliRYfOiS314EanzhECOvcjZN9MSisofpY
0NZbgqeQDGxeDUi9QKes2aAvwDZATElOZiQcZB0uP8dvyuSiSWYyIB5dpeY7WDvE+dyTwIyfpFrf
KimDzTryd7vhtUSPWueIR4bFXeYLPvhUSlwvoVXNCvVf/m0UMz1Qkd4tLSCCWdWHbLVHJ9CP3Kl1
MDqXPU/YEwfUcj8gJRBNixLUW6MXPFwIIGHZr+11Vffhswm3GTgOAr8+MMav5J3d9KGAuHmzoioy
rcMv02V847vyxK7Aluy/2gppMQdcDOAvHBBP1MPbBGl345BAS9x6RlF+UXyjrQKWyxJPQK+ZTfGo
FVpNVlf9mDqOJPcubVzDvIqhxN2Yf8cGIsRUALnDOzoZYstT6B8E0F/cHA6xOyXRewNI1tv88ZaL
xMAYGP3jLdGoSBf9caoDD373mvICbvzXGjeX47U3+EGLtFJxL2wsxO9LYxxMpq8P+j6VVsQ+BHX2
g/2LNyTjsVk35+Z3FnjpPRHPSolO9/davb8kOVWLqT20pg7BIefMsVNqZzdrsWMBLARwJuazgD56
lIT+N9UtGKndKF8LrSGtMLsB8TztE1x3kKZDNof1Yc3kFpv/sdkjWnT/hPf1lMBDCl7KbfbiDFcs
/Oln6mEyAQTkrprqRJTmt2on/yMjhwQo+Cn0ITXqeWA+Sa20aR3+Wp4Yebqc/BWNVKqler/pb6+T
x1TvYoqMENenx5LYmcI+Jh9HKAah5XqOhzYUe8FuFTDRvMTj9W3N8Ih6LkplrZs027yEtwgMp5Py
hhoKm7J8nZMbp3Pm74SUFTRsUPsutWn51YKqUK4vPEFCdTEKl3/P9kmkd2wi75tCK1wwwUnzyg16
kEHc9wNyHdxxalcmbtkw9rOfmGE49ruCk0ztZOqdoQGwxDE4Zzr7K8CC8PD/y3vUQNf/8sR3fspW
5mfUQlFZWPcwUYWpFvn383tBfw6F6dcYJK1+oY7bWeCuhyvwZ+tdZhsO31jeLvdkpjwPeDl5vX0I
7AAGluo+AeiaDd4N/bSewDE8N/Ltaxn672jptuymwC4Kl758YfxQNDtlaPOaDlpINGh6MCCTdLif
17ZRVH5oWHlmUZkkuFNTUGBPMN4efT5rvb93vo1DMUuy/wuXm4a82dBZy2hm75Nb91zXSRgMF7qu
WDzs/iLL+tGA0nTP9RurE3ltJL5doJ3rsUe7VNdvUT7rO+RF+3YrIzBvXBfB9ALmtmg+KNoA4HZK
bc7ITL4KvlapUMWnXSS+FwYZrjBnc90QtG3eIDhRfOLLNMxXSx9aIBCm/XWTqmw4dU7+uYIdIjau
NmcZURrQlPMxyjnZCclYdvPqPvWO8jtMjMmtg4YdzWbWdhNUhhbL4nWJ0gsgt699+f2WfheX+U2i
ruyzQRP4SQ9LPVgenSECjxuGxCui9PVY01edZf6kV1SbWvofJdA0T03H17xUICJe+yqArYvyKi6v
qpL9i40xEM4N9uJ6wZUtpZi9gipFQs2UOxlL5TqwK4qsMptkz8pcx6uS7H+Ua7DjCE6OVOzp62yz
smfzrJhL5lNDjAg8OLAS0HV7JW0dV/QzMc0B8XhAmpQ+0xvsPG6VfbyVqCUZWVCDmMAujJBdBV+r
PEKdORYsKgMkf8qG2h1wo2HjNaFXHZKT8mxraaDDexmbrKzaV9rZ7opng516DKU7dsO/NsGAtCLB
5mSP3SyRsrZaECP9TA+cGJC26ck7of7WGejeTIbWETCDjhRtpG9+jw+8LfjwCbt4O5w3nSFgkGqQ
goEsc7s5WEye8bdsgU5TIt9gus/7cKjTjUzIcJ1S5o65rc5pWL91u/tbyzP6vy6oE+xA2/AKk7t/
nQ9GanCSmcZaCxGURo826NwTnd56xCl6N8EEU9L4u60ef61IGAvpcm/u4XZkk8591REKG1K1hy7X
mpFcnCNzxnOzVtV/04/DjDCtK+u0PDcyCIA3jmE7g2gezHAAEj9BQPJP1hAl+9lO5wzAphFMlHZ1
BJEfY0x/r8/kMVob1wCg9BD4m3tKQvjWgIqcUy86Db7R6psxExMQa8HXR5iL2AkHz6jPR5liZpes
BACKJiczpdxVxdBpT08UI21hm4PosIaERVnePJy2Gzdxgf+VdsIeTblUM2QpqScQ3VoPoai3Qan4
MO/PRod4KaPT7LorJ/XwICdClw09Ez+cLyp2KEMqK3xB1+BV1Jx1pSfmQ1FyOsfBo/ITrUK/gadb
p4ZobP2go6n26SF00Z93ws05J0A/lO+CMBotqXIFQXngUPNfYlebPyZT6fQMEBurjvemUas14Jom
TZiNDv1u9dlbI5DSgWBerl4xFU2ebsqVTqBljzbMkSEtrW6tjhyB8LK8CZBKFd9RcND9O0mngWAN
CdQs0bYNz6qrJWzpClbW2013ISQrbVusroMF0f8SN5ril4vjnF2CKAzfwXHscDWZNULSNK5MPgCm
7Yfk62IN9YIT8rudZpkdJ3J+XWsvTYEz/E1aCss58MbJhm7SvbMYpIgPN0rF7VQE1oG92qzch0jW
2k0JAkZ1tcWbKguWbw1+o1phaZqBsCBxxCu74nWSW46BwdGjj9apb8N/i2W8OMsmZpvRDNC8dCh7
aBV8V7Z1ulJ6FV4Qpr2LXWn4kIRSdNx5lryYJdJUzdiunygMhoZFXbmyIhroayDba0Dk55YEhELu
tin2jXUarju27gM1vEKifHJGCeTUIK84LfLen9wwfvpRKblRT28BxY6dniBLHULk8CxTGLUxkFau
pYkYrH3r0GEdXUlPFJ6utAzDJdI8I3iTA96ZxcWbMyyQBE2diOQfTgngXXrsdQvmn+xAAiRukY9T
D2h721enaLUUbQYlkBKZuVRZVUvkdfnA31OEl+HTG3RzJJkQ18MHsXNsB9jSQzYFuMtJd5FValcO
GSPK8J9thKNY2lzPngYLjMfmPCuwZvkqIG5dkobw6LJdniMC/zDigA7CYAJA6PhpUtved+kBmH1H
5BMFUorQrdwQ6ohyKq4a+T6UoV9GsYWqWpusDnPUk6LabAjTYqj8kN6N/njrveB3uAYEP1Npz329
UZXwcV+8qyVxwk0xkf4HV1rjfHCacq/w/w67zFnAyuWsNvQeZycDjMHIQX6dBRI8XPWjzPp6AZ8+
Ubm3XUooKz5TPOmsy2RQUXG933X9quP1L8ZqgZIfHJhfovzT7/jypQOfn8vXrvZiWLgY04iE5RyJ
VAy5jLAGcHJa7oJQep7RluHajSLKbVJdJNVJjwHUmxinA1LnZ/FZLDLmw3qmoVfvMpyKZ1XPO3G6
ehunzrh6hg60i1JtriFJzKjpDLp5y6XBmNKdITKOlBrpzaVaXVbhDMzB3p6MveU//wrIuJ/vId5W
oH5LHzx3Dw7WZ77mppFrJp9K+LeK56uzppoZwFKdhKpFKnThBlRLvQyp4n0mbYRchqsrJLZVCe9U
+lVwczvqvXKiU6fasHSkDZv6eE2xswY/AyYcVtdal0AirbzgfhfOaZdrzEqsgCXXrLE91MlP+YMI
PWQYxtPILbE+WvcpkEWnxV5YmhG71aazBEgHlgR5SpGXwbc+KGBSdAtc1w4/XT5krkeHsxSyumIW
YzJ0U+Ika57v6AUklojNeJpij81BMlcneRrzRMgbZbPymm8F/n7EzF4gHg8OSKBwSBwH33mxtkHX
Syr0okivl3A5cNuvaVhBhQv531qpLqEfLQI5Fl69LIRQvWRB5j8ULCAhCn3xGs5pbBLpHoM2saUB
JnA4CAcMCV4C4H+WvJbz7bzyR5zgDPynRn3if5fvRThmgAZPJ4wBq/hmDvVBsb5QUSaBWIU+LBYg
CUJjcdNLl7QRehfDp7R5AAbROeWgQsHGIXvsA1wTo6Y/+PCkl5EFznCVdvA2syUGgyeGZiBCoh2L
wybgjhGIueQeNnhq/o1y1dS25meT3T9c1dWNtjDaxvwkr9k6DKYLwb+iO9h/MoLAYuDwXoco5FxW
zQ6PiQ4QlwtdL4PAmj7V8YYlyL3Ob63mociml+MHh/Oc7S0i/69Q4YXfPVD16GGJJuLHnLcxsA7B
BwACFqEeNS3KYTuiNUCszRJ8ix/Y3Cs1sMVpU38scVHwyRQ1K30rgjysa6UjVyQdbc7Ok3D+bYv/
wmpPtruNleBjPSuQaztk8HaRcrrzp+2LlIP9yUC7PMp2nZBg0Tyk5ZGxusk1YRC0djetm0MuRSLb
KnTcAuPBP9HWHTV1ME428bj+O7J8HATKvgvVo6lgoN0v1XjylwVtXOg2WFJSPRGBSRB08Yaulsfh
ruiqIlWjaAniZMsFVi7GLFp6GrEGGMPF67MzJc1WiB6STf1plz71AbEK6du9Gas9YK3gtxJfkoAi
CGocyQxsKcMeSYfkPbuXrFez824RoKU6LMSagTBioUNGhOlu5l5uixBEdp/vdXOq05nnCcE+xFfR
PpngAcHLvQS5UzFeJaQCoPG1Nb9HKQVaoi51ci+4GBbuG8dTJLZDlsV8rT1kMs1IeoSWjtjYjp2C
AAnFKOca/4tRUTtu8isNf8tYODIQvwW+XTrkhMgGQyYqRRqAgUCk0nmgt6Axqd8E0BA0J3BTO6+A
smb0tUdzuUu/bbKGOuFpu37hNMZxBTNNMeGsOPvkA3vmTdf4pQyL+lB7V18WxGsfcTBPj5xMgnN8
3hmaSPcEdi0vnoXOhLJKpJoXlJfZwlqNB6uTulW+/ZyiioqTypMAQ8NMEEOQ4WRXH3VIsIdjVmym
P+GtMp/mCtI4WMaOWrWRFKe4mnZonfgIlfb5PjjagBiXtwgv7BzWaX7YXeAgryTLjYH8jUg6+E+O
Vsu8p4ezoE6PIfbMT6Kdw1d/N43a8f3c75nip+qb6MNkCUY7Fuu2S2nV7Zjj/cjyeNot7TX5e2oq
11GM14CAaqKtm+4d9c4JDPzoI2XL2CzW9qL/W6IXgLbPpJB7yQJ0fCNUfnWNjQVSWRWZZu/UghUH
KHecjrf7YjCjxmNGd34e+ucr1JcLYq3JgBsuL2DSasjZ2H5BIOoDkG/9xPoMHm/R2oLdq9QMD21s
C4LHezpMnbYs44DzdTtF/+iEeV6GPLesVAMFItajJb6HseI7h6pC7HXvonWJZhEgbQXVabEWHd5Q
2lRYoZKE93ZsClmt1Wmjw0eZWHvfEiZj6ERVjnc6tSML4MWcQm/TGU1ZNG6edv6v8llTZsCcUssG
LmUhleT6lhj0uV6y08s9w48QENA7xUD8g0wblsgzYehtbzLqhHYfJaMA+OpgafmVItuq+xQ2IM6R
uAx+KBzcpQLM1rjwvXgTrGH8ItsUDbNPTSIOHmRXZQBnrKOkqJRWMstkfZLMUItEcucE1UmSyfgQ
PHjIZroEQ82p5SQ5UBrwOTO4TYvIOSMFkIXL+PUqh/Vi7iNraMYlYuUkSomucQef9EEfpe1Uh2oI
ffHvdo8GlLTi36iO3ROnuR1fY73Muitziehop+y9DJI2B0JsjHHOgjmQ0q7CPEtGK/j0l2oMgv93
hVGEDVlrmvm59egGudAPOeQgAaSsMB1mFdScFdyKuDEM+jRHszHW8tuSQOK3ElPExyTRZuxqvU7f
2wCJ76pXybqEvx9Exp/FsD1hzR5x/vyCsQoP90Tj0YKLR/l6Ha1U9Y/Ax8SKxvJF6KWHlyNRXy9r
Gtp4+WO1D+oC1/4OwT6bu9AONj2fPmxxl1H4AQhGOIXBQwYTlTVUiioNR5twko5qacW4TgxU/6wL
Mft4Vv0ioTYjYrK0+RmnVONaNX7bptvybUi0sZj+Y3tcZa41pWQnhvjjgDTZmhq59svFUmrVZD0P
mPer7zaCQPYkCFPl/brXn2H8iOG3SrcvZjft+4vTWjcz8E+FnF4BNKZ7eCSaY62rmH4Hti2/8qBk
+Hp0u4jtoHAPbGwXbOrAjE42xRhZrd/WyHAa5JPbuuKXnNu+b4IEE2PhRgCaZd3wYazRODMPWVHs
4omraKuPDhu9QpCFHMldM0ObkKjenVBt7+yLqxZZdmEdooCFtSQsFCcDlJfF2JNI/BKIUiu5MRDc
oAE8a7cegizqEAH1kVwzkl9aoVyi7EsWOpZn6aWbi2ana6rQ+DbeOslSbngPAyR6L+GEmVe0MTb6
ajW5l+C9UVhTxA8i2uEVvMxbyMAwGNELY+gwkwvfOcunyFdbGk7T/y0JOaHfh/m5ExswZph2NQKm
nWDr3VS3yG7GR/P2dF3Dc2UpTxEOwtEZ0MbDb9EyaT/0HdANxfqsJKPG12uCEcHkDJVJe+fCofzk
E1W1/fPt5/1EDZpupPrnGbAJatPSzI5eqcMrfZNcTjFtICRaihVly171x72lJcTFxw7f/dyLXbEf
CQEeAGPhS/yAuc/jmiohmqEWAoguWDh9CdCBoo3GU0lUZSkLrJP5SYPNGKveDM0EN8szYvFj950w
vAs4izxIgfyR7DZamrXYaNFODnQuAMvg7NKWrxZULcwCFrE9YSaMFeRKIwNMUZ+rF1PglMwSSv2z
CGiW++a11ux4f+dRejxH68woCj7gVxDdxB4iUuNyZ3R1WAhBM6GM7IrKekjlgjIYsjqOhoCE/pJX
PUySeTeA8nzx3s1gxkPLG0bZ1EqVwci3dxmkmp95ZsvIMWjK9uDEg/7WXsO+0x0mTOrBugA6myZu
LmLoc6mqirCz4bAOTehdfaO2wblVO0ZFx+fRoqiiqPu3+bGbpZT47VJjgA74lhR4PlmMm4qAm4rC
pLe0PnFIGyaUiJLxdOh/JwMDSnEYns5Y7Dyc1VJbu3APGyyQIcKOiJBWwnAj4BBPlip9Vuk9Mf9U
GBHOjAVRmL362+gB94DPlusXMBPBSd1XSHuIUb873YPM8F1VxAPuAvdwEuudiP1AGzZY4oTf4FUQ
hkOZ4GYrdwWI6TjOeqn+1MYesNBQ7GyCkSRJuC4gdor4MQVjgxk4ksv3ZvwuFYhBjbXFv4H5VrKR
SFb4M5BCNxM3SWIaA0Y7BrG5T47IZu23CLEn+4qRMIz9sfnz/+PezAfBLHtKxWURSRkKJoqYSYNI
dH2+6VyCX29qVOeCIwc+ZnNiWsZ6mfBNb44kwFRSHHyA2uR9LAQG69IT/H0d2aYgB/yZF+dFjdDr
YvZ3tFmLAnreWqvrgRnJY947TbNFQZG+YaS1bWsnv9iGa4cd99MUGKL3km9gci7HnVJDRYaVMXsU
K1mOL1JmCZuFOUHndxOavPxN8akx7YVhGqRg4d207q5aEhpMRZoXhKWQJzdJjL2VajpYYFulSfMb
cTD7SiKzOQq+38+p1XOv79/2ssdeh3MM02WUBYc4mI/joQXgkr5PqB7u7Oi4P0XguSzJX/iK0PCJ
2usl/YgGm4MTgJNjj3xQqh6KbAVTR1EtRVl4c6f/gEgjaRsee4VM6UoqXtZdd9Q/s+TxAtVQ6rv9
lyvtmdy1KmTf5/Iq2OnnxhNMX+fzMnqgAg4fhvzs0lo2jvPzx40MbhqM5H+vLEyEcMGT6lk+ky4V
F44cTxe2YnVT15jig+kFz05pLzNVWkLxbVPmJTsoSEkG+TioktF+A7CJFrOKAf4z2Os7jsy0nL9p
G/WZf4GVc2HcHJhWCIz8GICIfxxU+M8xBfZLkWC2tfdLfbPqvU7l5lhqGGOlnrOoDBwIlHDamiGU
SV+dEACOMxwo/BvQxmUVsI8ngUTEfjVyPcUDzJpssEFfLPsPjLEK9wX6EgXvU5otgyuJl/DC92Ns
/f+xc1Eti1MJBja+UxK+wMrP42tZ9pNjoASiicZQpQp4v+IDGFhfYmYSKCW2m0Ec/NFajiJ9Flva
Lz5TX+55lDtD8FgGg+IaCozv69Gwd4YJUBfrgQTi4umNikDyplJmXIuNt2SBcAxMDOGD3QwHB/D+
QC/MDzCTx/KOl722boMO1DiBZavaWcYJWui7BtEota9C5pxafeE2BD+fcsumBqarxQWgpnF+Du+R
BSFA5Pvd4Ki+RLAskN6gC2PxCfotZATrf9JuyvnX3mrlfRk18VxhKgTStB3m9XmKAeEPGm/72QLv
KKbe3DJuS5a4BL7jVD23EnmZzwl/QgauEo42lueOiseUVAwvLLM5AQLTtou85Vqc3gPH54v61lmP
SEefbYBd3NlqD1vzlyGYoiyRV+2K1q8Y9g++z9M9aIgfKZXR/rL2sUzuM6wLUPozcC/VmfFkdxmc
ddLOpsoqOZSEsO9G6pHW04gmDuYYiSMiorMbgpiYh/7myEa/zAAhmLrS5fUiJpWClilk6/SaOo9M
SrOFjKujHRJRNg4OpjHzXHwvgt8nFlt6h0hH4p+nHHa49OWF/aH7LNSrtkesG4faP/rJiOuy+9zH
pOFDsxQ520VcbwdFbUwG8ZPEzKCPj+w3Bz+WOM9qMKNiHscW8kiX61CJDjJsb9e5h2pdoiblCBuc
cMzoI5euK8SLw8Vzd4IqNvtR5qhVftx+v4PsYnZXJ0WfHbbyz5RIdhg4mO8R+Yfh0wpoKCpFO7Mh
0T+VBHpZIl63ffgCS4r90wSW3zfTiVj4/8jKBbFrjJo551mD1cksZKtwwxOL9d+M1z7iQPeE9aKi
PubNDdsOambrpjsd939FcKTl8I/3Xz9ACfKoEnXtXDd5AqoYNJUuCHR7zA6tmH1TmvsYqkG7MY+0
DmjTkvb+Fw3yT9et74/l+BKoMMKlnWR0e4eC7dLpnYoHzEAqOAdlWhycgv9SQ+Z1E4/I1u+UbUBR
vzlJ4mX96tU+jGrT8/2vywdYHUvmcbEKOzjdazhLaBtDB+l6XoOE6clz4av2bpVgl28KDN3fQp7d
Q35EwS/JKXoYFK7Wd6hLGPLCKyTFCgY9KRmsCpWcHlI2UamLWkl5RbWnRhTXi7tX7t92IWeP0K53
C0HGadGVQnyJjo5N/yD6HHbdp4iJYYIKjjhXv7+smtjCyjjuwXBwwSjlnRFhD15u0w2XtbhCBvHR
EfcQhBJtNZd1qYHlXCBy2c2otYHG9I2+8eG5Qo54gdk3CStq0jm/2yZOuoxa8Cx6x9XH7VEyEJ9w
vayJi8iynep+7Sh1ZM1l4bh70spDezgFJHSu9f+KsAxfbn35KpUtEsM1x49mSIpz3/TraTGd1R9f
Jn2nYUkRcmqrEBYX7Q6AhBH8DaqH1a5V7M7OdBmRv6sBdg7ds9advRRZUKuiSq/ACsPlQ+diBJAj
iFhfiP4ZHOQIqku4FudLFNSLzCN7vOFjTUFAvv153dnRo0cYS7YmygEQIPdOcCkwuXAapkkO+k78
uMTIRltzjaoE5xaBfgdGP5W1zW6chWm/5A1Nat4/ylMyAzUO35mENMk0n+aX3nWQzNrDOJUmztG2
bruIpvO3Slg/N8mRxlB5ONdm7f8Dv/QmsKIus1KoJNNDdEcWs3JMAlAaxTCKUvR+JinutJ/DOXOd
+wM6X34axD6+/BoSW+aPDf+Vkzm2CsIGwDXFvnxtd37g4GJRTl9B7E2oGHzzsQB8HOUuGObAaQn/
Al1VB3GKLKUyDnXrgg8hGifnpq3me19KpePdWxv/xgc1mhFzZubuMVDGg3LMKYGJrTns9LK9Cpt+
+mKTLBvqTCYvj7lGYphnYOAeMSV4EhbhXn1kjWShu/L01l7J/+tSJNxs5332xHvcDD43QUQOY3eb
vUm0/5PbYsujKRv80nmoJPVwAV/p/kQ1poGUcMOcDCVON7yNEwEtMaDxFvc2Pi7NBiuC0S8TH9ey
Gm5N6rz3HUSEy/19deXuRASzj0OGnB30VflPQk4HS5n9Pm+cjmb/OVAbUt31FZRCF8IhXnGDUuwW
E26UDgNcgIURajK/lIrirDkMgU3dKwVx+CMue44x2+qoVEj0ARuaqtWPRdvJzvYjZ/Rs8Oz8oLQq
NYI1YZDHBdHdIIRtNsL1vI/7fciqj+lslsHcWf39CGsUOBY4EP+I8GS7CpFLpyu4y5iQgWou8PT2
eYQz/yx4M2uDS0vtp2JTLFRPeGHgFxj0SZM6uwH3lrv10Oy5vpys3hVOWuMy5JiX+Np5fP/IeTcf
CO7V/SEahEUDdonW4cAf0kARFDvVFV9hblzk31/eF/W8DvfoHR/c2Nep/P3hxlXZLhfRX3T4QHVD
4e35EGIZrvtVYVRosRsaRBPKY4K+cSdbIDt2aUDRUyyC/ywbcTt0smRgssHRpw9kEqqQaHb0Dhik
WVWz8PoO9HCC+U0hZtUwWGuCIKHjYlfRgMedpow8j53lDmuhxCSQjmb6lmgS8YOub3SQ209TqxSP
dWx/mMDnbsLW7t5uAmLoGEXntuZWTotgJW+Tk5ZjxVSp2xhmbb8wwuWaYhOzCTZYcCXdoN7B5JbU
9a+I6AXIoirILe51xFx1uMxN+Qe7uT+e6f/bRB1TGbXlTreXCAEkyH15PXux15+mQ/rsA4vXaVq4
VncbUomjQkV7hnfaoVaNli/kJdJf7o/g8odpEN+a7lrJrsn5qasn0ovt+gy9Wmk7xneJnBmT5kGi
zq8s+kbcc08pS2MhkjpW8S1Jb77rFeXlQ0Ai+w2Pc8WkuMuFGIKSWHGLIPJZKxzZVYekGeL7l4at
hkuGyhLin7nB6FKFxvITvqyBeK8dmKWgfNeoJY7qLYN+kF7qw7SWuRracEZYB/QkKy/gdaSXffMg
CNr53EAXfxFQ6X0ObodNFYJuNVk3hjXETE+AXAnoXPwdc3xxLNsNLT6WWURQ2lg3gH8+1IskzDc0
OD6esEeLO/Xd8+SMHtJP8C+0paKTOJnVu+K2QjvMrGz4ugzjZMdOYnIqPplfmuQzrmTB0mXvOLcA
AaS6g/ixAGXbDytjYkenBoCBY34LKvlCKtrrxEWLuNAmis6zn9ni8JJ7B/LxQcgmRsIWSXzPljqJ
XEiY4AmpsOaCH1z6jWBAZFbOFSX/aHkc73GxCasF+Cn9YIa7nDc5kemDw7gJkfZ07JPruP818Hkf
4hhtqlC4JPfts/UDAqSpErrmUP+yKnfc8YZzs9JCRzbln7lknjBvF1cd4tInu/Vv0d2ciBR/H22A
1+IcSWjYfhfoWwFYrXlmNLrQRMSGTbYYljQC/tsD90MaiIgQFCqikjlORuHI75mT/Zhc/1VVX4ll
DdbhAs+5nOl3j+65ybFjAfojbPO8PYKvZqEDstW7ObrRXBWuLVDBMEKcHAgpmZskzNGh95eORues
KFC0qlekRXBrt//f9/7OQL2shMHTHUCJRB7gFOZPI+oJ5zrnLEgSMgb2kbCxGdI7NwAas1Tyu/wh
dQr0aQhjsvOcIqpxwlcjWalIA2olhsmsVM+0sMjEF2sz76Bv8EY/iYn8TFRslpkDFdUnvejok6MW
d8Oov5Mz4acxvWsnTZGL8bS9nEDIDkrrJJPdbXpXDlrhwlc7hk2uuMTdmnC2cO5igS2jI4Bh7dAz
GIcQhtc/ktNyO3KEb6P+8j51TCjou335c1ScLSclqicNM/SpzrNoVa8nXN95dtFwXdtF1aF1wlDN
HaudMjVzmOO7Zfj54E+tvT8Uj3CfPHEcYhfEXLB+KyhImKifw646Qyn5KCkbnKQDa3A7sIGTV7y4
XmhsoIpTi5I3QuG3SIHVd95db3Km3GBCieXtwjlL2St4P/0ri6e/QUJImBwWxGud9ZpZWsPoDsr5
/9BU/z2NuGiRTAf1dv6l1DmoaMYWiiJ+Et90TpdHhvfrYmq8E5Oodo1FzSlStICEhO80o+RU4sFf
h7Xu94HzbpDOstzUyWWuE5cUAyzo1WOYLyFKxX+rzXkUjVtrxjcOOaDNwhu/jx/ypRj65wL1OPMP
4I80fgeKafPDJvwaMcon/53/Wqct0l4Sv3jsU2/Se/dJ8vBQRAPk0bR+Jxu8qr7TSAxQxu4dEQYz
xfuYJvStWPmwviMLVNvoQDVDjyzjfR3Pfa+71PU6NgpLyPXmmYOy3/nMF6GtYGuJ6+jhaeZC1j5N
z4Dxd0zpTmAZGUeUwjBPpSIQusl3DZmboYLJvMSAwwpmQbC+4eccuB7g0kMEKdUq8sdUIs9/lNdk
YhaObk8Ra7Fdrgj+3UZq7g7bJgR0cxSXyucOqBFn4KD/EzCRDoOTgxbzn1NTwHAP2F06v2h5IzkW
143TPYlqjlTIQ7mrkv+JwZLsQ2gyhHZurmz2mRfKX1lVDrHiOfpTYPPgpNO9zpL05rCRXx3ZzPCL
mR4psYniEv0tRk2kwScpml3VvL0fFx3bJzm3RdBuvNQquxUCVCR4QNjb+uRzIDfy99tQ8F07tILE
Bb92CKFE8BMg5oLo8gTOQ+sg0c/1YkmMR/FlRODGi1MQi0tYDOqtNBfQiCf44QruZdrF+k7+oQyQ
dBsDpi8waKR2AlPpXUh15pDg0iFG2+ZpX3e++mPFCUOFNSHHvcZPLno3J4BaJG53kAZcSMxAMtmW
y9JCEB+uMzKaSWzhMJO2wsAIgZxXH5q4vI9e2YJ/+lSFyhi74CJIUeac69mpO2C11ByfztYHIz3e
dTzYRfeUn1jD67C7+TfW5AGX3+915GZ0tmOaDZ+GTkIbNDy7y6VsBba1iXz3nAlRgWoqElxWyY9q
z6QleMXXdkvj7aLqX9kJUFiYPrm8zpYTyDy3/Umt9/W18IWEFwQDt2oTr15cMrLdY5YCQiv53mze
NNhsgNOd/OLRAT2/7cTg+TcJuCnp1B9Psuc1qXUXJuNwcQBkI0K4GUzUnoa7PgVIhlKAwFgKbnIR
ejKbcVQiKslQAaEMLbruzB5JfsnHUf0vixoZ6RJv9SZoVMk0WcaNfmuWiOt/PWUTk0MR/HASYaFg
u+oyyjUBmrg8AY4ifpAQTlEfMFSN9/3xjri9vQYbPFKoUAfpUEIVxGa85V+rkaIlG9mbp/RdQ++H
cE11GqgMADDSB1VcV1hcpT34+fKcXbJGI9O/fTwS7f2z94LCNT9nZOvCiX6waQLDPvDnz5hXRTNm
EMxm/2Oc3OIvX9E7xh1b3I3VPXKhwmA/Xn8VbjjEg0CaevQRwBYRXt0zhBVYVYA9MW3hnUCaZ8sk
jpOYZj9LUY4pFW34p+TgBSxPCmOLcdQcIEEqkuP+NoCTYysZIWszSKK0NLzY9Iukqpo4GiUPU4xJ
3A1S9ghDVumrvKqJNbfy1SSgUOtT6uGSWeHJvvUP/wxwZEDGrD9JFugYhrih/di0/DljkalZgL5Q
dBmqpg/Z07gBREat37HY19vGxcTKA4sOk4vUGYbkatPJIN8HRiKZQj9FAtd058jsAxEbY+yKvtd8
mp/Ww2Y5fNJcXgs4Ve5yyq5lmCg63Hnet5UXa7JFsQ8rG3oyjc8G8rpaOOpfE/N50dn9GxYMqe7z
V6YaVC2Dy/Mj94IshCc/CYA7Gizc2Wmlp50gcace/K52BILtqHxYIRKi9VaAEGkszl3L1HfCD97X
qUpcDfExtIl1P6cARe+gTn0wKXyspXsVcIJP211vtdIYJd+X/yQYU3hsdhekkAlVmBO29WkDq4Ds
toAVDxFWqLanSxxnW7oXw1wFlK4uYQnKK1N5Ix0AzP4HBHwisSpQi0qJPc0wv9FIk26VfUvGTFqm
X6TaqgBGM3lz3WmcF6Vz9A87PEKJ2uCrbRj5OpAmHVvrdwqqCdHE1CeGpsIWB3YEbsNrfkeiQVQJ
MKFlPzG74h9rPiQVBljiyF71tkdepYc5Hy6VwTgQHIskdvISMv692xoeE7HuPutRgxTS/tT/zHkX
Apq+K7F1aV+PVGd0U/mGdnUCmKO9TiqySB7GrjleRuDg0XagGeBSAt07B+kCU6cDWTwSVDDSvKmk
f3agAeO3QiwFoSdTiCul6s+jxaE/sTlHH8CTYAm7Fi977ul9K1n4fOo81H1K8zDtmDzRwbedy1vw
FXBw4JoSj752PrHYiEGsLwaBnYj4UooHmBZTLSK3qXv9adufKKrEmhv2vPnpJm7GVItGktKCBWGh
nT6+9a7U9EXsfTt2qApA3Wl9zkT8b7zruI84DU5LADyoFJge51WoP45JAGWDvLMH7ocWwcOOJnr2
SAjFwqugLWNq4BvzjMzY5WzaobMThETZJyQByedbHAqfePqIcjLOKvW62JU3T6vzALZ0ZQ8VjpEZ
cmHVmH3kGVUnZ2q85rwTSr5gp68MVGORW8zipoYfelg42b7gQ/xpWHO9BfN1f2R9AyB0ObPEDIeJ
sDXOeitbkXzv3Kc9SwaIfYv70AklnrsmhonUlTHmRV7fBxrAALDMR3DR93j9Tv5jd0kvMZ5jCmeC
DcOB9R21iqcipp5xoaQOeblJKBtSXejDBuFAZzBi+RU47veF3qMw3HdhNW/bq6IetMGBj0zR3H+r
CarqX3nAXBIR2LexMXJNd68lIL4i41jc5KGex4zbzRBvKwezwSi9bWcAWZdXkHAOoUKqYqpOOSQm
M3s2BcdW/0xaFUSMCyNamXM3V9yty3Ji877KyVuMzrf4dNZyO9rsmoCg+x7i7QJxyGnWKW34RNrT
qlz3a/lQGCJl3zS32Cm83+tPvh2xijBjYfFp9JwpFl/fYqVEBebnzq9SJHDZ4Uo6EqtGN20/ebUP
2RCVWicjvvAtbPM+3+l+1d4ZK2q5pNenILcb1Eofos8o1KHtZswVfimIJcnaH1ux94mj6mdH/49Y
rhUTimDYHfDiM9BSz6QXVeoW+zmF9XXPXk6bVCNpD9T7Lq/YT0kLXLDsH/M0zUiyFEqWBeDCNtCh
iBq2U1Or5q4Qw1hbZIa7WM+wQA8z7tqDcyoqNWtdxIn+8SjJg8EiGKpQh0VXRXs8BrWz9j7Z7ldO
2P+K5PgHATBqnsRONFQ4mwRsloruBXdxtKFb2UdpGm5Oe/aRN+3TCsEcT7CW0MsRZHq4p3RLk8bi
3oJFhC9MtrOB7SGf8dUwLuXwxyEtt7D1Z1UuT1Ew1voWw2Zm/jHmmr0cBZ7HX7yzzbK80W4NvtAx
B2rzRqdGnH7mFrpprRQBWMGhaTQ5NltahMauCrV0L+zqZKVdDaOdwSOdVzprpPLP5mVxZ5wZ9iSG
C4gAAsOZeuvjtNj0kMU8Eg8ebVIN4HmQZcYMZhqaRkGqN8J34VYlR+GO2A2kR+RN5YW81UluKuV6
KAPxBDvMprcVcbZ03uoCCAFpTp9g7+TWmHUtNpZ5LhgULEXhpLxaPlsbnTyYKyiYxt9P+MXfJ4wz
P0WZpFGXP6FMsJFXvtGNkoXWk7aznEZWfWzTzGjwbNQ3NZmL+g/8nXCL27XGWgI1j+EqgdTCrLqk
XK55u0uFMDN12VJcA22quWZbzMWiGRSrJfejtAzo8moGuSOrk6GW29tLcWl0JeLS9jMgsEark1Yj
mFFakZhMefN1j6ykACCUlkyahWDHFvzp8J+uiGyME0vnbPYPY1R22MxeCYErv7YqB/O3SHPfgNnB
lfUJI8GtEsXJJe0L9NU8govEhjUTercErx8NouJAOrn5noqQxUCuKB0baRVGPWxxpY98t78DEwuf
pGM7enViRRN1LDSc4WWtrWGRvO32yX5R/sF8MHr4YpSdZSF9ripi9ih7e5pWngaLtTnXfZs6xlbV
V4nftN0rbfQmKKWfEjH1a5VYAJsaXIvDT2vjKFGoU6eYq+FJJNwau+t9N6KjDItO1OkxyLCXtHSf
+dapAHoxsUh3peYtWCiIFiZw8KIEFgL7Pmfz6jcHagyPkgcLG+M85Vsf9L2ilid8d61SimHanRRs
zVMsxLXVqpDCtK3V+LtplGL3Tyss+VzHOl2MKJg6FbOAwtciAROOzFFhCxZd53vk1qe7Wrn9M76n
A62LWD1lCBSi1BpV/jIX+udEM8StjCPQu1wIoibwbbIYNNYxmrOlF8Q/V3Ix5pMT36GMPAFjdlKY
8LG7sWhA5r357gvvDAEeW1697sl2rlTAo6n7XjHX3GTfIAT1lr2gHUkJHUY1EmoPVJb1mbDfJs4k
dd+z/z9Uvyy2QEUz2DL8stwBSCNv0b5FngGtjaiZeSfWFDFbQYOZxeYHjQYz08sLVx3+lNfoiZFO
inr2WSvN1CE/EJ2HHmjqDb6Lc9n4Co9/XKr3alL6+x6Qx7v8XuIkHFN6X3x6jZloTm9BP06x4Ucf
eSolOqU9soCY2Uic4ymOb947Ofc5mJtRDWjiAmAY6Okj1UVW1Wd/qeuV1hDb1zpef8PfNUgo2LIf
lkvU2Yt/R8AllvYsZDjPsLIf0o2ZAGywH8w56r6HkuP/hXap0nwH8DhRCWlrMvGPhH4KqVsbDy1X
pPjNmJuOoJ+zTdlAToJBOky3+4N+5E/EbKWZ/l31JPKZvIEoVV/XLDFXno4HztDOH/HPjm6B9NjN
OFA7G8j5dGnNL2NPoWVe93WCyg/oR47LI8ihGmOtgbKlXOISUst2srixL+F1Qr6hC5Dr8O+lIQ29
mNbxoHcVf8qf/N2BMGK5JeggHqLD3iAwpjUlI8uToCjX2q9ve8eZAjPVwR+MyiRemN2JUNe4xEtu
Z0NieHj+wP4AQ4TYVQ9Lvxft/OFdHzjoQF+49EAiPinfkeD9mRCpXwh82EJdHPyAQJBlR7QLtJRQ
fTYqY+WjAIoiycFYqIRkM49bsk//hY1zMhUmluch//7W3UTx5kHip/Ir+gSQ61rQ7PNcZBtm8e4H
YVUrK96woQ6yAt0nd1/WcyJqMDLds+1EJApr52SvtnkvkzmoDIzi2R6ktN6NbH91uShFMEXUZBvb
W6k1SjkSc8rw0Lt87BryhrW7Nw8eWTs0N01dC0/tFCcNA/tTVuTWnaBB/DYckFgidtSEB5sgweV+
fEzWNkqdQcuvByaWl7HIfuPPIaBlAyF7e5qcyl9miZMgOiaMPosmvLNR3Z4dn3h1PFrtkaQuAcDh
nPv6nGWauQPRlg7+pIyQyMz/ON97E6VcF8ANQsZrdM6c0lyZRvJyC4+uDqR3Y0piwkMWQWmW8ZLW
y4Ox0zwSTh5EPatwoxY9RiaaCpcEhWr3IsEKlhUL6/bMftYcDwEAnwdWschu/vV7lVX1PmjFfIZ8
WRyLaj62VyEEVD1wlwNQv2Rbxt2kBER2U51WU0t5FPoG0IBTrdGM/L637WEOZo/TNDRrScBjQS3+
hmYsSPip7Wp8zKbwjVg5j39OFRo29ne3rTIGBKNtKyeW6ImHL+9QPUf0qG5azv8gyrpfr8QSve2K
KR9rNIRHYcSsVNv9h2/w3lkJqK0fEAbt52bFUcnVcR3HguH1HL2TtOWCrUrAMWxRDPuAJohxzadi
AqubjwFD2U2P7WtQm4iKEeubolOgHTBlD9u2ZzlQ8tq+qJk8gzPHn5y8dyjSeV1wixmlXWrk5bGx
Dh+pkWAB/A5YKgCIpzg9XyM/gKpLywhp4h4q7yO63DaaDDNvK8q1iBOvIn9QfHa/EzaYyXEIUo2e
d/Da2/BMl7QA4ELVAjRHtYPEzFZ6FC8AzwfoTBDzVNn1LYbJjUwQCtGDHl1ziSw7mnSI24f9ygl5
KfKRlxCCLRyZfVUhdcsviBO01fKk3RwNAgvreCxMHvkC9y1YTpdJVoAOaLpZanFGSSdujmClIEUn
u35njsSa2TMy64GBdCGyYykYHFD4nPbAY7uyIP81LAZ+wgGh3EKtEPxFyAvL4Ks1oeUvh5CD+eax
FIJLBPJ6Jb4PWz5wDERsK/wXftZ98bGA7zfoL2nuhvCfsJ93Nv1sAaCfivREOYh80h0cbwoIMAq9
doplEkRZoiMHm/WFe6H3y3k3TJtc6UWwH/jZ39mDKUKlJ0ITXxqy6Os1jCr1mAvfr+FWHr1nE2Fp
ukWzm9bhJyHCYO9OyRitS99ZZH5QZuIrETaP8j1YlOqhx7BbUKglruP/iEnX4RFTed8bc+C/RwzZ
IDOQXFLJMgiMBAw3bvZdgIZY34JYVVWyr7xp+FiBlVK9yCDwp6rY/Qh1Gnv78IvkBbcSd6RxxHmj
tEAhvh9cIYkHF3ubRf1KydcGmZdoqGEwvdgqA8549mDy16UhX1yMlmkzCejpFrZyM9nGxBdejigf
KwzFEER/nM6HSPK+BipTF7HtpoiqOomw4dGa4mbl8wRk0Lu5a6PrfDkgz5mOa9egmlzOYg1PMu8b
WM1X0gBlXfkS4ksy2PM9sDxs6+Rko8mN13NBK7ihNUNykSJKrsvDFXZ242t+bdT1PNk5JX/eF4Eu
ltUoiFEtejwBNkQg2+3GRnD4UOh5OHtXX5Jj6EdP1kmovpbSKIRQhy+YDJMkuO2mwVIRLMBJl7AW
zrM+fPMEGE1/UOsycnR6ywxr9dJYmOCY7T5guqiHycTB97lnTvL+OKJDN4cwuDNE9xmJJOlEzaDy
92iY24ivr0OPn0svwNthCgoeWeoXY1aiiwqJlmiQNkw3RERjnvdFoq3yOwIsLg9cBaPkqYv96JLP
pNTkwZ19IuKavhztUZ0El7aNBwYIQAbuRRyN/cCDbj1iq5EAXRH6lZp+7Rl+ngqCCdZLdCv5cAbj
/0e2ZZRag7S21airLpvvXjpmGHgngXA2nekiA6PVMmc0H7ISEB/ZIOEIUipD29LKCcXXHh0WKx/k
8e7UF7y72An/wO3WAZ6XphEuAYN9iP3app2xYUfwP1GxY7z+JSxjrGSW+K5OZx5PLL7pFCxuN0Tz
Q3Ev0E0M08qURiSpIFXG2MwbbcsFyrFbQDkBx/WS49KxF33w82URKeg8KcWA4GxJWVlE6pC607H7
z0PfqipNpoM1pWTP02ZK/Sl8DG0R19mqeWT+MiKdqTE5JQcF7dk5SI5U1wPCTDVSZM+ii9BbS5i7
z7mq9Liqm+XFkI//2SxbYqrNlDz2MAKRqukjsCGwPLyN836wgxPq6eqeaezStIeQFcEY8iaIPQ0d
UIewNNxlXleSc5OADMXvJ4614QGvKVHjHkuUBboojUGL9UGjOCqReL4P6fPBn1A4RJEUsoDgZPEk
85/Gdx4ZrlRGWJK+g18VzYbsKK8ew8fSfgAx7eKLun6FL/6dtNvnE72c4KIXHxYDmPwalDoE0yit
XiRUDzsS4Jm5q0PM6PUO4fer8hK7igRVxSwrEBtATKPdHvvCcYqN5JP/jKOV8rxBgpDCpuOJGVSc
VFUqql9BZZQi22R7HL+atzfbTxhvUc/GnPko7xXmPwvnbORra92Hg0+IADTAPeGWEDEWsn6d3TMr
9LbfqfjNUlqWcWyEeH/OssmsFafRWzV8iJHGo8AQwCZBO3MO/iDumhQ2RDjNMUBIzEwsiyT1rFyR
H9EgfQrJ+YobsHFb9erAuGgP6d5kFQU5x3uEVoxpwBM2EQ0eTInry68h3NN/9lExMG3liy7cqKiM
FwQKY3+6ZHrHvp/zQ9F6fA44s4YvStsylYZSKJD9+ifx98LPqTEtX6Zl1tzlTyhyGbU1vbRhYkNJ
SAlCKeDLVZ26k8L4F0UmHBUOe/Cp2wNljtZcL5IN2lAiRr40K2e+fK3ZJDcFiJY72tWH1+FxHN7H
UVGohJ1soOU15E1kPB9eGNGfrTSCUOutnCDJA4X1cojyigAfeQpSBGILPvOCcVewpoSsaK45nECK
9mC/etP+CESQW7gYIKV7e7XrrCklgdVkFL658qkw3yDuYFgIHXRlsTIslfbWzlAf+uvkecyVjOyo
6+8+8O8B5XfwkTZP5khtSL1E6erM7eduXP9qwzZCeD8ox4vagtK9y1m1baIgTVE9oXH58XRPjm+7
1qw1Ot5ZWf38PoJXPkunY64UX/oCEmXdudBvF8jiZjP1Vabf0Rm3s23/mOnMR5QUIPfEPiuMLH/1
16thaw99DynBB8sBkixdxlG41TvZoVqBHlPimVafIjg9vTW2Vme+n0YsLHGwVkBRn74bkyv+lZqj
+DYfhsKfIOg8+veOr5jj0vIPAF+tZUnAul+ac1DxOIok6YPMfxE50A+cWseOcOhonrrpWtnU3Ake
j7Upy8JoJdQok6G/N1uU40R9pPFSMwKB+uwt7cbvXinM/PHJetF7H4IvJQdy/LsOkhrIxYUsTBA1
m9llw7lK+2BqhzPzdl76BYcR1E66ukGMR2VIxxyNh7Qalo4xu9LdknA8P9VrRuIZvHNkBdF7fuWA
tRhFRMn5F4ZvCcnZKW/SJETEv6o6Gs7OG8X+S6H0GSfU5D5EPLwlnuojEHVlSbs9OqT4XVoEMFLY
M7jx2pX+1UrchbB/RgTONbUTIHCKoOZODKbKXgFZEhZ9UzwPctb+BR0jO96MCvM1IRNSjR7mYM5t
LyEyMgvikvWGxmO+47p5zB1bo4NdnuoRv0RhWjtdxyiBCvxMMjvbSnABdq+ZNPD5q/z4DxVjq4pr
Ss4KAH49YIUXx085I796EczwwDB9xjQMkakKkRoHwod/u96M3nNAPjRe28E5nFmT1fJ/ikTqas+W
5Fin4H/dODYN+84TAi0//lQ9iapLll7yNi5jGNZC664R/brdFNKmnK4IdjlJ4bTZU0UgWQ5Am/SM
AMpGpO3modVpI6omyrhR/23AR/QK6unJnE+BpF2fHa2KpdOMupU7G4fIZjS5WzBukqXiA5XhPa3/
41NeOhP+tb/nD/bZWb7nc0CwimO8pIQ3pkNBz6ORlfBVwhpJQDrrFm4ey94jVduSitslSiiocREm
FdIfiz7wDc/maRe8VHX2p/GzSrKvoPf6FJahfsUhC1uVPwbga6Z4wMWjxbJYpXHbXEq2CS+echbZ
bQ6SEaVpCheb1Z/nAmg7tc6sTLuR0TDXxkxuZYImxGb2Fo/VMlnBf3c1ofodTwV2BU6FiblZELzQ
Fi90zntplYtNBSceJiu4Ubm2+lohy91k8sqU56Ta0USPkXeVrrzRffUvCZgVSwHbSjyUsQUKuCWr
asp4GwNpfzZZspwTmZcs80Q8Yh+VnjxOwLGU+Jh10wAqo1cLJz2sW38osEbNFTb0BKXc0SInWE6i
jwJkkjcDSnxn5JL50JocOQtnFwlYaRYA+DtEu4U3hs01tgwIjHbY1nMDRKiqboJD83Lw6wjXV+zz
OPnLQa6LllfyTUd00bF1iq5aDLuFR7LOQeULoOxkJOcp3HY5TnO28cvef8zS2tfBQIHhV/8PccZD
HsgA+I0hQyoS9TRxd42JhCDxyoycMaEO8B8h2J0uQcfA5K67j+yF39g81Gl7kZdMwqh2BMrEGIo9
HojAkKHyN6neWGWffzvWlrcN0mKi0lwUURaj5IJfHRG3y4+JRmcctbl/dN9brDucMfvtfmBbh7EC
Bq9DxZ0idrjkuAH03U7P5MTmO8tfMHyi+gRd6GfVgDGclBTp5nNLi6e3KFPxAidLm4X+1RX0jHNf
mrb/v/9xJYgITOoRtQbeGXdWZbuJMxbbGZL1mHsE/tz9DsIje4Qq/7QI/J/W+lPPk4VZsJhYhdXg
Mwg9ErZ/mmGpSmDCuxbzwY4nwPdH1sz+1iGMW5Uq9slVnYC0W8L/puRTgRMwqTFWpA+rZCVnD4D+
SJ8dRrj2L8D7X+eo+q4/GHg7ZY7lLpHt7ukcXU6t7X2tZpF5n1gUoNRYB6fUqZzBJsnYUjMzVv5P
lwbDiXeCFMd9AqBCe+5aP2S1kDEgVN5h0oozoiXVeJNXTI41exRmJnWp0rLdAeE1/hA/zLpg3p9U
dsZcGZIx5Qm3gFqriweNg5WCywly4HdlDF3UFcr4cSZl8caHwfokfrN9RWKvMchenJlokLaRdtvR
13ayCm2veJKHdocxXQP+5iKonZqVxACyxRzAT+w+pGwJRYbsfC0Q7qFbv93nKWIz9JGpxXS3sVnw
CzQ5/zI6PmO4RZC+keIQVdg3Xb7S2TMUkCvQLVZ+2BvDk3mFW44oirKrzOwqkn0e3Ysj4JrLJdQm
W7TtZripnbHdwEf3WII0AlH0SpVmBUAkIZoEdmQNAZu2bZnjOTx7nKNa8MCp08TRwKADbrkHZkwr
RT9xrngPIxJ+B7TiZgSjs9okXLiWtBR9s1dowDbZ6rPZOsRd0TWgBj0kkFk5ROYEsyMOSF/4Gn7Q
kRVD8aZT8iuCGcPgOzpjJY+8WmvD/4dmdp5GFSosKtXHNAABS3by86OVooh8JwX3GhpfTAJ6Gawe
wnc/w5K7o+mGeZim1ByNy0mhmCFLc8EHVlFtnxAFa4sTFqyhuVftjH4ukaM/nwZpXF1IQJNv5eLv
UmYAO+uAbMNg924ZxIbdqOaAPuhJtUkjYzLe8pE21MmAR0ZuIfsK7D+eRgzRk+SLxa2aE+zICZlU
OhTF474em0HqcY7fkNXIRZ7jiDGLe8cM813Ou5Mvy+pvb3nZ3dU+r7sCFuyI/QmibFikai96JWBo
NzPfxq0/alPiJxVjs0cEDlCkIh7346FE9pfi/WD8OlX8aLCUbXOgYOvxBjQ4tuoWSdJqU3H/bVcM
3llEKCxA9mxwWQHYmk97yVQEP3aB+PwaJN/P1Gkc7xiwyMAXIWIdQS4WP00cx6DuHRwaZ/9hZKsO
QEVtsTR+EQ/264e1iRnEBgV+w0y6UkynDwL5HtEtZLIrXovyjlHeQbVhVdbefVSiNWwd0rkn2Dbf
s9Ul9iTnKBhMVqwy6sJO7YjdClVH90g4ES0ojENqrNiSJwgSFqLAHMzixDewK5aRtHisWil8ogxN
Xa1aEnLGe7U7HVWZGX4QWB6cCpETatz05zsMx5vZpVfM36ePCS7zyFjV/coci8Lmgbs0AuJL7cv7
rwinIvvIVuH05zDoyW9s567orJ3BgHvQn0c/Nxax3i9lnBmw3lJel2EELw+uhdFP4uYWwAuUXP+l
Shn39o6Y2PZaTRqiKXdvm8a+mx+K2ILxS0giGx26+S2J7ZkyYLfZwyMRADPwq8iQBmsZ3Lk1zwn1
GK329dmOZGCTnWu0H5ZAvp7w+TFRy8YQ8HqdKzFZ7LS8xoSimahLul40Y0pj7t5x3kYVygNyc2Q6
oiDLf/NHgVih1hBkHEACASG4PWPeIf0QJANRyk+G6npOMbs4eQ/x1PeRjKAX/F5+z4GpqnD/B3Kz
WRfKo3gD0oSWEeogOTkvPk9mH/UlT6KD3Vti9WHdtmLkC+Ag7UNz+cMV7dSvDO39H2ZoWS4Wk+aa
+Y76rGeSBFucE/8VPryTnRHA8PMPuYignshAu17aQx51JvJJQedAU06m13OqIG3ZfQtDpnZ0ogCH
BNzzYS0vx99i46KswJepQ7uH4vwH3mQwJGq6tBNzESkXlEWi0VwSCGO8xn4c66zqzz50GMoF/RhW
qpn2pA5SZoH8LRxAEPhKbdrr+9Mwhr0D8LfBNjX215vzpVDkqVVBXZvJOh7Q6RJ4fh9sHUXrOHt+
cI8BUJeaN8HYSDwyT3ruSBNnKsoYnwqodZ1MrI1tui7VVctfKaB9BqvpqRiZhvyicq/Mc5VNCzJT
3UxWUh3A5H95+XzT/ZBXDcKcxqBksOdoD9n6aDTa/kCFwzp4ciJ2MFhnxr1fzugdBjcZQuoLOzc1
2/menWU7f6TBOKN3lYf/Rg/3XKMwf+nML46cd4TBYnhdqXzPTjP1don9mrNTHEVsBc+rrEKqa+K/
JB/OnHOw09TnTNcuhukA4Vwb+ij8zileIZ/1EHthrMyG4YUyRDLEpODuJl0gLupxtH2jqAx3+Gv/
F1fxy2BeGQw4IlBjrBDe2dzx2AnqjARTZFe6AzZfhUz63Wb3L9/IFG+XSbuRyvxrHXLiuTtG9738
+lH22rY5RFOxdYaG75QH9dBIXs2BKugXAzLTUWnkp/m98+tCfAs6n6zW4xkTRDEeStr1N/v4vX9H
EC1B7V7HCEfD+KFZpMAMUgBpJ0hdoC4BWhFwWl3aHlELaKpdFu2tCv9AHB6iO/26N+wcDh+UnhkF
uQ74c/qRqfjO2M2tQ/oVwcOFy6ZD7sYWPW3BdhL/df1+vQTJieSY+OUPTQUTFAI8jG9X2bVpbg4x
i3v/jGZbO/EvN7l2CJjjsybVFRZTuBeDS4SRKj5WSKR5VJM7J3tqQQQtlfw79MBVmxhXBEqz+82J
Y4Ndz2+U1rxsu0pGiUp707UivgkUbFwQXFnbs406d+M0vLFpNI5XYh1BY090Uo3Jzv52VkDfLtyp
NNj4ZNucWtkAdEw6qBq3nzGriVoOUd5rPrjQ4jDYeE9iGz505FOPHxmjzQe8Vewhm6gg5R/CCbbM
FUxszJiPXL1p4iO/SzqLDVTyJeX2WogFDHMLQ9PQyCQ4C4TTnzL/FstxKRZnrNpJywNUECaN0ue3
fjCC474qxtByNkaLVg797XSB6caAt5XueddNEIEdjgyLFqON/0ylbiYNXVoScf5G5sCpNIpLZVWl
uoNsBKg3N84PAwtlhdrbOWtabqSDgoc87v132y+El7Bm1iGyjfZUVee+OIa0msmwQZb+70IPRdR/
HxERxz1a0kxOtiBS9tRpATf8rDTsLAey4CufxJ4voFMRPQ4lvV3I4dyAUywPEbJRiGrAMmge3kvd
dnFB5jDnEKWGpSFkKcpyYkHPKmPFb96X8127Xi5PKnXyIm64wjLTFYh4UqohUcaqPWwE+jaXBMV2
QunZaPJuXAOLO1xDVUMxtomiexgphcPFUtfVuHdIcwzIqqKcY4b5482cmUgZObUjmy/1GHJ1yy2O
MxKiYHyx77hoO3Fr7UsNvmqyKLf5jTGyG7ZMFDJ8ig8gCThC3W+BYQ6q403BZ0JKpXMmHnPaAUrh
tg+W/FD46AIa6H1jF88C5auqBJ4W6oVhKwRSSa/bhFVM/KM9QlCpNn8lw7sjZVCfo8Pd2yE1/FLq
FeRMTRSNL0hXuDSH41pMCQaRp6BcPLMq8M3FjHpnT4C6Ed772+n5lSMVLwrbk23+X0Guqt/01WXi
MOMCOdq2NGCxvZi55L+6DGAWyzJa1AL6aqYvCTTE3nS1QrdcfFurSpHsnDEkTJuorHDwCbmDSpXq
5unRfT3LSvOouDZ8smXA4CIRu/IBufEtbTu6HwC+/TkbhlFXdze5f0K3Hpb3740d8bgnQ8G12yJn
M3gp5cNWg27PH+k3fmMr90T6RQtnfhLbQNX15Yh+VcEFago2G2YKhClTDgwIyY26dOJGA/nOxbX8
VtvL44szTBqvQmkzFEi9SwSR7y3ki0cJWcQqtNNZrppG1M75ybkn+DSC58fi9h5nj/1lHDfp7rKu
D22IwuekqQAB+8PhJrGhbYQTiwhNvAJK/a98DIkakTq+t2AeGWEHHBDuricJ5+yPe6iT0cEOLYg3
/9niwzf9EZk7KJV2OdlFD/25KQxIPL58zR1UREBThV5Hp+BtUHc3Q17F/j78fcyIENSlLVnXmp+u
WDSxId1RdB+3F5uTdmbQ4W91RfRRpGMFRnIQx617QIYOa9b0kq7HUAHclaDEJMWIdzBbjyyRCEfl
QKk4cZyRGvIsi5taHrSzPDCEzcmyuzCvasnNbOMVWaR/78++cuXel+CLZPocCKKPBhANapaehk9G
fRwVqfHN+ePZGX5XZjX0Y9Dcrug8oUuRul+0fqh9+5HKkq4muchDWX2BXzqcm48B7QPrmHLpeXsC
/jMX2afrej3ZL5oGV81mqRJNU64LEeCSyaHUKtC8eLKsNVAoqKULbXqL+qFplFk0glTrUPo9MK5N
grtp1iq4OrZyQeuiKZdgcIqsHCTkcmKeUdYrkGc8qnFeujI5PH94dFOjnC+3vCCIS9nQVS7WyFml
4283n8swbkYBrn9wWE7KCp1yolOhi57aWSGL7z4haVzyu3pUVDEfZBNBQzkxSxg5ry9RZs4aYmEA
+AP2yEj5q5ha/m7T9uwlPiA1Mwpq0pcte4UCZ0Svr3jxNaIQ35Gp+tjL2eJmLOLJfQltKlpUfp4b
5oTxgBCrRwYGT2oZV8fwYCoQRHzMRIO9FEWnIc36E0Gghz4yE7JuiPaMZtuTC3F7uRswmZtGnROb
zg26lDAyXJV4GuWwsXIgPpiq66XLNovpVshaSHD1Kly61Qi7KdYbAf5IocE+rpoY75svq9236mwe
zT9re74L6GpRlabT9rq1EsHXqUdpYF/E6AatR4SM9MDRCSLSWRM0sc6gi8ZpnCFNni5AhsF6NZTu
v2Y+cko/HJjgjuCY/sI3LGnw0fxTmb/sT5nlG0snQ4tTOyOM9FcgHKm7+x+v/kvtwhOdNze82vGp
x50I8dNhns9XCf2O4oPtGPOPLTxQhASCga+9A94LH3PCJWUd/VTT7y/Z6HUg3UUPVthyUrMEJxRn
q4Vhd6gxAiN4nAb48dJkQC8evFm9XLlbs5cxKRuSlwRAKd6pDMjzSFKbTgMTkNVHfzzeg2U/u1qc
qsfXfVia1J99bLyKjMIekyZy8YUF+dEduHCKNtOpXWoefko8yDQXRfHt4Rjf2e6lWEHgAGyZVE7t
C1EUVwRdD5CbNXNGyTpoMyyh0IF04z8XkqbAUqZiYylz8v6Y4aWPv6lIkWnJEOqcWAzqTl2Y/Cig
NwwjAayAMbWvYufVjrP8jjjOUOU55u9N5k6/4OH5rUaA/JKtAO7yQLvD1fMMx7GC5dWc2bpk6p36
3+PmogN6a56LheR7DbROOcXxYZN7S+grn3pjYqnV+MgSjmsWIbENIma+X3NDun2QdyU/G870Fl3n
9KM9tDRAbhVZ36IfAcPN2vVLHZ66WZls1LP4aW8HCQSRl31PEJ+gO1k9R6ywbQVRmERUGaoqHhYB
OQQxcGCbiQLi6kiadCSye003m4YEYV6GmjnXKhq0b7xkiobtia3/cQr2czlGQH7etk7kduADuMvv
IogIQE2ttxjafP3MfIzoLTuynjPDyrFd3NP8PyykJy3FA9PAhqMX5skaJ0EbI9z+mwc81X+cA9DP
rDuHX7/vhMU36jwlqNW4NRtZbnRM5jbTPclyB8c1V+gwVqfot8Va3W1m3qM7Y1sVM9/rlfNNT5KS
P9bwuCkadUCYBiRMdSQn25B3OBsb1qF/2xcJR7K1oluHXvuN91TUddVJbMv3GtW/UGcoJzORYhKa
7PMv7vSRLDGJ81+5y8ivIB6ySWUO2zRCQRGHjIsPJRIot/QB71HewSSjYerpJiRJlDz6YPE2o+fc
/ZYRIKACPcoOf8bIqMqk71UDyNiwxNQI9ulfl/681ewMtq8ENSnC5z+PkvrQkRw+xpJulounQl2t
7hELlhKdFIm4iNeODWKeVILFcRXUCV+F+XYuWJWiHc0yEhLK5Sjp3y4av+q6PebEziGXlzyezLVE
f+7ORpAcgYEKfA/VxqxQSlqPeZpQsZ2KQjTGdDfgmXseTYGi2C+mpaBFTnkhzu83NklpPvxKtdJT
WVZNbApOSEtSahki6vDuBZ3BOS93LhRSUtAJ3rnmOa6VQ0hJyaOeLuheOwHGJagGcafZu6Y7/kIO
aYVp504TLJ49Ey5T4P4wzVVqtRk/50KCNsSolloCgAkecXeYeuRoSwR54kX53hU85hlwkn7q38GL
IXB22kasiS2rZdLpdQS4CvegzN+B2McXad33GUOeFllP0OgcS3Uh6HtZju14pK0W2YSuCeEcZetK
hiiBgTdCTY+Nb79/a5U/jh5l4uthjaohnt0oM9kp8q1lb0E9tPd8FAtNwtwjjPPJPfuDcyTrqvLV
CliZeAc+j8Dho6lGMAOpTjmuMvUrPGQdTArqFHfD2Qibh4a8TL39V12C0l7vvohwa+NDesGzJN5g
zK77UfoNX1lvR9zelEepkH+pFHe3WnosBYPDUkEbd0wEyIdk3pZRusod8VdPXsXHPBNqzLckpqh+
0vjF1kWolT1+dQIBVTuCkrUmfdn2Q9J/gQbbDrBNGsk6BxJpCs1lcjA9yDLSJ2FpNCM0+jAmzygu
8EcoHXNmOk1zUrxeN6cYwV2+GAuGip3JpUGcMF89JaU/52UUzXG7OUrEoe5E2RLKwMysAqdzBZHL
O/OUmK5UEc91PnvJKOl/n/uSx0pVFcrixATTaMTsIkkY49b6FzmvkQ5TDhnzALkwjHy0eg+7ctUr
cArdQKM+cZND1na7PBz9wodvpqJ8KgZg+H8DAgF7Ws5hHjqCkw1IONUNpcK0rYfvx7qh4LsgdU0q
mgJxYe3IzMJeQb011zxeXQjpnj/VS9Vjd+leKYjc9xJWROIGjGBKy8HHA/aEQ2iD+kPN2nghhsy5
ooyAT1zAJB22fcbgiGRxlGxH8PqBTONAQayc7JRzAcBbj3vd1PbctjqwQ5/HZWaw7KBRhc/wMdmQ
bkLZBw7jDfOec+XpsOKY1oBXAQ7fQCPgN2ijodVIavVTLcEYa6H5sO3kSCnIjYYX0HzQTGqVzNOT
nsNpmYId6ER6+hFnkR8JBOVTtFWBmgplZaFVeqXJuawzuqtFDNFeF9IYEhu9Y13IsrWfDUuv4r6t
A5qlY6AUTDRJAx7pXPg2802yQLObCg7B2/0fNTpYKPDYEYCvSa1VTrBcH1AE3nqLdJf38/ZB4AGM
RciFrO6uNUwhrXafH10DQCSX4Olvnw8Pq6UcpJYgAP5ugL66PJgyXPak0VySQo4S4I7XsXfO+WPx
oTEqS0oY/K8kEyVkfE6rSy5aPVSlq98heW5D3n62K7MkzOfu9EjM3ONog8EieqVqbx0qmW+wktN/
VfHK59vhjnTtQSLVcdK+F5JLt5v7jglkLJKxu2p8VBPcRyEqUfkx925vEcYkcJYzS0C6SrQlQvSh
rZdPyHjTMNjIj6RRXSMjYGaikHAe1cqjfm0CfwCM4pBWWeE+IP6ZoKMix7vSG4maF1ZNEsrRSFdt
Ea4AjAvj4sHJUyaCD5FyrEPLRDkUffX0dWeC5rHxl5iAGddAmO36/bDqNYKXoQCEptw/Aniunw1N
e6y0/WIniYyLBX/EPhm8wLDGpbeDzmDukzITuF+2KScbAvrmsAn6FjBC+1kxIhFV2UswPqVQbtOK
EaEzdivpBg70RifxW6F0CEr9ZA9N3NBv9j6GhJFan7iB1dZl3NrwS5WCUWcHqPMuMa0zqRwHnhd2
jzXVY2R7fYXTABxvhOtR2q/zqZXoFBRIPyDjtgXswrYacWTdKgSS8DBUKt+iV1VtCYCtLXHIxkzN
qdUODEjHNHPducpa2OTqKmfkNt3rd2TL5Dg5uQ+I50xSyFqwiea+MB1NzEvzTvyHMChBLhCx91AX
zTSOQ6fLZMxW7ke9zLfbchgfdwKCjDrZiY2+nSh8/FvmDPqgMSKHEPzTwzngD7fDSWDe6NpbqFkZ
/4FLBHUi52nEGEoXJZPb+KEGnw3I5RCNlZPZFQCxv7ZIeGIDuDTd58fvEOXtRsKZfBQUnVFieXrY
S8MOlG1KWKRCN9XlrRowk42fKC0z6AZ0oAZKi+IwNwpcSd85diJmUPbM3AqTJ1YiGc/EWG4MUEb4
QBFvDUQ5WjiZ5LF9gNFi//KEPP/TLPMaR7UcjAV54sIrNinRk8u0EaLW862OFRQAvOpXhMFkxSuR
WJtV9K8kNipKx6W/xPXQCOy2bCSb/156F1MLW3lOSTP3xAJjZbTKSZOOKWzyfIiFogK989YkkHmr
66wY275AE9BkAFoNRKFcdIYV/3i79APV46BSRyy3YcLfl1m6Som6HNeY4BQ3CS8xLUTw3zakxqw1
JoDfPl1tiOSLIqs3YN8wPa7yf+C9Gq58y+2PXYM2Eeyew4WKF1fz3U7UkmBgQlCzSLGAJNLNDlly
0Wn4t0Lx4iIen30cGV4Hae15zYd93Zrj9wKTZqUuy6A3HFNXqU5G/p42lPbCSiLgZNuN1+gj7H+v
AFZp8E6pBoe1RjzopwSRXZbpwfBEbmBnR9x9TQebbQNwF8eCo04wyq+bSxsw8CaDEWkO1t2r38sJ
RCcoiX/z7TeiyxKUYCCeuVSVSlfFUVQcoPgN+0L4hQTvS1OD68YYF0cEYEtiN2J5RM3bY1aFcagi
k92eEQhEcPXH4yOWUbcc2t9KpvkUxhWazaiEts1Ib2Pup7mVgCZ75BH1y+faiLl+t6T6Lol23ERN
pZpTOuwYrmpN54tKYwwr7lda74ZgFc2uagdAY+5J6pakbTgYTgs55DyTiUV/wC57YhHcyIJldEdF
kzzaW0zq1dMZnm+JqDiRHRleqFMwmc8P2we3P4tw2Ohm7iP8ipMTajycN1L/RBHQyMlYr3RFGaoH
57E5kc0PcHvD9mfcDrJ4Aqw1kXqCepT7C/eXoPMh8Mo56BdjntXKvli1wGAKT/jR4HLB+mkFR1gF
8hE/He5b0l7qh77GPa3UNeIWm5sHudvbe7JJ0p2GBIuzt3LO9ohCuB/DzyTTRvON50+RRqLcOfmc
3HuK/WXL3KJiLZ8Lfpo3P7aV3nyce2XDKdW/QlU5xj/zINiq7eziF4LA2oCDXhdpr8rcwMNIdmew
JqfVfX65iC3BpwoWfFHWLxZ2Q0DmCkfHnAgk/14dNfYiJvwq2sE8OFPl2W1eJZvWw0+WMAylbQGB
/bOqKqUCf9jIUQ9Oqep3E5mHjbR+yNE0wHnqp9qdkXXrRFia7NXNjP861hamnCcP8P/45+V9XIZY
xUhW/dqSf+cFHvSkG3ipW9XUrnBSJ7qI3SVhabyd7ojfkQSoFgPnANW672vP/8rfrtKBfO49N95j
TUL1ZSqLiieEvjZUAiK9NmR4SVGiyRbnIblzBPWD+9V6qKn095pxph5zOVPfQJdo/yuAtOHe6h2m
Z+BW+cod4P23ctxJAw8ajUm/tLcvIfShzQnxwzJZnUJgdPp48Qa0ytOoy49XBaxhAg6GOe9KVkBS
RfAbmb4ilFxDNeYnwM3rfcrPfVxNuZPxlFCAP2Hxm0nQnPUUVLxM/pyL1czdcm+fAGipT4KOx7O9
EYxS1tQd3YFhHI2JG97rccH7bz6scYdvQyX2+1I1YaT0EKD7k/ZeuW02AtQ9oJdwvft3T/oHZfN5
TdEXNj5WaSopY07JurrExxGrc4c+v/BlPcbu4RFUhkCHDnadWyDUth4Lypy+aftmYal+EgNRMCKO
CH/jUJk7ZBTacwMl7NgW7cPI5cfH6f3864pmYqCipReyVx0b3/6spHevvfHEDeOC7KpDHgvwsZCz
BW8RkbtydKbio+o9ZIrlVXfD+7QMi31Bpo3aahtnAMWzW+FuHWvfsdppiY45dgxqJWMjOo5TXw04
gXg9Fl/fspf9qjlbUgAIHLO7wDIXz0Ri50pP8U9vd5+uRfH/OGKxadEpU6c036N9OgGjCZHBTLBE
AEZhUeKDyQpD2LOBfSd0fBomKY0zjPj6m4tOygtnY5Fp3VbfND2Q9iey9m2oZcgrenLd+t4yv+tW
ezr/VnWocigkGli5Pq78S4LmVSDqMBaihkIETMSv6EsT74qPo/uHCaF8fx/80hX1fNHPoZYXpvtr
H6WyPK/n6Yo9pM8x2ToMIobKhARZ1388kEDzrfZ/QOdYDrVGJ0I4f6zm0jHhB2Hy76vSyDt3sOO/
OUrAwZHx9qeOGsU1KpiFOfriuCHXPTqg1j4OQMS8QGsmS1bT/uGnpGQK6pQ1qi8+YxwGnkDn+biE
lTPGaThtN3vXSLTAmRKgII2m89JRCzuUT+YGw4dDdEUZoSskc62T0jt0lcb374cmSBN6LxlPpt5V
vGSXoDOQ9rlzLHrIKaqgXw4gYERpa/LbWnZaBmoAch2it7E0ajT2I8/ROaK9SOcgcUlbrMkya2OS
ricKttB2D2PsLtYnJWRxmygVkuNVmx5ajZ2gDPZXJFbguaLcUM5deqao+lFTYC64zjwOCmWW2d4W
HRBrlE/3gl8H4Jc1qhYEneaEBUgsutwk/kIvSwoX0k7VsL/s8u1bvjLUEzeOBNqx7vANh3txhRaq
PV6lTtOfkCZ17szUsx9lV2Mot0Xh7FlBiOu3g8fSAubfUpIVZcmrAWQrik8Z1tQfJaYQJxO6cmua
O21SJ+NYIL/P408dcc2AvEnANzuvWoeR66LHfPhpUuzyf2zxEB2rE+++kNwEnBPo4OYVwgfBU6a8
3O1OizvfFO7X1QqoIJ2dDYRGYinX/C7PqKtTrKhriNJ6gEqBq765TiAkdr85A28GEbe4shdxrdto
IR/hGdMeD9z3hvBQJzOER6SlxD5oZi6Jj5xCRvUyBkPuiN19Ji7YDdIzZ/foL2ZNXFuMfeHFKy6z
St6WLRG8qUbjxOfUhj2mrzVPdRVxpi3LCMs/lyS9PZ2EqF2ChRnB9YHufpuqC6yBuCHxEak1zK4I
nzAotWyKlqRiFfwCuslNGWwME/1SvrcP4/kfut+EHQ/0T0ekv/0BPxSonawE61cUwC5syFbppSaa
4Apf326UU7WfB9mW+fLkCe/gQsF6o7W7uOZ8eN7AokjOfl7TynfeczGql4keK3FtfA7Kp6rGrG9W
5CKPRFOQ6xmRcrju6Qgj5NWl4t5T3L4vu9RAYW61G9Hl0cEoA3QDHsO54O0QEhWZb9HgTdp+fwNd
TIGsG6a2V2u/f69tfrqOOfjmrMEC3GJXXn5WgGRHuTUalSHd7nseTBD6wJumeaP4pRQ9Fs0BUiwb
VJlpicb3VivyaG0V2vbw2cWg79HS2DCMyO0D7MNiK8pi0017jZFJZOdvxa1e5qp2mTDq+0Bmx7sG
gPYvqr4Q73fyWyK1qEq4TNS86xlG4p3XeuTC2WE0GFfFkREZB1Dp6/YpKQ3Echmnb6jI7pv+Ayit
OR+1qRvWrZ3bEn2VF6qsH5QnME4dsNHNTmDC18+sFVSWbB5kEm2dMcX2fogjhm7W9QG2Tmqu1uHc
jYIJJKfsACcJmtKsOcoEcCQDlcl1IHgu2JGCxOL2j2g1WRVysq0prU22zULqmCkQSGxp8MtCI0fc
wvLn0YLiIXFjMCknHlvvcrboeLg/RNai+2HFnx1S7vVkAiEm5o9WgbEwiyUWxUO3HaamdRyDPTcU
PDpJvYL7HbCSnlwc7SYq3Q/tip3YZmcjQmg/5R8XW+71m9aeBPNAg+Ot6qdaE7Rg/2x0MaVggl4J
7+oD+gnvx/eCZbMbuyp2eHd3gqNuKH0O64/7OlUri3IS3J6OOl4ogu41OfYMsEy4n0Li3J7DU9Qr
zTvyr8UmK9ryVNoytAMx/Y4aL5RkNgAgk15ne3OwLT3Gl/cQ3MNyRuN3/rIrey5bwuBESNFh4DBX
Rm6tU+Ho/Ijnlbtqq2Q5xT2oWEKH3qCJnoMuQOeXCvswUZaU/4TLrvA6PeiJ+KfFLwXsx1uUTI4l
eOgWCdGLMg/fWGYZvFKUtng9ekn0KrxPnnuDawfQwUzrAqxYJlPzMDHmxiTEqMj7LrTT6Jv5ZIhm
f4xe/D5hAo7l+Gnn1OrEQANhXomiqmFiSIjLltHrCyQtgmlMh4++sxSqzxY1ujdIihch6DsWTY73
pvjxXsAWaoyUzce+xXOvB1IH3CO8c4DWvTqdkr94d7ZiX/n3nBDALfPADAmMbc6FaAIsuPX+R4Zn
VSK85S0/3pze+kvLBdmgBp/AKfxPHpru/uysBGBb4LNZLZf2ws5pG1ieHpRsYvFxtQEX44dvUkdg
cTQ0Z4tEv1EOKcQwnl5Mria6YoC0gyhP+8GnNrTHDrHd9Swn+hIHpMnaPx9p9ous9qoJlte6C5Ck
5McZz3f5zjB2/WwFzEh/IrpBnjf9G1WF1TbRW81Zq0wn/9JSUSC8S7uo5d5I8+o3QKcp5WsNwwNu
bm3tV7Tw5X0mVFd2HMvHaUQW8vpZDhtVgoKKl8EVsdfw308WuHS8XF3x/GrI1kwDaZ9BqArLj+8b
yVzTfwduID422xYUowGFDYWzDo9KeLsKlfu6uXVzxshH4V8IKQavUAhHGHYA9lMl95hELuBiGCD2
nYmhjhgaFi1OFLrlM57yHEcnpF+k2gPUqwk+yiK3A//arI+WLkZcGF1IrybAn0ztuXdOHnvSoxTl
ikr7xOY03daSONA443bKMVQaNUOLrnXiL/mIusFHTM0IcS20dPWVeCSqaInb3thruG5YzizVhmxZ
YsgJymSRK30O1sbdFlzCyuGjO6oQqFz5s0ns0Znook9ULr4ANp2eEbodrJ7HDtjTED7Up9uQPAsk
FvnIZQIR8SwP5O3Qe/7unmPDy/fjKzQNhDh7KKi51uPeeUXeSmZb4ntu1PsO1q43fA12vMGXrq5f
2+mDjD9wY7Ry6k7zNEeQ3hF1Sh8me3SGJo/nNMGG0pMb09JO2rS/+kkfLfWbg3n8dz50LJZjHom+
+LBvPJ5lk9My820CUM/dIxJRV+l+2xvJtDJFMePAjMfgHv1U2klgsFFfBJ8PvWBCugnXJGBNr3c6
NLvCzur+KbeIJqix1VdOJGMA40LdGD5rvIzKpSnq+g5za5Am9+ma2c6JuJjh2S8yUCDJnwA08mRs
K+HCtTbesDPoCPPnKqOSIGyFJZAlaw9GyoyVyFckHW7nDTO4+8TVE6GLtLPZ8ehldot3YtQZToha
aB+xf9L9UVUZhkL0PZcvkdOXooWqA261m2mxmED7KEqmZsetXed5GyQORA1E3PP6mflcT+7Xy9kk
Ayy3B4EdhgbFb95uFsRpN4SKqCXrzMYKJfsG/zp0rw0buRGMi7OOvMCpIq5rWmmF4z+1AJiE5a8M
LiXehk/bIyxHScEkShrtJCmwVARnvmZWiakihx/pTdlvFrcUqHS3HpsziyvRhPw14go571F7XMwD
CS7C/ufrTnI7cZ1NbL4wOgeWdq5g84yju+ECuB80GgB5ulxzIDvWkwol8I11HVRkAMx+13VypZKz
fYVAqnv1Mafyb9GB9dXSPdhbT8qlSG9frs3lBTc8n7r+0MCNj29JTe2dCikGtkW8pkwGogFQH1la
ifkWCMonGPdwR9IUxYlA760Fyhc7CHBa1/zLHZxFksGalQMC8Pe18fhaO+3bVlig5t/d9CdJkchr
vj/6XdaS9tK4vWfPn6M0UOIEqGb0kzp4SEdUQ+rzfu9iwNzxTXolMzraSl3qDp7hOzM7T0xwXAuX
WZ2vXY9+GGrZqcKuxbHpXJfBgwlumOyDRQERjUCM3A8jBpuJ7LA+w/MSfdVHm47KF4cSaOalstWe
VPebvdewn2H9a7IQ3WiDqKPJMXLDVU25TtoAEJrjseH+o3SApVQgtTRkDbMgz3RmcowaAsv0I1SG
Jmdh/ZrX3BH9DABRg9Le1jsh3PevLpVsayyAQwLKh98WKTyxh625D46bGz4QFewpLRNH1Ahmz2BW
Rt+h4zhYBBKVRNMBbJRMGqt1ZjNS1GEV9XEtahrnR+BwF/OUfrbP+lvvlAaCbncCdLL7Ni4pYvYU
3advdGqJCCmPI0OJ+xaTExvICfMD4h2wR2NdZvRZwBmeuxh9mH+1jz6zsJUBn4jw+WGit2aWLHoH
NJMyFV9l8C+DjOkZ9ytzsKlZ9HAWgWINyljzTCuila9Wf2RNXlJuwDj3HK9/MlToVLh6dpl6OMT8
ZcOEywYZcrrBNyJpChXgiVM2hcTGUFxDv1ayEYW+q+F1kKewQkkduNgnjx+zFHFDdAHbyJtVdznG
BQMt95P9n/Dkrtv3w/BbJMUwXihnBNUcFIvC4jh1qW/byTnGUGZnnuTrejxEy01RNXW2dX1qQABK
4ZOy6ajJX0MP0b3WzNUN2bg5N8BorPYRdoi17jH/YiuGF9+CkxejZFr5Qx9iHtYHoxcw7duJ8wv0
sJNDvmPrPVn3HpLPTadgRnrsWNwBav/c9yVG2pzAMyh6B4LjDE49tEkptGc8Gy7AXbT8/FjRVMx/
a2ImdI000svRomsDen0Jwy0dA9CbgdI6svj1hHBv4cPPsRrUXuiokM6JaTOroZJFGITvbT/VVDuq
05XQQW+zIq4LxhKz966LmNOYh/xWycnA8wt+wnv4sReat7cOH1AVjQTyENbdfrcTSNJIQUakibg3
66VErKrTOHchUTMcnEyGq57fnO/RXZjOYS9Vra4ZIrAwn8kqszbyLswNH4x9ILWcKZQe2vOTZCsG
ibfdJ8Zo4ITjUJzJUqNR2wFfOKM0q4NO6XH54xjRDnXcDKh5q+JnR8tUx0LVNJfw53aPRkuVDbBq
2cAPd2yVjewUlWSi9VyacLxw7NbZoyczhc2YnmN7KLSzpAtQbU/TeMuCLkQVnlJwTDFbCKw6aUlb
Jjb+NBe//9laanhTg6LeLHxSi3SKgExRZ0H1huO4siebdUzMFTFokqy8KgytAan9p0ezxdWkdPly
RNHxTqo6qnvwvdRW8lP5y04GJBzYleRHl9PXaYF8atyxAhi0sJLG6vhXfcTpe9WLMnP89haQH8M9
NJB9hJXAOl+oRAmle5FV+FB9Jwa+oCc05YXLkCSshQkZhx1BTYeqkah9ntY7d4ewyynWKUejfAdN
77B13/kNtLpVJ2Km/zajy7eg0w3aD9AKmShkOdyqyhp1Rr7sxaSInNm7HNnG8ae7ksTjoKTnh8eF
J/tUT4QdfZouMrbAal3+3//hqwnJuGKEM8s73Adqz1UPJQBk6aly9GNnw/5mWB7AXgEeyA+6Dgf4
nwV8yosDEjWfAfwf2Dj3yRv8m8JlzI2U5sOkzpPJOgWeILjczVWv4qXlfG3qjpktMTKEnxpEG5qs
uPZxj5t8NtdEP8gqojFbOK/6nrmBGhYfPi/wT3sh2abNOISHDL9yC+vPTB2ZoYJcY4XLSfKOySFB
O+WbKcpdGL+mNfCCGN0eY5pCcYxswprtAIYOnVu/HV9zibXKRbeZwFGaSi3olFwV8I82CS5XJwk+
aFt95tChXpQDPcsBms5OpWays2ZsFIY+6P9djNFAtiz40wVKP+ak6nKCgXj2s0VVcj01wh1OJf/J
HXYU+2mMsNX9V5txpOzQUgs1m17JTVnxL7vwzbGDi+1BmFgmUKJlpZRJsQIz8+dASweHZzCc8Zfj
uJLBxEVL9/X9HdBcJbj9Q1PuR2CV52Hcv8hzTV9MlLF+pUbAcmni8Ay+2xACcjhUcUszWgB2b68a
bUZXKMnJoWsLho9kBMZTzHiTnK5JKhHuc5YAroxdZFnHaJ0kS0Wf1ubdzC7Swe0QQ5//wcJY9uVv
8UJGlI+bETkZMuce69uRPo8oEyD46KAEACV/dMAU4tMd23VjOpiCWcdRCu6w/TTEyDt9AWaTIMzz
QxiUYVgl0Ejf8r94Cqy5/gSATld+/dhdaukis5LY4TVK98AFyK95CZuNR5HemnWl/RLFPyH81TYv
t1eGgKRR1R56/DKYX9fm2r4mdDlpX2iGDX4XxwFjJqJ5pLE/1uJ+plVMV/3EwpIKYUvHqlRAZppv
Hd2DFODX7BfEqaP+zH6I5w5x/xLx3rLucRRq7qIj1RH9UWL9olSOcBXfx6v4FQMkZWyniOYcdjYj
KAONwMYUCvt+Dm57jPq2Zy+36bo92u7bgDwCcDc4LgJm0j/RunAqvIACa/DlJ6ecxGQECIFTrZNm
7tD0+/PWN79FhZNVYsw+dwBjN4Y3+x2YIU5JG30hv6HxjXe8q5aTS57ls70Ue8rGwvtz2Jl8sjSb
FcPg5eyaljery2o8wdqM58lU6DZgYeCf08FLi4zp9l0JcxYSav2cTFu9plnLasUPPj2k/3x7oaWO
6h5gDvPFM2NecsNEwNHFJCo72wKIEa/YBgyNObb7waU8w60eZOi3cniWdDg+N4Mo8hgFu5ePZa/e
1Nq4q6EhQHpfcGNBbJxGoIazgW+yg8O3L34ulH85CJ/5/kU7H7okTMVfWZVhKVg0xwcKC3CukmR+
zmPSrnFHZOhRLm0HDa+jJpd8UEEnnj1kkgLFmNeSQS2Yp3l8h5F8HxiXNGGexjxYPELOocWh2981
eJlzLse+RuiC14Awvhxn/yhiQdLOPWZWi87zU/WbxcmmcccfV4Nlrbe1aUnrznqMz5mKHBVNLzbn
qaTbqUgrSP4dLElDPxmVKJ0TC6plHOt4G2bvKAS+D9wd+dwYfoM/ScbGcLt76Ag+9bG2XuBScZpr
cQZe0ZKcIZxIRWvUiuTha5raNu013lQp6EtIc3p03VJE3QuNMnDHB5foiZtnMDk3GIsQMGycygOB
PdBiO/Aw2tV8ky1wSwUMkJHxKytIRDEH6eWJb4gzuGX7iXMYHintmH9JQjh5DSj/NyHfp22fCFJG
jh3vBofLV5Kr/DjHAgFRw/lJposqmi8LY+9bbS1tVCWyW0e9IbFNV10BRCTFQ1G5aBMIBF5W8i0r
ZZ6BPxy+IVq0XR7w28MiQmLfNCvW8K4HFXL8ajE6Qwsol+6Kv4POBTvtbtNyZlM21e2gWKw+0uD2
8+FQU+kX7onxcX3Aln1hHcROKsKNb5ntZGHaepLFwkQPkf4SMQSd3KwbU8y4HCEzSBpteeWLDQ0G
DvEoFG2XcezJ8KKmNp8LIKMey/zlNxAlwCSH/wH0L/D7ROM5IXxo2aOaCyllLRyoucUGVhEUMcEz
rEvBo0K8BDDlMXPaRIybNztOjJVlO00ui/dzaErUdQdXyNrG5uzMN0W+1Gmt030iW5wlbqeBjUWM
SIzJPssbxzAcU3v05bsd4+Pdz6utpp2VkCPXdW6Ehv6Jbhl3CRGa8q7YvgQeDwxSIsvNUmWq5SkO
MxPE1uJ/yXLsbQTZQCQr2m/10inMD24Nq+m2VxY1SJX1l2rptdCYIYoTES2jnQfevUH8gIFrY6PP
3mZCBUvW1gDb92gR3i0PtlssYyfJY3PETybyEsfUtLJfcZku5OViaLt6Ip+ihhFf2NBkn4fncjkz
e+jxdjmlabAbH8Oo/pduwzGIXrcwUIt/vueOstEG/wdMwBSeASL6B6uVkxIztflENqOPuXaeUK0Q
NbcsGcJQ2U/9ogKXfnOnPKG5ix3vJZfErErOU2TyCWT72fJVnDj7TAA8t9+WvYaMvX02wzRyDCh5
XxwBMQTmNCE1TMew/cmUlGC/fR3lSNA9WcSdkNOx7K0zgB1fg5jSNPhwZiNyTid7hfoC6yBqNtBA
z+VUhZUp6RpSQXlEzSuoS0YM0AbSnRwAFIjWIegXiHkK9hUjF+RndjjUG5lbAUMN3oXUhJ+5zhQt
aXHL/W0mLVpLLt57eOI3zHzeyFQe0C2cPQboAmrz/21R6brAhj5ew1NrF4+AXw5HAt+wnUBa9Okl
W6n8LgUnvNvl2YPzzTWXft2yqsikowLLrsOsD7QfxsixZa2drfyVhOJVk3OG04Jn3jv8CGkzi86Z
2LalWz24MEMHY578oqO49lhhw8GzKeR/Vseoru9dmtLRzZ1lABzwgXgdxYCQ0B2pGQ149qG6dtn0
AC6Fo1nDqF4qDHmNs/5pXnK9C6M5tvRCOEHCjq3yZnWvCiPMxBACn5R4JJnqpeS9lQ4eF668Cyag
P9bc2XbHmCZcQAet6n/95c90MmrIJSl22EDFkasJLgjCFoypQwFtK2SulhclKf6lgQen/cJhHmN2
iB6XF4o/SdIptb1fL4Vf6zpxhLOUQqQTOif7/QHuVvK5IzbpGPaEbekZYBZrFbbJhWQJKB30xze7
qbmbdraNKvjsNCafCEsQBtxi0ugmIFKg23gawYkTROgU3Pwy9jeKc3T1o2FfbZ0wfQwMZYmffmYM
oMsSPgbaeeR+Ejbnhv3bCUtR9ALXoxVj2pYh3m25KiY5c3uubCWjpthw075p6N4lY6+KGBFiUrRw
x1upv4HrOBukBUcE+3eF3zE+fND2Sa9Dtp9HD8h1JEfDCHJllpSK+imBB9gFrhvB39TkN4lpxcn4
fc9EnwVa4CGbZhIWVzM+MBI8GBy5tg5JzLUhlzlDLrkpYs1GcQgsUXk7whtXPVaql8E7TSViSpc/
W8jQd3aTGMTh+dyCTOyuGXSMWReCc08D+Wm406wNlAcE6ILLsRfuiGc7YLrQgOgKYYC/yV4Jq3/y
m3yVFjftYP2iXwOxR60VmrO7fYTbVKt8rlre8c78PEM4t7f16BliJab3pLM335j6mWaXuNGBgjua
n1341wZhvNmWYG7chnQhw6nJavh9Y277fleyLJmr6UR+8LTq9J27zKkCc/qZ7nWRiw7L2BVDVsSc
kfz0KQpUE4/xwxxQLzyAkE1KjMFJZ33zc+njRQZuQT8Mq0ZXsw5bELb4hVOqJnw+kcSXl9hUExvG
iRxcXj8XYPZB6G3dyIC3MLhCnhTlUs1MScusrcBnMy89dVxrkLLTvZkyG7SkPJ7ZTyRjGcmTp3wu
u0w0sdiwhGSlfXFJshwakW63vAiVTYm4024ulcSledr52n02miZT0ppLDH5QvE+P+0Zzy6zfPq74
J+pGbOQ1Iru8kVfYE5OF25JpJhPjC27IpL7ac00JFxMG1Bg0VsXU7tWyMdT3M121lLfW3v3m/SpD
It3IAgJCNHG4UOLc/HJ25lZ/qVXPeL69dsF0z2/9D2qXVMI5xVgBERSPFRe5n0YMJG0fDiH5Rz3D
X2nawU9bKuUHVoBTN/V7ECLij0OvVQeeoS9361ySUuK5ALRPXfIhzvZz4lfyib6u9GNBDhoGZkN7
BYd7NVD+QmVyy6goEckC4GaEump8flLZ6LTuOSiRavbMxXbzQvrA9RXHyflmlaYtoQjnFQA782Jf
tFhV0AcZWQw3TfpC+uoq5Q+Jcw9+Wc5825ZzZvbTGyDPwMN1dqhDsW3yYxYvhayWc0XDc+uXp1Lg
Z+j4hvvBhsHaiV/ks43Ziqp4Irr12MCziD4Jw31TuovOCEpaAopa8JZeXok0ONN+kr6dnA+OqqlQ
SwQkc5YxXX3rKXefja8izBFGf1XadL5vz+bmAPgr9Lv0y5d4iyvAgBQ8j4Nlyiuzu7xqAP9RLKCF
MTGfyWDRNMEMm2EofJSVzst83aKTYj4L3GnDxNKYzSTCX1W72YFV4aaEiEjyEuXngjkJ0uxsQQi9
VyzYux4dyI6366tQgyJ25OdDV6Q23jM4bUV+pt0dIRM9L9kfGPMhcY2Tw0HjLB+BZmOuZ3NVpq0g
XE+qvPqqYxjwWKoXeiN8ktaLCbMTAv4sDJ3n1qcmwxnStqCR4lrS+P/fGwQfw2jLGamRPS6GVn18
rt0aggFSfVw9x2AUgdnZNhAfe8WHpfHvn+yHfGqbbzECjKEiQlV/8aXJPmJawX38xOUyziDG7XPR
aLXiPwDqEL4rqHna8ufr1oJTFzvAhs7+dibaRKu1hKGPZUNlNyhY+ZraBN2G0Jk1n9chvd+Heq+y
XL+ilbv+0i+emNHgzVk5T3PQts4hAzSVqys0rJaAhz8H/2/eLTbEFDkTfi2TvKbjLx1IHhETSNHQ
HIrQwiONxrYWC4Gb4yA35hdug0ijTRU17p8sSJV7TL2cqrBU2hMIct44JpzAfsE7jHyGdOxfYcfM
b4v+lIudJV/63bevJGkUAuSf5nc3+jl1sRAgRfXpOtyYOJXNjC/Y5AygY9SaPtMADvpP2nCfEGay
qZNmNRm8lf4AjyDCsuCJpfVoBLGGVERS8+4yzMpIHtme9IIJFGuQXIez9tHboar1pkGK+2EhNOw+
dseoepmrYVmqIvulEDrdbNBa0sMJxsUB502ZASEJpylpolGOdwlWxqvQ9zlzi+MDhCvIBAWKu2IM
SVDKb7+V3vZQWGNP/ZR9vA1oVCM0L3r97Jn0l8O4aVNXE43K625Lv8Z7DaDzvyiWJdXdF71D9G7e
b3DPPhC8RR7W28oeJgZaEsf/0z9SmxIw366n05ankrydhM4GOdyNppb7Ks0WQ02nq1Evp3gwwIde
GHAxYWc5uLTZ0oscF/8BPxV3/fhXEoJe4I5t6HzdHcOR6cI7M54SqOjrqYW5Ra5qDE38idWfU6D8
2nHyDtxvoO6SyUY81qNVHeN1My+GkNsLvFxpse7QUWAf8HokBzBg6odVPLaYiiUgKUeGcuzMsbFd
ouSB1T8UUpFccyKOVa9FetNsQc1lTFplLjJ45c1NWSXBQAJULWu6AuYZjTk1BQeVTnd2zq6OjMVZ
H9welki/6Zacn83gHZGMRb8Qu5VTewlqK+kri3euQWwRXuijzlXYSOiUFHHq0mOAT8hxE0ZDgmTt
iHnM40fAkk75darSFk5T12Nlq+PkATsxuctLyGUbKp3jPVg7gb56rTUwmD8yUcw+OxC9DFVQoFds
PygF1I0AqGf8wOamQzmDt2zu63NiTxVhzUy2fGnwkcuQv+33NOGAD+oAQSsmHSCK3p+1k/GDMGTz
VSJ+vU3z9jhEgxQgq7ugkAEOgMmLssvrfi+dm4m5zwfKoWLmFaGRhr2SypVRwQEm6dbzPAZLzSAK
fQ83z4FYCINoNdyD7gQNYDcv27Hxy172x/+UmnS6D6UZhfLQnEUOlJ62rtwYriivca86aVRQT248
EYhdDISe5modldlP1KSknE0heU+fAZ0w/KG1fq9RLAh2amEzWYNug4IQVBtxRM0qw6FJa4F3izAh
QghVIYzR3MVlkVtj1dCklPDCW9EsnsKDDuFKdd4n8ejVN6GmgLD6o7uTsju6BFab559Ip9x5qJ8q
Th49L/RLc6DFzZyTWOV5iDgoJgQuGSZE7f3S1nyZ9TfYyh3s6urRRwQwAZLOSEG5qbItsDaqOA2U
vufWHM4cNj9TYVw2fHD6autysHwmMIVb6DMkAnqgD26wF5Q9Z4VAzf4XoDJmjKyKpOwJ6jJVw5vI
r4iJsPrHjSHhM9Y/gB7wuRgNqJCOYnSPiJF1sCapHJimELnF68bYWcqTQhgZwJ5c3iSsfe/96l6u
ahIL9Q9EP2+ll1y8w3knzPJxteNKwhFQqxJnGzH1dYRx9HoV4OmZp4Jj9ATMpGAznKjodGDtqLhf
OocV/oys1dBkXsx1rScnmQ4qxctAlDxNoqd2H6kWQQnzw9+k9a2KL1HgL3Aq+U2eaolo6YT0TrsW
Fey80M6TpBs9ID56z4oiEc3wm3lFdJv+RFoI5HxrhAXNeVb2Zzds0m0VygApQx5cfMDYyZNeUoMt
dUpqBdKZXOpv0jiVSXLdwBjP1SszapQq6L8plGY0u1dB8biwthj9ceKNygvd1M7AMBJGVib3RqTo
7pd9Kuz369sXpRUMSfxxWiozmtJ5MJwfTKtG53oOqDJ77bLHnmtJHsMazijgnQZrd44lNKSR4yD6
4CxUM/R/5jDjbJdGQ6QCX5xOKPPgZ+KpxO4NnSGtDRCVQ2A3tYv1z+Lkdw+OmYD4a9RJNLY/zN6u
j+4F6jyi/OmnpQZpbQO9X4Cce6Kjp96xyi5IAJFxBiDpfjRWZv5YeTtpJlxlOc0+cW29NgbKSiyI
3H19p+U37/idAbsWQ8M9jxyYvSNpIgZdMqK7+n/FcWoaJjb3jDaYLubNMZw6KD6dGZVW+yGtrEge
R/nY5yBWXQUop8poPRXaba4/mfagm1xkQduwXPo4YrfLU2OYXHBnIlXfKj84BCLRuiTbyGWO7Rmu
uevLSyHCu/zLWVW1Id8F11W2LgDdmRCzj6drJcN7NJFXUT7VsK6QYzwyFd4W/P3+MEjmdhHu1YhZ
JiBAa71zebgKL22N1UsWRFvbIGGS4mcT+6Pnm7zBViloZzT1PkCnaZHJzCjiLXLmllyx2nSi063X
1hBHjYqsDjyrFSMCoexLnLn3asFi2GrQ7B8EMCsY3kDGtmmdNmglSwqag4HZwOfSxJyE9gXM93BT
upIF82fCvGA6fND/ZzZEOl5IxFO387FE8jWNl3GxVI6T27JNhWTYWg6XVN3mTVA8GrOqkBOGfkH5
n1z9MEBuynmyE/S8J3fTxP4JOEAWs8Xfft/Q3bsjx+/UHmrriRmCgwY2f6Rau56a0Wqc+pWE30w9
NVP06IuZt1v5A6QxIDCOMn0laTjPJFjxhMPzHI+1/XsR0NWkEP7kvXDj3T/EH3PX6wY6il3nO8ti
aJb6xL59D2lLEvvJIBy6mVnR7IFRLY/iy3fLi0M7UAvnP1iVMY7ODEB4LnhyUrt05WRlQ0hnj497
uAoZwKDnsFFSwMHz/exAiqi596UJjKPYqWJZ4HdY43/zlUX6e1kw/IZuMdCkqw1eyBRTl09SLB+1
zopMg/QQCgb1OYX2xcFZMctSQdgWXzVg4Cq4/xzxBfCZGWgxHzOacfmcNMQbQoNKR23+01J7VJvb
/lSDQTd1ZFd9jXKiymIOdFX7griOJzKCrnUy67kWNLpNFvMdbN+n7sRIihAmB4HdohbOSD9QNnb2
VsTEvNphmVV16BoojnXfXrQNcUJ95PY0VF/dD18fhP6KQq759Dg1DDO7E3jcFthJUu5g4oB1NJ0U
e9+wBzsPFzIN8J6B8XVURPvt3R8uUONPi+zapfCiQZqguDsKt+YTMStbP6bZ7+wVQCsLUjqmdkXS
ijPLEgY3oXoVtGIi2w/dD4QglNes7ybFcGnr0y10or8ZvPVek0Xa9PxhQaBO9r+9Ieb+wLTm40Ci
xZdgnqvjZAW9fhCeS20OrcT7FOh0hLreG4zAZ1+RxkGgWOUMSmKLXJ/Lmo5q2mfrz05SQEb3dkDe
aXxEO8RPsmKSBOE5BRQNAAdC+H3GduT7FEYwj0U2adr58BaRWADxgza6gKp+kRJD6fRNgW1ji3Tl
DL2YoquLFyoG5qaC9eOrXC4TapB+3bWWlv/c/ymGY6rnQYsd5/sHuXisiiaQjmpu9WpAaBGTLgCV
Po52gg19bSK6hkBYu6GOua24R3lTSXTkyn8ITjDvQ7maM1SY9z0WTgRyNM3XXe2Yen/S3Dimih6N
TQ3gkaFinXWtIcasgS4cFJIJ1W3kQfk71U2QX1M1w4rZtKOjHEvZCuHyGlMsFgxhLPHcCWoHXcgp
ZvDmYMg9wSOKQKBihUqR7gHtdqTbbIAiZbCvgocGVgmt/xXMSUpY+7f0zNO3JUgqGfg7vIJvL4D5
2ClGl/Tee6Jyq9Rw9c3XxJpBMuGMiI1U8ynlXo50u0ftLlvGJtfC2548F5oENqvgCXPiqMezVl0w
KsmEYE9c9kyA6IrIxo80WULHiCZ33+0SV2a7cY6nqSE9/RX6mkhpXjN3TUH8zkicyzGQWsll6CX1
R0nZKt5zxqf9zlfGJ+SGx1M93Wjdwp3YXxtriX6rdZ6xqlyi+jdAJhfi0CXDUsCJ3fH6Ngdye/1T
H0Wm6+DbTkHqzUEDIylNQg6SeJ1uSnhNEpP7agN3bwTqk62VmQYOkG37Vupi2fahp8rGwIE1570m
ifYikHJxWDZTtaO6pynGBpZHrPHGt4C1QTSqfR8Yj27BfeHLxiEIm7KCEO1CpwuP1Istlh4QFL/P
NsTfIbrzo8G6vEM09C2YEVifQlgA36pNXfoG9xBLrFtBjabHOnS+i8Mlc8OsVLfKrlRJnND64I4A
AexYZxyPOtPob1j/JmpDJkkRb/KI1hfmP9QO9tv142L+abJG8fjFGeDXmkX8+QFVS1pNSzca7lSo
/r2sFm38NDFkFnYj6s3g8pSvLGtt21aj5jx0rFGIfbkP5+nETAxxfy4CmYO8Co2q5KoGsNqVXS8U
t05s3ky8JGvb7Mk+jZixoa8CbsihOZdeXoZi2+BR2HXog+DQZXaLBKhfABV3v29cQyCPP/6Eob+Y
5NpaC4p+3azk8pmnAyqsJ3J8yc+9HspxpBppjf/8h0vOttleYfq3haba1LVME/gs6qA+jWun8HSs
tVQ9VgYcGwgUr8kxSBOgSuyN2c3mWCYhmVf5zveNOyFr4uEVEvPEqsuA4NvQHje8KPahF2G9UXv/
NiIw8nmhBukK1c9brJ1kX1cBAQT+xatzrbxIHhlRYkDAjg6AdosTlIybP9gJUv4swdtzdCHM4nLA
T4t4/wgMWketELOPhCbmEIjxz6SdOdBZTSBrnj9oeht76kei/a15w1eddbRhUHGFyfNDi7aSN2Kc
uYGwO84v0kWm1ydqAFt8u4O4MO6hcoUSVUyb/Eaf1L6mYN40MvWcYy3cyldtfjhcEgHuQvoekiCh
ANVd34Gb8/PhdfVWHMZsprwMHJlZpeO7WJyN1KreubZSgdukjWdkQTKqrwg3SvsBIT0s0gUKcB0K
pdYj2DGtW7ypc5hUjxRRD08isp9E/LqzXkg8owK+/8RFLlXXZ06VU7x+zl9S/pZ5VgrdWVamz772
9OyfsimZc2sXElXc0Qn6FalTZMWBw3B0CdW2mkmrXOYofq/W3xKE1mKwoVmFdKW3CtLr5gF8SKfQ
moJKoFUeiqjnwuFJpnakdwE1SE8cct1PDKXVSCNaZ2+IvDbKd1vTJRpbKhz6pldadM8hkMb+Nbhx
DLQLZhJBjBa1VU90sESsnCmua1BNZpo7pqJDzh5uoktLn/aoUrChGg1i546Bob9tUqQMJt3hEBzI
2BbeAztOwNPbYTG/uXWwB11OHrRJuXAobyUGvY49+J80bNDJiaNVnQQgRbg12SwE0I1HaQdoTd9Y
r5KAgBMHfXteoykQ6efZALtTvNtXo9aER6GPirJDUx4Aryzjt2ZEOyG1CRHZ1CwVC502QvrxThSO
BnCFEAn3egKVW32TOADV0O6HWCmfDFuIFglQff0PaJcJmkjtcR9WhErACwC6FT/N1fDKGe7gyuIx
A/o2yvPyesn4M6sR86YB4wWj1xmV/OvgmKEnVHl4B+l7WKIdALPI5ZCZJ+0k6UnwBu+BTZDR2oio
yPrn3siGWWf/A68ev0FesFvZn0+donQ76OQQqse6Nb+wzbc8uEcA/Jg5azG2RMTlEOnK24atsyu3
vY10eVNv7ETURL8DDVltoTePV8g/7wWraegTREJbcEokTZyvbRZNh4oV8u3EuANZQNdKXGHuNoQK
WpOlrtp/yXqjAn3LduInUkAvTB+TSXaFJvlKSHDPlQdsYeST5KJkfNbmm8h4Nh9Pt3tJ57Kb9w/8
bN/Zl9rQdktVdGwXtqTCl188Fr8IgxNRcb6uNcHjIX0/o6MiAGJb77WMuu66LjaGw46aAROWJ2gE
cTTEPXifNRXpIfR55F+AlnXqDqFjQsSFA4Q21QJCCO1rv1QFXPv0vS7F08ElMit5CsBZO3CPpKXn
MMfCh+tSSmFs4+op6/gGkyhc54iaYtTVRJZidFriKBYICIKynkwsZLglshBeuV6Ge6otb78esd7E
vC65QWFiWj0w1wKoXhMVJnoc/FBt3RyKLVghvFQAgs07vP5jzGVzt6JK1E0/utENCkNLbVsFrYSO
NJa4efk4VL8DliYwJRSZETJ8bKLLZi30K56XG1Ka2sjU8mhYfkNvxg3Q5DKxqgo0HB4H1p0OhiZK
o8XbUIGYCwukHB+HPR1j7HGVk8Z55Wp2U/29+OXSa84NQn1sbLTj/3787ez3lX4m8I517arz7EyW
vEy4FlelAVe5frIllycjncKpbET3iNJpal+K3Us4C4mYuCBDmjETjFwo5HIrpf0YERLsu+TJKJ90
cMqqE1lAk1yfyfGDFhb3KBYJRe8ac+j7nZT6LP/pNGTlONUZFai0EusPx3yKBLqLSjM6TzAl2qn5
QQ9kewDfjOrIKJl7ubf1pbChM6v2sNOxKViW/2L6OkySTsVDFV0jK90stIyVPzC/fq25jjctblh+
dpTDj9Lm9qFu344O1P2KhOmnTDX1PMvgQHLx+qnx09Od5znpMMgieqjzk2BpqciiSRlauz248R5h
HuoLDaCB5QAcUMHEKViGZJ99BCrPgCKomMYzx2U2O9fYfFODDhs55t2BwTVFmRqF3MzpnvQH8GYl
YLbYhMz4lQka3xkbCobWAg4CDZGNuyxRAWiaMAzl4gND6ULHPr/8NMOKXIAL1wWQGiv09klK4Mu3
tMqLrkjIwBvqTSALzo83QQLrdSsXp+gEiPk+Z+sPnBkbWOuABytXNHcfQmSWMnVrXZcbau5cQ49O
RcUuZm7adkponSjqAtCA280W+6yaDqP0WufSg0BcNUQDL+kRradC2HUxUJK12kYKbM2aSbVYY8H6
56N5MJMRSPnpYvZH73E58qqnPEW6IWkgUb4nM/XoM5wx2st6bQ96wB+QvN1uuKGuPY/WJ6ezl4lY
EzM47HmYQ7tV5nHSIRgjEhhDqJKTBTcPBOTRXgLlcke4s+HAUma5Qdmqiq1AIPdXYDm5ZlG90cZ3
Ape+SSsEUg/EFe2YfmS0JbQ9XauDltSkgRXDaZ7QQTZIPM2LnWL0CQCTp2c+R5EppzDaRuV+bks8
ExY7NBbktG7M77hz99/toWSG5E7Yh7gfQ1HL04JsUEBOUh6ZzrKPn8O3NmxedVOhdEL5ElbwK0iq
9G5DzL4EfShQOxEH8pK0fnFSBPE0Y67r/CwVC0RmpTVa+w2yRJVVNztu2pweLL08yoZP/1DMHcMM
QsiO5rB4UeduRGJg8p3xCIE44wiavUGyJarl6HFa5W4PZGULvQKA8oo7LzkiVUpWKWrwxiZK3ee+
S4VWkp9VZDIcyMzu63Vbn7iB0dtf5eZaKQEEjtauDh+cUGWY4BRiCcScYDFqeR6qX2+eXpQ3FBWk
/LPlZpJZPkrrfQsAlQK0ri+rbt63OVqIan2Ly7vSwfzm7wlDAudu3tRzddwuGjCS21cA2CpLZBmE
2u4OS6st5BrAI9xMR6hLOy9RsqiUwahVoa3qQ217TevsuvmefluHuPLL/mpGekHR4cv7Xr7DXa/O
Fkof0x4DWIdonhNhJ/WHqk2B/49CJOyHoUgKc27t6QHEO7hBbFtcvz+aeS9SFpMQwhpPAhD+OHMD
LivUxftHXuoouXIrAWExO5Brd/m1DYS10Q3YOQn55Qdouq6bsHQVdeFAiYmL9gcz2I5FuYMMgaDK
ypUYwJ4gl9Rr17GRTKYAw5xYBjiNeSyR+ZEqkPFkCU7ba9x38zzeLoFYSYB3CjBc8CzNQ6HbFtjE
ELpR3Br+3BrExn8Qp2DpzpHkfqVC1wDFJgW+Ej+7A9cakWr9Sz5zfOij+fX/+nYlXm8klrsyKAtU
7Vp1Dq+d3JVXUG+EXYuUabnt80kSv+Qozm7Iotlicp+/bNs735jkEkEsqqFVb/qyGyFPnJCg8qHJ
tULPDExhcs/jYcXO5jizVJTWfovMbk+ASHGwCDSH/h+NXoGAcF5KPN6t9uSOgPnWf+yqWov1/PJ8
8Z7gIvTXsrtXpGiX3NXvQv1K3ZbdufNUxbBFFEnQOWsaoCmTLp+vtS+S2HFrvVmJ+A7fLQV0HAa0
inN8foWfagGace7O7+XFIY4rxTQRrGmf5jch2UIupujBoDCzfvLBcuJR1tgjCp1scSM5skMx+G/+
hDo7ZMKnUXdhnBTwyoshdo+/ts9pl5GwdS55ZtIMq1yTm0cS46nAQLFwgNMH2AH0dAqGGa98ohRo
It5/tBrS/veSHkmVm51KIb/4wvKBrWdczFwrkSLy/kn3W+8MnLBVQPEcyqip/k3HKBerGy6oYCOd
QP44NA8GP9V5S9W/Zrms4SgLNA+yLSCDENCAw43gmJrk7PhuoK/Lqlxzj4kngPmRoYhDyC7Yyk9h
6t8plEOhbHovSyksk2b04W8mEYjdLWn2oKKCSEp1kgVC9K3v3QPdmxheOzDYZg9PXcm4zzowLTUH
2cA7IY2nWh+cWvvblV3KJI3RYUWxf8n+stTHQ+G9DjSSjJ8XgCxu2RwoI5sqdtKdRxrvR4Ps9Hux
VWh4NA+I2uKnenYrJQp0I5w5NV5GMjQfHd/VuNbzoT1vxCdTJO8Fj+HU4WJRjGV0+9imfaGXvicL
gLah89GkbWIeiXE9CXTeGiJhvNd7PN0bw3a5vLGfZLcaFhKqUFUFU4OOw5eaO3UGyImUPur2kduV
k2oYAhbnqvA4mz4xMe7LRXyqcAUnyjnGAU+rAlXGh0APF3Y4eGi36k2NViTGwxeWjdC37iBZUXrG
jB999p9islDW2uGozsB74dM3Z9tjdGUKWyzD9iOSi1bGbAK4rvFcD0jPRfCnP8La9lCP9VwOisxp
0pDWemV2EFKLSs1bTBtJR2t+sGqrKPY9TaU7AnrUMtqJjya2T2neWGkb4yxMD1jhliTnONZna0rV
jeWZqn8UdqGVsgmMyEQOu46SqId3S8nUdWHhFmmXgz3NykZXhHF/pLHs/6y1fkfTcC7TBc0VjJG1
irX/jQ8GviA2Z9YxYPXw5/B6vzorNm2xgWDU9jkx8CXx033PMTMCQLZErK+Tywo5aOvLNG6ux0R4
S5CtHiJsIKIFOg0FkR3zcmcuFlrITyQufLjGi2D0fF5vFjhQf9cik/nmr0kTjZ+tTd2TrS+5ZMQi
LtHyKtDX2DNGS6k+VpydENeE0Asv3hv18tcKbZbTwPSSa88aqob4ZcT+mC1PzRTosfzAuEowTjXt
m2swTFEORlXHQFIpQ0bDaOJNHn8ih8ByGJZVwDe07Adj9O6+7D8JoEPAfjkVJfYHdpairb96pcUn
iAaxYaeYnC+34FT/b2kpr0NDc2pUCpP/d2t87/GuqI9+VLBzyQ8SaGHIMQbD04ytQduFsfOJ3XPg
MrjNjapcn9htHXAoKZdP9UhT3Ycbp4ilkjHXCyznuOUqZ/FNSKpBQppbk/8MM5nBuXuJzYhLliL9
TT+jmviGWNgMqje2A5rjYCRQdQ7vzlaXOCrJkBHxgU6puJKbUWdECMAc7A7ZQtOC0kxN5uFr5Eyu
R/AyND3rFJop7xMi/CJjq5k0x4ssrGAbuR7pUYUas3UizV3ITuCRexxd7DbGqpSY45du7AJxkh3w
0jFItePOtjBXEnEpSvbTmCqC514ZBuLkrSEpAC38udHI+nQ5HTuUp2p5HV2QDqP85aAcYsCcaf80
456oQEVP/POuUjnHZ9xvILw5Efxg+eXi6raoZxxBhbaO4YzZBuUlrzK0S7doPEmiWYYcLQCAlwpV
lk1mP8WFve0luUGA6Cf2dmErMwMestU4i9RWrFND9V0E5jqIIrX/QCaebW0OH3nfzMqSbtzGsR4P
4jEZRzUCgiujpWFcRlojKv1/XbXqOZRAoYyuafPUCHCLS/GydINLHO+Q3lo7rmO6sxuxMS2nzn/N
UCjX3KgKO0+JpdilNEvY4FSQibcp5EJZnQ1lZ5rPh5krsXfaD0SoTk+DyP8J8yH8+H8w8a8Ppvb/
Jjlb7xNIM/zW0+iTj1Qdbt3KWt8BOD8uNEr1/y2T/eG2AEoUQq/qqhl22ewn/+CnoOozdCxwcn7o
XKPfuH1EuMCeZqDzEzYAcqrDldjOTdSlHrZOekPAn+fKGkvo9y+vdvoT4RMYFW37l6GdD3HAaHfq
oerA0fMeIZ+C4NABx8nIG8KGUd+AL39957Im5NoGP+weI7zUYKRFbHOwmGWq6EvGR1seigqe119t
oUfpngoBvObxL8a5SO+/Q1fKnJa0/j08UzU8I817/zdCMRQutUmx1pOs16Lw1thkspI8oCFTCagC
mzqkKGcHBZZ5/4p/bBEvvRJhb5ogd2y3Xp+lBAjQkw0AdPr1eXESFOB0H8OEG+kErbZKp8NjnIIj
jqmNjOhF/nti46IYvTpPgOHj9z51nXgGXHNWasiiqfvl9o8Kt+vZ18Yn34Ym+zdNvMAFYlsX1YEg
ZWaHJ+8eAxYaHc0RwnXgcj5CmcVVTUxntIG/UZ3hicZ+HBubOsUpzmjbl4e/xDPANiCw6RH1gp6U
g08beiHViXITh90EnphDnkWaUgxzMEx8dlb2i48TMH7IURsd3YTuSyktbzhoXfQxYBylGdejXNUq
bCesaboufcyqHAK7Nrchwsr3OcDzWwdLmUoZlbNQNu/34odaVXpx4g/nx3SPJinCECf2Ndy9Kshx
pP5UWJdfPobR8pP3KN5fggM036PhaO2QVnhy/xvTSP0+VAKtME4YxgAUs/GNueiNBqPSjWbKyUtz
BJtA3EenBUxP2w7PlNL+P0zhWejgZwRv9FvBEORaCTwCIMjMkRBd0l1UFJZlOOfZThb7KIVGflIn
s/OpB3Lq8F0d3zYJ3828AE5AI/x9lAv/bx/RHdKs6cMuELuYzrKlyJUzE8UKfPTVZTTk04Q6rN0S
VytVti64ge3eNt4Nh7E31HU+tNpPvWwj5jCaZxQwzWyuaA9APEzeO+U3k82ktsDNKtpBC1HBrTU5
x52jLfBhn6zbjlJMwxVfz1ZCwpX8nqtLHSQSjGcI9B6SN1etbQ7z06TJrKHuBbLs4khkPnDEpDnw
mCti3aLYmFtxomgZeCF+rxilOlt9BeSzaleBG6dGktsl3MyesZIjt9Qaut+MuePkcZdt7cNKj6CP
+3Yh1OJMCr8tRIoC8AAq+XLJm0h3x0iELgLJJphhiZ6QoLu7xo8I5/e/WvyUAxunr9fYWt98JBGt
1ShhCEIOOTA1O3kvqQbk2HXKCBrNuu41U7FGvBhaq+UIAK8SlXE0o+fkGPk2zTakO0DDKguXZEx1
CmydJ9qxvjggU1yLP3bhjDuZFMzehm0eZ9mkHSzngT3imp8A5d+u6o3QQl9L8ioKmn92fZCrE7WE
FRYNZDhE99ZhHih4h+uBd8baVQKB7pGu7wMAyxMQ36nex+gDurrknp7Z+UJrEVqjlnS9UfMp9XLh
YMrx1dUIqx5jndRfhTPyDqfoQl3vtYAKm8zHXeMKQGiBGGnmu4HY0v04XkjXK2CFbMgX8Esz+x7e
hK1Kzg0T+SVfbDmqwNkmMmyo7RqiHyx1CjabhYEeLdK4P8vlw7v73ji34SU2JYBd9Z+Gy3/hdFw4
XtvIB4ToFVfhVeJu9TNU4Ct+dXwyn2ZI5Y2KEweHDKip/9fvjI4ei9GMhrx5YjRjkjlMIJQtQqZ8
GVe4ZehkmZ6F1ceaaMb/JliPeDQ6Zf4FyOuwRBNSb4VVjsDbVXpES7sYxzbhJ85hP8MrhGzxcrCr
72VKB4pg15xRr01apEydcl8VFxXSTsJTBe/Qc0il4JP3QsyW7FZ+0sgiAroqyrI2sgoxf4g+3Z5u
nZ0ZmeQ4Tejir31DUaGhgTtonQp3DbqAEKcM9NOXPIt3HYh9nQDt5lWgl4IJNtaNQjmseSjQkBQB
0LzWdrNgKphGk4j+x7uUbhYb3H7H390ryD2IAWAXe+NmOjqppETwr78+bTSHjgwjvzWTH3VHcF75
uEv4IGgcnfiIDiBFFSP4m8ehiHmpR2e+3nJWYneBpeadzoQQu7FwkQkjTAFBFTokRvs46NVOMqbP
IQl206qQQsvyWzfmrYuc4vBspRoTz51eKA2tKtmUuY1Z0r2stJaFfVIWQnFbkFh2rrYe88opmZqs
BCv5oS2H482ssmDi/CJgYk38GeBilDFTAkSdjdgwJ5eKjjYRN1sbU9LxW1S/Y6mJNURIk1MI6lAh
8YOXLOH3WhJnes3YyHfl+aF1fZA+JDnzZHdiIxcunPQOwX56vJ0mM3hgLooNJYXRcH0c5p1cgCo7
1LTh3JY9uVXjIgvpoLqc0zH+HFTPcEz4D/cK5fqGDxUr7RR5HZQYYxqZkjR/pmbPbxgDRruGIOno
euDvMJUzQq6LgGwQwI7DOFThW9i2ONDZLtUD9H/aKyXIT+8HxJmgYHvcTINZD4qAnP+s8h6syc+s
A5MpqqPDaOAo5O0OKOOQxahwdRj1gcVxLviyIpGEz99CgBsZOJVICjBm4HlOe3eMtCGob9fiP//9
xQ+OHxFbLgcmUHKVf/av5JXwpMh/OOytb3NZEQs86xm0tUaRFy/N1m6NmywHwZ3ZBtgeQsP3m6jl
9vw2Pv7Vc32uMqp3Fzwtu/1jjHFBelX/OXZHhmlviGqw3DmRStzkNwry9RkOuXao6YFIRciQ7n3z
pyUcnCqDJJQ3zajARB+sjPL+uyOjVkuGW6sLHM1Fmmd2RNNpXSKqR58vpQeGnof2ehn82rQK1SaD
QNfnTSeMLOQIKZBy8IHo8/0KS+dTArwRENmDt/LSjRaMrsy3h7W+TflwIvLrT36mUdDEePNqYCKP
EbRTXEWaWJU3lQaozhm0HdrIZ7dq/dH1GRNY5Fa9EuAvG9uAQbd3ht66w6bkUbCB5tkJP7CSCAp9
FKWu9vcu1S98s1nNOyODQnKqD0Ar4bA2s36jrtxzbOG7jKRAFOnZbp++jq45rTWDbJJfOCj17e/H
K44qXgm2AJQM4SQhGGimNMonjrfXb+2fiYKpUtGlfMiSMQgHMI6PJykFinP9EPK2OiSXo+Rw/v7B
R4MlrJl6Z97oVOEj8j1khaYOlOtWvdnTnK0kZ4yUQ76UG0BHoV3RqosFoiEnbvygw4Ig2zQMeV8H
QxtkDfMlP7cIWoKulu/BV6DdccVUhXCibrtSIwNMj7Z+f7KYhvJ7YqwvNK2AwhrBRfyW2IpAwh0r
WeuSUsIwoEox9g0YSvPKS2E2WQOCJ3ZNeau4wDdnvgqDlA1znoXPy44N1Q3ZOL7fJzXbOZcFNjdh
KUoyhIM09r2kDV2qk1OJ/KPXeW1c6OiYc2yRVorHQ5AjmH+LB5X7MkxwYwq83aLxdqGfx7ELWMX3
Spl4neB5ZYzgq24ewI55xTCOvmfUa2Rk3PDimXqNPJJ2ngaPGTapwlQlc5wicljWMFkZGZ2X1pev
4OIJn43cxj2/6ViynbCyz5dCNK0qI0jFFqVKrpd803cKYjF9p7U/F3zJwWsXSOOttHhJQYW118wK
H6aJXXRFidoi42h5dtEq4n1l3HPs6qVmujZ1i0+3jGRkTzwfwvNdhLB9nZ6i7uzWZIy485tkifbN
3lo1yXjWeuTcfO+0qKWaDupc9cz1LDpsyGONZa1ssMeZhLnAhQfBKaUqSXTJq0ELKy3hyol4YTKY
+98aNbON2YbscOMo8CO96Q/pNRxm3ktz0hkwH5ZdsHunYVr8HYj0fE6CVOund5/N8lHqd0HoGcfo
VkcKiXusdsRzcpcQQIo6rJGS5wVgD5t+jEq5q+jXhAar85hHGlBzC7XOPrSnUctEUcH62QoI5mIm
ClUquzyycn5IYJtu+3W/edtY2PmIyv9F0SFy9weNqYOt7OXs0A+YcbTABBdEpwk1cNwtBGJuqmtJ
J5LL5T+GKcpvB1m1zVLblyXfcW7mZHReS4HQWRer5Yy7VYQh6fnj+e4zcqqiPefsC5vINzpKxNso
mCJ4oppcvkMF7fVRqWEAF8pL6n3ucqcak1+J8lfmRH+45JdOuVRZT5PEIUoETetQeAuv4ACYs22A
Sft2wlm3R4TPVmSUnk9Ascp+3QBH6Gapy6QtWM7PfR5Bxr0A0+meR9+ecn3rG0GQbpZZhkmqE8d5
fUa4e/SI/Xk6xbc27hWqfzRcR6l2VpMDBLansP4Mk9QehUlR2qMhQ94qUcORADyIYRX1qBZyXl9S
53SzVpwkfdPZda5nxGFUSwr5/TKTAMTw95XxYMdHij/jQT4D4RrGeWU5lULZrP50NOuWK6aWneL3
Du1gKA3pPeQmF315Sh8a6woLHGNPnRseZ35qe+elUcD5WJq7B0fqSz9tnaGRRZsFomgW32+EfNjX
O9aIYhZk+2NK8K4X8QaIs3rbh9ZxtkLeRBtclJySfSLpnAx98d9OEK00orobnC4ZJLbGYLRmSOYE
S7IsPa09F1Go1z9uP//aWlOayOaSYBzBjUgDObIH7U/sCgwmQzoGZqzhelAAIdQVF8DlX2UmIhel
63R+JODvPi8ADPLge9yVBI6qxdETWbjGM9lN9yUe69UH07bX8Xpqekzwu7tZpMPCp6tks4qaVchr
3fHE6yO2HkgobnJoMWBo5Syu3FkPhl8teTKSw+Q+U5IJ7aC/M/lfbxrqmm4DQW6SXjyrkT02cXq9
I2OZrjRvV+1c3A1A53GjOzczJ7wu4OU5aLXeA5sLqpcKtSJedgyGHd+txE4IRxmzs4bFDMJWPjxx
pM2RSIWKueNP2PeqWaa+J1YbDiI3jJ1lSx7iUp5xuKCSNiO3TFN3QXGUggYioeKiuDkxsIYnL6j/
dka1zRxTDJLNuIf80mP5i0+KAavZo8cDhmsJ7FZWkoiLveI/YYlf8x/7qObJAw83K2gAE4LyMLNW
D9nnh+rUMN+5V0V6oxoIifElvRsK+wimy3UkXo2IuUwvNLAvIh15GvpLf/uqQu8tIftC/A0LtiNc
CIzUESNBBsr3m1sIyk6O1stYs2zDrkchzlNu7gpiFx3btH9WkASHs98vG6YHoU8tCFDeaTTP/zu2
gJfvfKVlYhmDEi1zVDBLagnGGo5lJh6HDX/ThAUdqITAcKMxbh6DOfCx6SLx6gv+mqiK/U4GU+Il
nIT4KwPQS4twGvc+yzBOM3H9451F7c19lYpW6cUreWRl0ATZHnCN6c9LEJGk+qkPLNqv8Bc+PeNk
PBd2CwYOb4KcyJ9U2k2TI4VPvq+HbyEMUCgpNRa4GGpRl4rfhC7fqPBp4KpDWCTIgORE4hCSn1eE
KDX8rFF+sjHJQR+X+rx0E1dld9ZF0Il5kvnu9mMW83hjyex1jTSQbXBghl+S2DVE+8ccQf+IzLK9
+/k514A2atK7UP8y4uZT8hCCD5nlnMIpYLKzeV/6D+catI/MrkjYaws/XqJNTp6p8oqTYbVMkORo
gApmIUiT/ldHjaiuetvVgMz/CTmf9vllJidOYPEt+RuFO/AQ8epWkEj3S3TSBfry79CuptzugEvz
FyTzA61DWGFhjlilLnkSF/ZYstKXD20RZgSk9tX7EgGDiEvXFaDYEVbqP/4iCA8UyJZIIPNDnDrV
e5sqdZejoBZwmBAXU0sAsoKmsc7s/ykkt0ZupGpoU0woM09lmyd/yLf1T2uvSd0yNYP1zegZ8u3K
XSMCfYdkRnrgtT2GCNSEGiOiW6yzXzdgb/r8yG9VsuWMQqxCgkmuazlXX7itnlEJi3QIL+q9tMxI
Fz3YTDicubHOeUQNcVpn7wFP8cQKtSX5fCHcXCTiFc4SKGKVBwxmU1E5MCDQ5w1eiV3mWjszXQRv
5AVZSTUrqOlW2R6x2HAe20oXRMRj1CKP1UN0ypqwSVIM3ZUEC5ZzgImfoRivLxQn9F3xBZ1a24XW
arU/xgnU4FvFn/oNVk6F+YAADChFQWVBa60QcEz7p+VdCcWFki7/VA7g9JDiBngnHCJlYkzHZ325
Rh/brkhHA9LJmP7vOBiwkUlmmNaAb8/LpTbtDG/jIGQPsj22hT2O5RPSmg7Lu6BLfnps4B0OC6+1
7zIv6Ydlsc6U+F86R0WCPR16h+SEHLsp2AuEHW3FDZSUqD874i5afmo5BPK/gTOJteesILOqcWs5
+BYyfLIQLApUi1fzTTHaIhwlYeIOrT1gEUA+7TQF4MRMG+LOlPux/2I9jCVwaywKfMRD7o5PBa7o
M1rbBee1P/Dk25H7QB3mCeMzkH5YUhd0Zyt9829HNe2+z35nVuekspM4FyUwz9TjMgX/srudTbZn
E+VuvhzIM/EXGkXB1X/HlUFCptzoESOL35bF588Evw4HDskVxaUR2D3/zIl4+A9QLhG3qsYH/Jka
yb4t2OYvzjXYJ9m2FxkQ0qdPLXO2cFE3xS0c9C4YC2Xmwb/++QDVp3PYQs9Q3yWr3A6Ap24nbBZv
9ZfuxfxhRYWmVCE2YdDIN1UHNMkghyRNaNMcSJx0VUNer5dq2Ix3Cg1EdsPrkz/n0zc8rSs0tA5x
5UzedCAsOtgkdCsepRLb4T/8cC3BRJyx9HBaAPrxrWIz6jFcVXg7twJCGhwJSrcOnCWqaDcFnIfa
olrmumftoWx4OlnPiQmJv3ANe37Lqgysg4Au+ND+fuKRGPrSoaV1j5G1LCtDrm/uy0I6tkuXHyo5
etI3iJNukm4wRRhK8WUhmCEAtdITTo5BSmjxammz7UrHvY7HfTMuQfrlii1D32mNeomu9d/SG+/w
Fha3uDkqtIZbt0ZYt5hVcikTIhC22aq7OwrCnQLO0N+XrLtbqEVOA/JbWUr6V3A/rI8qacYn8aaQ
F3Uv/fHMVKmu4Pud4+PIY/7FIzhuf340ETiVAnqtlE+Abc8T1SHckH0BTaueG0jfgoGbWDMCMmBW
bZxxLo5B2ppGN0aLInzmM1Mz8J/CfGgVH21Ll2bZQLYRd/UdjiISM8XfasqhfnDV5vf3N6zqvxZr
mQYzD8c8zGce2lxXxALOpKpuuMgeQs2TLk9nUgzOQ+aBu73f9QrvpmQ/txVeRIRhJvcNpiJ9qlsy
dBJKeh32Q63oLhvMuCYz5iGxwucJrgPpwrf7A6mcWTF6bBT617uErgrO0w/ZZU4L8Z1Op59AxLeL
SmSPVxk+7HWqOO7t5hY72Gx6QuhsFy2W9ux+oSVsTuymJGxGxW+SZuY33enNQI8e6paD2ZPU9emO
q2dlBVLO2qIxr215+9OsULpSHA3xKzJq4iFqFU+q2kyua1cAgbQOlUxKdrp70FznPJGQO8ssaNzJ
iqMjo+J+ecJwOdCTRBofUhw8uMNr0c2WsWA63EF1TBH0deWdqePfxLQsN+OFFHILP7p0iQYHQkb5
TznrSVXJ4FoTIicgpqFStO1nfQLp6PtZ5AeYM/jkn9zMNdL5VwcHP3HURZKYfr1Ocp7rUlRB+xXJ
CdHdtP9pT/9y8FppoZ9lZrc7SE3AtepgExgBlB4iHPgmcAdEaYmKu4EjfnzS8Y5WiQ58jdUUwZsu
yWGLL/aTkGCP+FGam1PbgkiPnhQ0Nl3UfqdmSqXFINZBfIVzF0gOWmiepFa4WtpHzOvMBhkV9S+K
TZCXbXrIV2XvWFFLzhw/R1sDBUkNfYb5liFyH69qq7AJLJ7/XCReAtR7GsQHRY0DTP3ys+A78jtn
DRP3rk4KT/CQid0OjMthk7JbL6ekNPDm5wtnisnMHGp97nc5nmA5VmxPf0t4mvbnaFD4auzyzgcF
6rm2fMNPOiQLUz2QJE4dRBUDuYqRFoUES0OaQlRnaO5g9Eq15CjrAKhJjbsW+eyMYHDM0VKme6Hu
lXIsNhjTiMjDUwnKUpa0IOaAiyhUwdS3vgk73WpTzvLFQZn2mdmeBN9bycMPr4sYmlorv4ejj/y0
pBmdt87AMNADDBS3ssNRm0w+D4k6USUuZAqfhpm5hvmM1w0b9mRW6B48SggSHCtdiAJTji9ZhrGv
f72HX3kiV5lHqVTcxw7h1LnFZumeavSgCRQMyOBT1Ee+yuRDnjPtvFm9uaUWizu+KuWfAMyaibAF
5J7ugDn/odQRsDWFnLEN3IY8/rFmfCs7GRJkcVmQaVWui0A1WEJmNOj92eOuxi8L8d3uJvx5ze2z
IDoZYlk+LTx09BGT8aRs4XHnoHHDpx20VpYb63vZld3FaoXSFK3pD0JVf2WXVTZjnAbiBb8e9mhC
+XxebTou60wY16tJKBb7HKFvig4gzwEvGiv1JU61z815vXujla+3eeeuJWHlOKdFK6q3XkJ31n7W
3Jl+Uvqdspq2u+y3vAE5So4chnWZZE7kMIQvG+3jtvUjS/BU3pJSXVB3HlIbmNRD9A4CO0mtundD
8FrteHXkAgt5o0VJ0Mry5JGWB25CD5cqnBLr7NmeGxSo/vt64vhxDOi3dIRmqR7VsbbQhoFQAnmZ
opAbhAubZmr7WHg6M5pJm1R+moemd3jR44ucdS6BCaId3C8EoLjAbXDJh3U16FhABwIYR59ZDoBQ
CElWCLj2wlBN1niNLytgi4GZv925oRNtkiGOT9xF1ABafRfrGxDY7w8D+P9hBoinuoEEJ4PBXnqL
rMQ8HWVeaMvZRcmsrCvlmbxgTaFtEeZXAQk9aU33E51qakEukBukFFdNwvJbQLjR8V5IZnF8meq6
fAtDNvl0fOZQLjMrZdHgKTlpvZruirRNlN2z/cuHPVTk3dffovUVUBDDzWlfkExWfF2kTN7zU29h
EIrH4NFqiRRoo60imYuOJkvT/mVn96ZNyMWZ0IJd2V1PKhWtwxmgRhHzFVZo9OypVR6YJxTzYx9i
h2kN1RGATwXM6FUDG1sWXyldCn6uN/b+10V6Fmi61niaiXnZHwf6Zn354NmOVbYUaCvSAa+/IYCe
0HPX46HBEK8mqS3rtZIUO43c63mYKHBwUrC88Pk1+ViIbNwj54dSgz9RqT4ZKHgrNbs4xH8uPQZX
qdfNoM0YWh+MDg2uQH/G03DMD54A1GpGvG6CRvfxf+n2SpWAT8dEq7te94SC1RpubbvqPJN5ZYEz
JeWlqM4ABtIp4/oepLaQyTZbPa7M41EUzfwa8YzK8/IT7TF8F8xKn25PmmbxSg1i/TscVGe5o5p5
a+Odek1+WwGVql1l4mzSJGsy2cs7qjxm5g/6VNorXGuB6qA7u0G5l3j08S/cS4QUxPNRbexDcdrI
PKNkIaKQOosobJTzMBBAKKbas8j62abEvdPWWtx2yEmFrBkOFdnE30NIiLEVXgnhff1k4HlFgRp8
gyQd/MRVMWYGootUnfbkB6QctpuEz2paX7JZqtCbZskUH4tbqTfspQvi/Q98+WcTWj/MBmukIKlw
ttOOs/68mAFwdLSpmtT/+W7FzA9bhhKNBOe0KpPXMSddG91i51dBIo07aLThSDMp18GDCj9cMCKE
pezD0VRFosc70fHkvGoCpp8OeX4/me3Lsz9FiWQgWvzxLs1xrraHGjN59Q9vLyBg2fzmu5GhfGgE
HEdrMYNwc7rX48SSKrCuOu17iA8QTnk5POiGaaX3rozMsj110mElS74cqAa3OxucXmycpalE/h77
DoFMOIZL7QXpnYz4CASs+LJPKIsbkPgmGtPzvLQjyNC5hprENf44+2czxrtuORz0zUlJZn7SOpIl
/yvPcmM+SKJUQLjU6SjbTcV9h0V08C3kn7KkFOQurNdBPPAzVL2gu6KtCJj4qFezZ38a6lv/4FJQ
0pCWgqhjBDqaLeiS/e0g7cU76H9WJ7HkoVXk6m6jVlfWOZTL3E8pH1EU0+CnIhSI/4lsUz6U2O3N
+x6r7ia2yccvY0/YQsuoLzdTllprTi9oAfWqp69IGKNZ5Hq2x8E+qYO3BnEwenx8BtPrV7jlHFJl
qDYvckxf5OEM8obctMKQmZako+/ml0liiHaxquPVYUR0Jpzf3LYvWgzyq9Fa4+bxpIDBp6VY1X9y
Vk+r5pHf27g4+lRRkKNgamj84TEK9HUxc/+FazGW6hsBIoqq0caKlXjiivpAP4qCxDqnhWODTB0K
o2TbjryecsKI8OrDwLINr772DhvMyi6Jc+TmOJ7M8iS52gzRS73rR/LlrkPF+dxTlAJvlvIZqfJ1
2Zk/NVW8s5f16KVlrqodwRIWfKNhWzylDWxccDVT92s47LevwxKJA0fW+C5UaZSAwdh8obuRiqET
W2+y4LR8I+bXI7AgZ+3+QpbRQTjyVr5ti+q+Gw04qRfzOXKm8BOZi5WzPIxL7b5qLUoYF3GlQYuk
hvfcwBONOmhOYCNIgbTPW1is6Zn/8nEiXAk8pPYtTwqyb4biNE3Itng9k75nDu5RllrTimI/F6nZ
BYTJ6tj4hcLOgGhobJ4yWzG8I2D5LIUtf3nd7gpIIN5vUWQzjMVHP56W9eAWWUYBJN0WQz6bvILg
nrvTYcMi+KUOf8/qm7C0CJdkPQCBy9eoRp7GmQcXpQ2LO8Y4DYUvoqkHdDLVEB6yzJWKMQn8uRcI
38gp9L7zqcNLbZU6hrOmfKFyO97bOx/r6VF11ybEF9w6K/76PB9hu/nYY9RPBYFBl3a2pPyg3GYQ
g6kCyY3DbdQk0n9CimULGuK1SU/1jckoWxbpPRPyT8LukmLFwd6pDKf59n3sHAaJGnNSbxWUbLaV
TYjpXPQkdaGaxCwrgb5S6mEEN/AeMTwM05mu7hQwMz7eqIbh4FLLJy1XlifKsxKUuZUDr5RWvnMy
nDQRWA6D13Jh8assJgBxGi5v8v03n1iMxwuT+p1TcbYVw1to7VdqgJs7FfZXxodyodA8ziXo7MQ7
z+jdGqUl72AyPoqg8v3LDXWjtHFQf249yPLhBVMNyxfRZkHY6Izm17D0xnvJocggmajiW71ufqTU
NfjCAF8p1+/+nrXSUZom9gXF5VwPJppBgBOQVkbWI84Z7UHF6SjzkK0wF8bGph8l80170H/WF9OI
YVD+RiS0lhVtatMYAX+hSI1HM3Rb6PrnnoCR6vvneh1zXZLHaALlwilHkvA+oZEmxwczRMDTwJxO
5y6VhKq6q6Kf9+gMCVNnGgdW1mb2yR9ZRx6n9mHskvyapJbkyYbWJbRyQqVRNXB27g39+c29BR8Z
JozJbhCMi8u2KZKRRe3vYZNij8whGUObownNeIz+y9KOu0x0FhL2AoczJEkgsKjQwojovrLtmScc
GjGG3SDil4s5T0Ou/Ht/+Z0gpAjNjEFJUlY+60th5fFOYP2mWshYP4H/Cnd0+JDuXM8hAVktpsJo
gd2gVoCManS9nPftJUvWUdQ8Eq0xdPOiCeTkohs7NbXejwrN673WqKsrHiJFoN22aiDY6qxP08fn
0PU0vtanbivQ4Dx/e6a1u5ZmcNY+tqBMFBVCDUyCOMfCzlABKvrC9RultsWh52pZC6K5Xs6LeGM2
XCNMZH0MB70SkwY/PqoSi0WTt1VntApKF80x3MgjD6CdfMUN7tGgja7hCanuzcNxYX3hZIc1BxNt
dIZXQYow72vAR1ftyx5g/XJJZ4XKXGHQWvNTK7t0zPaZhSEt3B7uuYmQY3W8FOB5wX7pqGu9Z9cz
JWHj7nutY0jlvAjFlakSoEhAWrGA/0jjVlIm67SPCYh7hdeHkVW/OpIGdKlblno+YldJ7ObeSUZE
BYcxNphN7gsusaUuwpFlHsb/cfQKczIrvPzMCuGGoSsxmxwQkQIIZQ5IVi6TZEwLQ3ZaqgaWuLjb
Giql6ISXK7Mz5gD8uzuO/U4q9MPnfjjspvuwPXE8yJhCSKLgXwpJ+ai7AByv7Ewe+aVVZNIWHz84
at/N/90Js/TmWLrVTsjjXq+IHZL1RnbXJbAEFDb+ksVhFn6++DD6qL7A2QwhI0ELk45P/hSsIJo+
Zy0RHHl9Ju77Re5IjsdZuZ2No8W7tQk7lAhoxwmeyOwVD4LTihURbhkuM+vq6P7C/00CKUZmxX7B
XISWS81Bn/SErJf4B3EzMLVALdSdzvq5xYRX+N4nrlYefimMGMQRdFY24rtpMm0TBb8M25LsT+Zk
ZFspN1f5c9mtQkubRg5kYv7hkXXEQJeQ1zIRnxQI2mcTJ0kE5GOGALWAhAJfeOyvuI1fnpAagXu5
XC7K5QNlp31BUJmjtUDlJ3PZ0dhp2tKUm05mh1D63OJMrRB2IDLMJMkeZka58bVNacw6FcQ0xiXz
agjIkF48niPvisiemKeKdsEVZ/bq00d6oJ00rr6WQdecBs0ISmkuyrJE2W5i53kdXbsxT/wUNFzH
LEYTHrKRfAZ6IVWnmqvQWUjfbrJ9EeS4/Cv8tHf/WguhIZJme/Uu9HR4R58eSXKOdZe4Zf2n7iho
GPcuFlnnsObpNOv4hCvrm4QjiqO4cG8HjchPZF27Ip8kZm/m4fufiyeI39u7P67f/kMIAZ9sHUhW
VsHQHxf5Asm51n0x1kFbpuGMfAgJZFhrQAJj0keUvLtonWPfCa0gf1ELP/E+fFAPDeJ1aAxw6nND
CnxenxmBwxw/EFdcqVMmHJic4JUFokEXCTvH1RSoqPOBrhBSYZK7b3MVfrpAddVh7IC9ndeUmuSo
XVGirxtpUVDQ+CwLVPliKrCUFItgaxEsc2S5OE4Yj0n3huJgy2vmbwyb+AczvBfNBc5EAc3Od/r7
3rP9dLeCSxtyGFJxhBKRjzZ4O0UmyHCrspPKAgU2cFqSOVzfR3GBM0GEhReU6MRkmTexilK1zdGO
74uaJ5ImmBMjmuQdcZ39p7Ehhg4uTDJVsvaBG3jO7iCuUARJTWYiecMzCrSEDdJHbGavujNwZpDP
bFTpuuc+Tv7HEK296br6t12lmholk+GFucnDvVe+PGILux/FC1Lm6bzX66fTOejFARlSaWiBoLZj
KcV7EqZEPrTiY0CfzKxS4sgCMiqTYqJOl9V5Pr0ntZ+wP+BQcICd7stNFo0yA5CzNSTMvE275ZAf
C5/C+4/4ahOOIymVSutqrQauQTmwvj5pfRaX7piOqiWqIJIVO6+s1qLsXwKHiT1CWsu9BMkwFh3e
3hAfCBHsEfyNLzrnAPVxuJtvSaSiMD6Jy5PWI6NvyPayWpXkNtcyB4EkI+BxNqXykwP/jOHckoQ3
HfniAEqR4EOgS7UHRpsrgL0puwi0EXAv6LIGXmxqN4EAafuJfOp/+MICK+nyGIUSuzZuXC4i+WWT
WzDhmOtcPKKZYTGN0YXxkRy060s/U9iDTFpmRmeiSJyaZV1lFUGCrBRF5lCC34MmJ3wcuXiYvmUp
6oHv4LrOodXCAAW3vc6GONTGBGrXYOO3QcyBsbygEkcMlrakwiKZVJDHBYKnkBNevvB31eGlRt8u
T0n3ey9dW8u18q+ja740PCqp6/n3PMQpalOvSseDj9ImZoEizZKZuGDPCZC3Vj/5ZI/dvHs6zXB9
mBhSiPyX1RrWBAF1K0q095WMLqUqU7Sr7A76vIPQBx7gz1w+vZpv7rXCs0Ryi28ia2JFeWvrN+bc
j9BzN8bAl80b+xKk4SKTgb0BJOvhP2O9FQbBgtlyhio/8+fed9pcHbJlH9VAQ78kHb0iOdx7R7Yn
MnMk28k/2Ge6afk6OWbCY/8LldHfzmYdqYx+MLbvLuWHtQUd+8u1pOMaHIx0xLYyscUPycDppn6k
Xg4xQM1Go0hwUGrQA89F6LXCecip8BNIOrexJ81MBldUWwGmay/y5TWjUYNnJaoCmRimiPlExjwa
eqaers4FX7zZUySqi7I/IPQajK0gDCrIf9R6PXzBZbtverZf78ZQ7sViEWxLtQWXzarXfszvmhoK
Lyu5XvKLzlMqrH3GvyyrLW0LTs/oyPtTr2PocVGeMs7WNzA50PkDZmgp57O9dp/tM/8mVSE5LT0S
ICVqXAkQ6Cdqd1lQv9RwBtmfiECsgSOeDEhbBrynYCt1o3ZH70rEAAz3cVrar67xNACXVo3i6bVS
CqQJ7U0vc3AAaYq3juYYXk5bWwwGgi9mg0VqVnqaKm0WGipjMnpYzTABnARqfTup8NqNCgLVUZmj
9kzm//2sitWV5zhIHGH8IPfCtZh38cW5GvXOp5sOfaef3Agq9an2m9QMPwGo333cfyyRGtjrF1v/
nhMNTwK2M7javfx98Wm87epSd6xxTdiuNAiV65s+XYRveugJfOOG1WzFBcnJIE+CXi+VdLGm4z5r
Wkee2/v73B8ANaZIqoXqLN2IzlZoMIehfxaStpqtpbrh2JZjppVykKs1NPSZR+epDLFylkBHyGsz
4vE6bVOHcWORDajZ6CVDhYfCInn5wmIwYkOtPmsBOxaVPHKaRjQerSJx4yAsueYAoM75+k+omWoD
tWgdrY/repuOvcH4Y1iQFVBSfDlmQRNq0Rcf0SfOnrp730+z8oK1oytHq3p9XY+IrIl+irHJzTKp
CzVEtaFHW/uqpDEeHcrFWq/zkUdEFkLZBjk62zsjBQTArOLr5NTpAN1NAEgplZI8i5B4HGV0CgtI
BtrCSMvDNskWjffn/87wXaqsaKeIJhEngzCq8go40Eo8gOXbHAjlnHiW6/Dk/cEJTf0tcjUJ4Pel
S8t/BPQG1faa+cx/mLx20DyGzzDbEJD6t3R0GdoZFFGzxfPMOsp+GPy8ZurJxMeUxIxTlj8yyLuS
iG9Z/0d6ixwA7/xLGxC4tSDf26JwBmaH6Ri/9MBED04+RPFOvL0duNgGURtnnh7Dwd4svWnYMaiH
vzBy+zNYQlFmSKNj0IFmR1X67VGEoScAIa86E/AaJQdzUacUI1QnaauSrFpzYjUsH41Qk8T3jVXK
qyKmzbPUyVKko7729THraKOhRDV1AhWYaxD/skmJHUx8XrXg/I44NEHjtO1ff+lPc/uXM8wgke37
Gel3PVUsQL5qi7bYu3laOydeKC/ZxsbdXodzcxgmlk+UVu2C5aYGJk+vZIuSVnwrVZS1f/3U5jMH
bvfJ5heGzFpK6UHXE9HPwbfFeHNNlVIrfGv2I7rvu4ms1N3gHNNDQtBMJn6CGjfCR0IejqRPsHWZ
S8qlXOWvRp0Qw1+Io6rgcsDyGs/AClNqsOcqT6vAMPjor0AUnI1szChCcbgO0vplCEuoDecW/gGE
yWwSfBGf3TF+GYlXp8BDFoYUGuDRGWwiqFTSakWqI9aMdUbb/evXc7Kf6upjI7OQWRvGAZNUevhE
l4Uhc9JncISHQcI4pS5Bk98PX+T66uD7Qjp3r35laIVmadRflPdhZbDr9jVPtFQvUrflrs7HsVnF
LQopfHGaUleYD9+aAw1Ptco0h4ARG1eTi3SyXi/fyAYlec3NAeY88HvsIP6BJbJEpaicYqmqROEO
h6EMndkq2ewt4qV3oeCeftZ4BSybQXJxPjUqVfbuI0qtZXYWfFWpNUwmlYk4HzWLjlu1A4/ueTBb
VgbBsSovgj8dfwPrMyzeWYcL9ElKEpkX3RlOUzLxm7DHCEKW5k+AdNzhunaBzCHPvwJrDJu80HKk
6xuXJGgcG0rvY/Nc89OoSA+m/zj9PN+1qxUAMTSS0bgFlasathLULvQACyuqT2tdn6+0R1dFzdBW
qi3yKPbkoRtBrMm4KWBPjFaSlc4w5GsD5SG8n1o6erI5Kvb72xZY3P6id4w9WLAfzLev3L7pgYg7
LM7bQrUVkR6qKEn/umF1iAmOVM368Cofk+woqHV9lo4P6Y5zvG2kct98ZbqEHtGhfpuLABQfBSDJ
gecRhptPo566elkzi7UnpKYL5SO6p3hLy2Hz98nKgDFnlrBijy5nmzavO1yW8nqmpb0wWiaxWN9E
oC2JVkZIa6zr0z5HQPqRdJTdULZ3y2qlssHgkyXKWiLM8gzstqMomhVcP2WzTvBHzQI0L6n/1DpW
H/VAyADo88aMujmyqsSjBSDKTCDshn2PUqED+HkHwBcRQz4W0oQ5OeCSZxPpcbHRw8uxnKmfTUV0
9XaJ6p0QJK44rE5bxlnoACEruROusCNArRxfmjQwOv9T5ICLUb9yQk2UMtfcJ9XCt7V8w/5qzOO/
B5zLEeRnEylhNS0fp6gfbJnNgbSssMtKhDM0u3r535MBqHF52vD0cohQCX9Zs7ZRl1wBXbx3YO3K
tsWq40F4JxtdoojqedGAOP+FQHbMLaJlZzFOea6+ONPUgcSw6CX2FFArP+T7LNE0aNBWk9JVJR0b
czYEZOPoyza+P1pjPdcpLrK+XzMfsmflwhwrSPJB1xsWkH1IF5834hjczxbpx9AhbeTakKNESyy/
q7SFYAGuMgL1O6mnIQp9LzWY8aJbtA/KM1N5p2h31uJlq0Nnyqvaw9Qc0PIinHxdTqnGWXTOGLlB
wQ1YUhelfo7Kc8v8POzanQJ4q0aXomt1i4/vwTr+GBaAVO25v74/792Ph9g2kYspn10vz7roML6x
d63tf/1ubQJkRa9KpCMVpBDpX7ZMben6WOIYMmCjN4E72NTPVMX3Z4pkmZwK4yoU0pWbe/Jc2UYr
NbBbmLYI9vM6xXjUiGqrZ6+puUqF6ClKcR6dVZYzYPq9+shD+msZG5GkTBUUqy2sWoY4qxoefgYE
hqZ6KnTVfUKTeEW/m/bir+QyYsPwpSD+/l7SXofMhm3dlENOH2MVdg9//lsaa2/JzjSmQhlD7jH3
cA8iRLEcyccQm9Gbo+IzLg/Cy1Zka/tendfRWqx9pM8XDHKEfCKFLT0uPqhl3X18Og42KIyUJZeJ
+uTHeXX6BIi3VTSfOxM9A5T3ZEQv/5xuyszaUWk7AX9f/7Ga9wxugboa0iv/ZUhihCv4Cbe3oX3J
jv2nfJMTq8rA+2EgPKD9Yjrq49XhKa5u6f2I7d4N88wzGx8OPq2BaIx58yW9lI0k/hGVw3K3+ols
CsxSLegxWT70wxPuQy9CWEmI1QmUrWzjH9pfoZQqZWTsLQKzoklxbQ432Bcw6PQs/7FuuJxL1085
1RkvnVVmZdjM2x0lTc6XxEhnJwPter2eYbvMI58zW9GgeUmFR+YAeSN5ls4uTKaz2Bkf6IJClIlK
VcgBEvywGXeDhuM3rZ5jAK3j8ci7Y8/powHs52/kiVd6Ijy+jkC7iX8vV+w6SmwIa3Play6UWi5c
2/g8TLjTF+qvs0oEIioVwyhiPc+rMatD2K1nl0S+RNNjXqWdZzu1uNoW7foN1QcUa2sCPDF2A2zF
e5WBlzyjejtGhL7DaTre7ubx+MjiftvYuR/OdGbWeBMX8PkKAC0jCHy/fKUWBxXrr/Rz9+UY+QXX
pMY/Lkr8bVgsLE1JrFV7psbeUFjMARAh/kjVMWwPW+AhqV4IVnXoLdNq1UwhZv+VN8/R8eAxeV25
pRAt5JHfwaLonZrC3YC4rdjjZnEKZlZl0oP6NKDs126dDgNxVES5EPa5PTTS2kwwT7Nqq994vlyC
8a/zV1IDwibNaF2xg4VzuT4S1n4TRBAxTqQQUt5a8blu1pE1KUCj2bcKIYhrdxxZ8Vo5fiq8TnyR
5AaXU6owKkTqafdV8J0qMbxXhfsmazGcxq7az+q0eJ6kSUVmFBbpTCB2OBAZlFNb1h8i+cdMkWVu
Tc6ppZh9+VeF8HwgKhudeLRvZEJMQiRxpHaa5FFiF/Lu6PAm3WE2Rjx+Hvs7ciua3O91yLkwdDSS
YU/vu3CjhVEfpXAkd7XqHsWXPmKco401kAdRLlEyKyYoicGpLB5gEXEwpPWLOE/Kvo4CPcBBrZ0G
mZWS33NpSFHhJmfu/d05qaYa9/jn/p9N6gXWmIom3pvgYEJkJaV4ZoONe8X5Gl/83yzQ+WGUoVgn
VUoY1HS8WFWpxHtLCAjGN8HoT890WLz0nQDKOEDIo2g4GssoaGGoVhmZAQtSVinF/AzdwIDFq5wk
uRiqOdbVolFE+tWJtJBLTFXQLFO23hiNdsB5S2N09ohfpnLXMgnN7oddq+eezWMTTponLWcBPp+T
ovPFBQm6XWwIGZLSishF/yqE6wenolqv9Gs/qNK8QLEdJw9pAAHu+9LYqnyGxVUQHLIk3gNqmt+o
f4kL7DFfDGh0fTTbezf+KY8UmBAUhsE7m03GSbUMDD91JggC70Sl+b6eaP9H7Wd2gfCzzJbkBCNj
ETMixGGahbZFsjyRjeQn5Ll/OoiYiWcEFM16ynNbTSt7Ho4dH3HJxQpASWAYkbTz+1s7T2Vw8NpI
Dtc50svvni97pNgAKB1KaNoaFHxEClUi994dyfNcYpgJDx0NG+HwHM+FcGNFf6HunHBhhnofCE/B
W8s07Pd8h+f/nvyHTC1mdUT89WQEM2H9WEKG69cUcOvP48yUAtOAJ5TagK6+X990bjLJhYbYQtDB
ySo+ww1+TGcnHRIscHrswuot8jAy3tNOavakrovxkzURHqDmfYlMKVRZN+P7YOr6dze7+LqnWqMy
r9PyfRP0xMfbpqWMTOht/V72tfcb9aZKSYgLTtVCKH8tyJHsiD3wvwQDZmMRGr/a3AeJKWfyBYkZ
+TrDGSnEwduKaonMOKBN6SAV5YihrWxd4bKDSLcLR61Xw6TX5vRKixHmwGiPrvrR/Ck3KjED9Fgj
vQXa18LSOOt5sAnf/3bZ99DzYAoGZs5msn11t1wgToZB1JngpEMxXlMY7AJVvFMxBdp7kk1O8EER
Jqy8LK0MXUvzbmYql002HdIGELKQp4b0Ejou4hsCQSudzJirxxeGHXGbHiqAj2Ebl7P5mRTc3p0C
i9cOKYiLg5cHuDlZhSbS6BeseuFjgbuSdyejkzlRd44K9xt3FX0Gpjx3w+4whJ0/pEvqXsnt5EkJ
2T77vjG+9HAp0hbDDkWgD6i28Bt4iJunqjuqt05YSdA40fkz8FEvSeSpLtDSbIFedA/lfDJ/1uyS
BEq7R0ABa0iMrodQ5Z/Q6pSu56Qc8pCFe3sRgrKIWsx+BPzN1JvtfyYYx16EOQGX6RNLBrXmE3IT
Y6Ner3tUSoo5nWEX+XH/BduDleYNiZDLhGQiJgxAbMkcb2qkr5N2CN3NX4Oh2/8f0RxsnNww8ND4
WEsx6/8EMFhLaiFlXcKkoy/p3ZWsFDJCWVfpRfk2xnh0LDd01a0aZ4AChGsf342lJFS0rHn9UEpc
PFd7QCoxgKyktm0HXmIAeRl4GWpHGGUlSMqha1QXtPhXw0tgE/+M9/pZtazN1WFsvbvG2HDoZucf
geposuYPX6Mxyrz+9AlxRVtn7mnNHgpzJvkgzC+94ZrWwAHL6V8+uTRRUd3DCtJMlvdHkLtHKUny
LrLLwdOYM6snizoj3fOfiATrKytazjbH6E3DxZ+r8JiSBZGLf9bLhWSF8C25stzpQ7QXzDaPypQ1
DKbZ6EZBBwfP/vRpJcMXmyo/OBdX+vxn/cLISluvZedyicNzyJa2/9hgO+QroMbBKlRHYaGf/nly
NnIw+IhpvHxS39+LSfIV3WSDy0s6HuQJP/SbP2dAMSmEZ1KoOD5LDVAoDL8uzTr6hQT3gdceG9kC
aIh7irlCA1K4SPKbd7TNtAa8IvVofq+rwqajfTfFTBdvrEdBrqfDwkGceFb0M9XvtTcNITus93DF
y3A6VNv+z8RkuGW2phX+mVIxRmMuaJppgiX65U1MHjdNHNXjU+S9pkd77c8P2VmsusK4DvhpcuSO
vq/+749pasuhAE1OYb135MsEpx9/QFAADVnAD+17o8hNMz/Fhlc5GFP9tQrsbhhnJ92Y31F4AUsc
V27IpSOXWmfPfXUQNovJytNg4WwDN+ic1kkeouvZHt/0QpiNkw+y4rwVk2io1+ZqHa42cow+Wunj
jQvoE34vV7VrFWW3KvYtfKx82/Ns4GrKKWZ6tzXyYCleivg8E3n8vugUewP4phzBu8Xyz4A1yTlI
JHPue9xeWNsGQe5giQozLxcYQ2Pz57fejD0ZRB5pS579g13nEUZjGb9mIYI2AFvh/qy2KozcOMh+
+wbmOgaZmCU2oFXbJc+cd6xPmh7DEV5tkwsDCHMqlUQV4ktKpF/j4boYV9uJZaJFSIEClmC02ALl
tI0Mmqyq2uKwBygHdhM8W086lNErz8Gc6QAnGAKBPVpb8MG3zgAIf9jP52S1nfXoR0kxEkuFiqlO
EVQhX3ETaG//phJEYkd15mpGmvYPbGKGdCuIrxQCCXNpCAjnF5B3bhdB8fTwl9lFAuw3fwgv1OOy
QrSg02A3hj1ZS27hGu2QP8Nri7GbRqaseyRMkoLqx6T/eArXMpdkxZYrFH7mGFJ8L5T95MyxYo4r
exk8YTtxpKF661vcCGzTdztjoF6B4e23ifAA6ijRfkt2vJgWXHVylsB6+yWffm4VbhCcI7WowvzH
NJ8VeZBFOdV7xscicuhqbKpg6vCb+0n6Ic0HRvXTdiUe20jef2OwtnDgPHP6b43hQzsJcFourWgX
fJz6Gz2+qkLvJ140Yp9bUwGjSmW0zgovogvWRdAEMnEcjgblEPvJmHIJhXHnq8AC0FdTQs0R4Z79
2xZSCOVp34dUKwqf1JPagDVxcv4bn1/18Ivgk5Op/ECi3t++vCUditWBkhCd7Mr8eCfO4pdgUquy
1/7vv0iFSTxgi1bI0M6pV4eH8JN5YHQMxWnmzSG0bNOs/lYywUe3OwdpM0o0dgGmcDrxZeIuQin/
9yNAuShOlg2XpLC4Gn1I2uLCfZ2xIh4/VEDAGQe3Zu4U5zHO8CKUHN4etgnV6p5wbW8XTXjqkM8V
3X6NHm143AfOggqtEhKpE/tKqXH3SzCQ+4u6B/9X922iXuMLkk1+g/teVkRhlJJYj9N7dJtj7BoF
t2pi7X4RxP2N+3Z0tfuhSwc9oqE7w8ZVzf9Hq3lrlxrhsE5mdH0g3br5lQtIrUYAzgcAjGohC+n4
DcOKjYQgNAEOo2jL6tIYR8cmadmNxXsgZn3MgPTEzeuAKrZuUexsTo4RjBCO652Bitk7g7X2SbIM
GBpHU3BHXy5Hho0/KN9AdrFfXbHbqzwX6TB8SZbHbKklh1sPKtKhTt73uDIpj2TfKYyMMcTjNiaP
EjP+DF+ZBmIIt9/DxaOPFAY+rizTrfL9L9a1cy38dMN/Y1YUwIBiHTCReWuMyaC1WzTnFlnGslYa
wDB5l3nAyLmT4Ieg6b0Bm1OSod0XpN5mPRz/9E8MJKyn8nIGPlVcfF373finbxan4m6rCnb7ZjW3
hVx3yiQY/QCwpl0SpDzrc2FSmBWQEHWGbFL47gXPoKtLbz/ZLOR7Z1bt1wOn3MwcBIM0RdPyFaLB
7rHp3O4wX6NtGmUcoQZdZjBjgZQue3lXoiM+8jJ1Fz20O+80OagnnHD6cZDLBVm5NNf5dA6YJBAl
GvClbgytfOklVwsDzwIlx0d6fm7ilYA9YQRJ13rV1nQynodYbbtyVE9UMHC10NSfVpXcGJp1mpO1
J9fByRNtiR/LA0hSh5bShCOM+HD/mkcLdfx1E/G5QlT+QY4ucJfq+2zq0s3DmBRanPgkmiHawOCd
YWbn/NXe2SQz1MwhjpVN4nwvjHKkhz6PwDD9HeYFj4GRp5CdTVJnVp7Mm1XmMfQA3OjE8hKam5z+
+TynGTnACLQmQwcWEViIH1uywOjg4IEAl+mAjkq3agg2/DsXf7CS+335rvqx0WhJB0f89/J2LkHi
CkG+/p11TqRyK/Lr1AEIJRSzwRPlGrhWrxl33ckhLCBTh8BYxITldVQmLt3cQ9QtsvL+lQScfBtq
doAMjNI0o56+PrQ6HXXYoB380k80KUJ3ojnDnJOacnUGgpTbxe552B7S9FXstCkpYDMDO20jOHq3
X38d2VD6RgqAR7/L1K9FFq+x2keiiiwej3VeXPVxY0GgmM1K2oL43u+SLdJ4xZ/Nl6D5WssZvftA
2ulQQ79tItXSIeTB2wM7arlCm9rhzKef13sOspBetQ6a6pByYcyEZYFbpZjWwmXyo5eZukyZGASF
c4Buby9mcdmrnGdaIogLhViVcHphYhEwRayz1CuufNs2q5DF1X2J/MBnVTT0o+lR0jrgyxiWcSTi
Lc2niW++am9j+ZyJr9JXVkRSx9unZJLbIimqSdoMNzHjxqHh+PtU3yalAXc9n8oU2Aguork19jxb
SAM9EqmBC9S/ORbTxoS/xNGMOgwzPjYIE57U/ZC8n08FrkxaFKJG/7smNNv98kMr07I3Q0hntXk2
Xz7BpKJKpJ62CuE2lytlLNQ4oYCTNejEpobOe+Cwzw/kH4Lb4Kv51SkJtieE7iFV+YnPd6TLdLep
WboecCloMOmEMwAELe+No9dMqyC6sGj5WYc1p1/DnLijSFRSUVsrvw6vH/Czhs0i8+wcnsBE4ZgS
hVGcA6E6BJXwfeBp0UDEIKEmEIPOsf1uxkNhMKJ46Tmivx99F0zaFQnKnBGww3jLv9xSR7OeoOk0
CzIAZOrW4qC99+wUH1LAiWF9D4dYUJzV096/ghIeidigFTZrLkJbj6d3Hm3SyAksmRnegEqT+7yH
4jI9qQq9A2GzKHDk2gqgLXf3Bmvm8G3FFqjkEbtXJIIhK8W8qm+gk+asIsb+B6GHjn6NS0hfvPWq
TEmoVPeAwF8iQ9EvBJ0xY7o5uFjcSlqazfIXTCXe4fog5hLo6+2ijzyIBCLKjIm/m5k9vkv5WLgd
Fdi1mIjZel/ZtESoUXr//x7hj6L3kqhHal6LfIioEZBsGlHf7vNiNs8xYgDrB1Jinkiwq/RdB3Hz
mLK3ccNANTTH4Z/bZ7SSLgDVEAPPPwhDNL1lBRta54McjaAz6JrLvSS/s2xBEw4Sx/qTBVl9fPml
KTkpO8zQbJBHeEdCyvTYE03LVEkSywM2Mxtsk6NIe1e1ZrXsMhb35SbbwiCVZp/Q4S3BV+GjkAHs
DKw83e4Qr4uYo2TOXscwI6m1hHdQKGmWjRZHuoeEx1ygqoPtgyP2PMl8TARTNNbqtBvdc5Dsew3h
NlUmfmE4T+4MStuI8C92CCbEBb7D4YiNAnCbjGUdo2WFTtVd2XPzFXjyRRi7kW9i8aZ8Ufbl/NS7
Do7MJ+oSzkkmlFeAVGwCsDbk1bmABvMBQ0+XwyrUG7cJhq6HMD4luD7KrCHncl65600SL6EvI0s8
l7zse1HLnrt16ZqNZ1ebIzlpMzn9HpU9RC38FomRlLmVVG77GvcFkG4SjqAMq+RXLwc8Lz28swpI
z5dp6fxLxw7LwOOSErHHMwEuyPDhrldMEubqIjiQvYStab7Wa+vrMqVC0fbh8nmZalSVGI6hqKP8
wyCmpYHl0w+NRX3hOHQMo8MdVVvwjCfjZO6E2qB21dlo7/LXZADpEGOjhhHH6f95ktxFr/m8TyeF
XNkPuoXdlnN630iIb8IPHklxlsORVa4GX/2liQrw8Kiq8sEqSbco3RcY68Dt7HGNbqkNK57uG7wm
SzXP1K86afyU8K3wid/O/+Jdz+n/Q3OyxABvKjwN3LfwTQ8bQrTjWerQXhRM67+p8TcFtTihFQH3
d12yojNkVnMtj+Nck7GtM0vQPnvChvz7wM72BQQMBGgCh+sPvcz1zEOGPzmsHZjtPPFjfyOuVtD9
yQKShe2lhKMh5ctccKyObrL6lbSRkogWNfgQcbYf1Pe2X8Lb4IC9OdW+tD9pywJynyefL/UCB8Mo
rdzLzTbS58ReBbd0vnM41A38OJvLuxlBkWIAEBwdrWdJLKzr8Fbt+eurUW/DF6ZlffUWJrN0SD/J
XwRhN3IqPTT8jgCErcrZHC6DQNYUgezkPyC8myA/6iky8YzKmL7Bam79dVdP5J2zuh0eqgRrjU/1
fiOTudYUg/EwumEG2jJr7dZJulDlUN+dXu+3BFxvQI/h24xMdQUfqJtHR8uuizcln+RCGKiuMdQP
//Dz6+BkOKFT60hKB1dnqJ4H9/tmzsxTYA4GEfeOcDNVy9/ukG7RF8COLO/ohflo/aCXcucOhVJm
d7g+3tOnW/bzjEAGwmVyJMGlmmpGE/KE8KaplmyhtySMicRQQ3LLNcqr839i5h+09uTbFlY/kZhd
wSLwc9PBbTyac28MUbqRKIm1W5H4PwOVIaDgpy3TxOECQeFCpqw8gYdXeNscB4weGafbBiDKtAcE
6E+9yS5IX+ucFM+Pp9qRzMR0ZbW9TrMXlwQ7Ck9mH11zIfKOjamcqsDEF3kSREI+E1IzGQ1rAukl
YpBJsaYG84gRDxlZB0DrcDJr0x7Gh4kFFXDDLhVER3RLMnrcyGsLiWCSapb7ryTHgB5QeQUcM2QD
Mj5KWJLGo/W/wg6i5NL4OUgvkxQgyUdfoUjKZgCYhbf7CPTKLes/vcl1KWc15wfK39ctE5j2EnSY
WCMwDzhoFb6aIqlx1YWacAo9tFP3uscgIpRbM5BQfZzI+zwjV8svCD60zmACoC1SIRLReM9eL+Ua
cO1MY9P9S7B9AHyaG7l766ktiJD7w6A/BzSsilrx9/yVSp9PE8014fdi6e6ZzueXjGHvY8/Bs+Y6
Q+2fDFIxHCsfewJfUSimCl88LJRs3hsd4WnFpK6d8GtnI3IuV8IFF5nOj+uHkz1sePtG6LZ83pmk
yBIubFUoyq64CbO2KKx5vjdtWoXuEkOyA5EM95bfDtogMI4DL28djglf5PqPfD0f0ARaDmF09EWd
h23vTHPHGZv9voNTncE4t6dUqzazDyyrYZHdOFbdLxv9dR96/RS4A34TWDj+FOOmSbhrdLo15My8
4ljT/r042rWZQp5IrIu38OFRmxBHP827j58g9ZCInjsKsbkh0XXf3ZySy8ZTXxqxWQHWlCG3qHbL
OYoBMz2uvKuh+GsmFhJqgfDn2tQ/Ub7aYa9p5GkuouR8MLw9bWSmfKu0hLUTsuEcs2lFRH40IQ/O
1r9952HkwofiZVYoDhvl87fRb6DlDkRXQ8ztW3A6LqMIAVwBxiSq/Jpx8tvXsRDun/Kt2EvTYS7j
dmX2L5m5BB+WKnoKModLSnQyu/PH0NiG0YV/eoecJr6L4u60eyeeNye5e5tLfGZAS4kXTag62YZl
3l0u7qi1n8HiUQKrh0x1piy13LFk2hrNaxDqK3Obx+LQJmsbtakapi8qKcNsY7GWW8cRjUq8KNsH
gNBJFbG8P+qqcK48KW82T03ZRK1CJ+gN6njF/WsX2O3EvEVCJEaPcY3H6KSVKqw3WatdwNqFKHat
3fWr2v9XsPBhleEF9W89K9fICQGapGmxSwHM7NJQ6Ir+MVWJ0WYaRf/RtJUgxIcMCwmumyDLnPIb
A5E8wRsqJ/oBlYQSqP5PBa5oEVbiaUvWBcBxPDtR0SdXGggCjkLmz4IB+aEgEVhuwjwzuoFnTeBd
9xbGu3rLfWukBvK/rjxRxqzf3YHRBJPIaqxI1eWewlyBxiD1yeGFcnM9ZaQU/24T+ahP3Jq7obnt
Azz3DYMBGxepKA7/KQC+tinimAWc29ulWT1pIZji7vhZ8nRQrrGZZooE72OAXQwuITqOEVtErLpF
zvOkJ6F3UfWIaVbzPK1+q/T+rtqc8fdPAyVReAW60JpxNB7kI0ay0r/J0db0x0+D21Px6stleBTY
manHxyU4YryCBzOa3HOtJdINojEUVxODAZ5Vg3Mz4D81ywUuY8WYXAt4eHVztAM8WWIvo1L2ZhRx
89aG5L3nWB3172QDBV24OwRLF5Ag+zwTecHqUrMZ8T6sINnap5kDxc3QcIn06ea4GXjJTIbMaA45
rKw4RLcBFOjbZTeLEjNUJK8yEBecutgk1q7yBhVFzrCjDTpnCYNPkkeR6dp/mhkDsErZPPBfKQFW
kJxyR17P2dfGX1JiVyjQNM+ba/tDc8Vi0UeXu5MCG65mmxKHY+MDzXtVVfwjYFGt/1bHP7KQDKja
R4H4z9kpaFoyoo6pYAkWWd+483XWoRhYDefxzg5OumssyW/VD6iD+Awk2qN8qEiE8BVvUj+6NUqZ
VhdnF7zF8wbDiWk+ntgSKQ0kUrhbEHcQsSmUANmmFJi8AmJd+RyaPqQU8xKyxvUie7HdtPWqa/tF
VEPj9DFo1Dh1rwu/FuLAem0cWamLfALbHabK6AyvDDZE8DfcLcpFDf+RPpCCdp0VG8AWkFne601p
JZ61SsUzFvqJyLm34r0RdCeHZRXJ9YZw5ZImi8CxIC0jT51FaC6fMfmOcBCNxc88A992nh0J3hy5
pkyap5gtTQsVuwU3+jLoQ3hK1qq/Fs202VRh1mAvKOUmiIqQGXMuQw3FpW1MpMlh5BxvMDsLEoKK
nU9CBNiYoDBmG0HZ6twMVgwi8+8tXqT6jJGhzdENDi/dbTdDq67ZTBGq61R2a/oQJVLj7nU/k6gB
8Fdnl4FKNttGlg9RRhyiyB564exVpX1cbhkTzjACssEnSmJHhKYMRi3jSzF85iLdUyC2a8LIvsrZ
Mm9vE8CuYK5HX156cALzp0T6Y/amnJmDtKQ3JYAfpp9HZ5T8hvlF1nkQAjx1gOm3ij2hdGj1saMv
VOYTp/4vRKxOSJgXvl5IH2fg8aSd2QkijTpT7DSa/QfJ0pJyDC3ca8FE6X1/KFIBAldJmQnFpjUg
UnEhG99eZznMSQzZMYjGctKfdyQSsNfnnQb8VOu1gGq2vQvAFNaCuzcsca111dWVgRkDdREQ2/ft
6YaZvquRlqkoLMBkxNEFCjRLt3OXtl+kTz174aifHuqjkpj8eENotVh5OLbbxwjOBqjNjybiGdoT
9M4UuTvIKEQ02EAo39Q9DWiLdv1RQl2Z7YHfjiv3mc7qutzhRiQ+tu2fMy2vicSIveJAuP1YEkdX
4fTl6FZYPRviI5V9aVSjxVix53GJEVfhBNKevM8n0ZUQyvpQwggq9YmDTm/9wRaCNks+lPmGRNR1
TP+woH++7knLmIUaiPPVB27SYRmm8zd9U9Jt4fPk58kyju99AE5MebihlRGu+jB9jDMTsConDctM
Jb/acg403s8c/i692Uf/CHufl2JYErj4yEbH6M3n1cvZeiVbxvIY3ZhrQWOPqgfSGjuGDGlZitpk
GhbwpaojBcUZ0+Vu5G6cl2fV7apG+EL78JeOOGMEQN+4Y/lqKWYLo+1g2e6ng8bkDZAD8o9H2qJo
ci9ylk00ELOW+PPXVGAHLGi9M95OO88T7AGtNmiWsG5PHVlBTCZwflqB2wbgC6i0+0rdFZzW3jdy
QXyc0UHv1y+vR30oFFvqOxWP8b0yx2BE5CWO2repPQ2BdWnf0zwdOhDHFEIU0WIco/vPdrNDT1No
ogWbnFMzNCNBageNFRLg785348h7rVV7qAKFB722wQ23ppzpP8LAqn1EdQwJZ1Qjq5eSIuGSnKPd
GFaTZIN7f615Pv8+cqmRowgTzEvFFQ2CS2kmrDs6KhZZtS75Uk/VBmYO7+j6/18WU33bRaWRpxYJ
8td4SpFB8qnqDGJEKaAyUWKh9P9xqB1A2A5QIx887+lnJh5bIdAZM70ap7/b0Ugcg65rYPX0vaxn
XEyviqkPYDZUOVsXrehuzVEemdXjxfdOLIl1RT8FiLhl0xUrRXBwxSNWLUoFvZTZw6b0mqfcoSd5
T2h5l6URQPSBiEx8IskYGPX9SP9N9O0oi99ZGxSWEQK/dNwI+2lMMbZZg73WGlyX3xdteYZHLf0v
LT9/uhUzer3h9pIENAoZ0cALQwWn3yHQX6wLVJxgWWAvdbHimpGoRP+uy2QzOtpZSTOpqSJnPddS
5Oq7JJLuXC31Fo2x/rIqKa1eoTJqYRqjtKfZsL9qhlTeXOUaoxrExUUhRGj2ymkBYiltn/cFfO2B
LvYl4hoHpHe6wXWwaMUEgIq7HkFJt4U3y9SMtCZPJOnfStTKreVvYRYH4xoKQ1a9LYwbq0fExSjj
yjtUWbkzbDUoZLQuAXjv7hgjj455jdru2qIEJkHQqohNVbIXtt70Fo3l7NZXXEEoDu+jHYqeyTjC
8oZ+RHgL+I6O//Fkg25Q93HXxGdbHnVlpxQtqQl+n5WAacbqczeRzcCtQ0dH8ssr/Y+SHgawWDoJ
BtpBaVVDG9NZ3Ty1/mLDTItL13jipIGbNxdyMLlyX/p3HptfQgNibC3shveiYsrOlEq6f1+uABjO
PZMFVT32PlJkSy7jGzp4+gVcTkCx2xOUTSG/aq0UboJJ5hehVO90lusWacIFbI3N8PmeqqMt+GF/
THNcDPOJszGSQ764S3A7ZM5YSA2wHoWvn3JEan/JlNFZw5OeYQqxK/IgTiwtsqX4GiK9MtXa9YnX
oBgXCyzzetw/Up0CwmKkJjwpIDgLCQrw39XcMoHD6LpFhzdfTONUlUX2UI7LBPGdO4fZ1MRXdbvu
lesOCNoDQ1oTVo2cPRWWCdHcIrKSg8WXtU9xc3RgFajPURfUp34LE76lkKrUjibdFfrGiYeva0ax
Lle0X+rjb7zDTD5BipAY7GFfa37T1w5Y8cTv89YtoiOJiVWQSJfq4WtV6lFqMrMy1b0xMGUP64nm
0nnbm9YPA2zXHnFhx0IcZQi0/4FN5OBlt1K9iqbXgrSHJ5bIubeE1GNW4CSRZXR3d0OsFwPAhw7s
30DpjjlAEs3VObXfaBMNplEP0DXI8iaepvF3t8Qu+TbL5C9JXuP9Gx+9JntrWa7FhiQG0zPT37qO
8AeDcl9q1H0nhB6LWtuQTIzuMhRS9U6WfokVQJIX/iKxffDGwdxbchvC/wwSt0jSrVtmPnhjvhZb
Su27oIF3tfESip8nhK6Htpd+ZmmLi44r0DAi9cUy6wirmUbOs8WUWM9Ygthxrxm5Lzk6inK2eVxt
C4K0EErgIRsK7TlpTViE+VgxN6X+16tFl5Ogg9Yq95cxsqZ4jlOEWKyR3PVaetDJuymAfrJCkpcs
ghudra+nxfjPhR2VXLNc2jptlSeL35EWz3nOpId0pxO0rmTLPWkOcfKOMDXx1vNSbImQe4kZa/tu
Aih0tbKmlpU/TtzvicPLJuJJZxu3UKzm4PPraVmMbP9C4qcA2eGB8sV5BOHCkTbeZ04I3m+S8X2Z
T1VmwRDTXL8d6n1hlA73WRQB6GxVmsE+8OL/fPZki5L2ci601SmgDaI1zITzen8xpNRzR+q9wy+q
BiQYvtjp8emgllWobt9SqcFbc2a2Qd/BibPZ7OQh3TAl+yEr0WAgvyqJWkdN2KJhazdc4IRMdzzK
5NjIFi9RGUM6n9dCUFpTPT7PsConfxxpM+s0YBFVsVdzyUKbzPUYF9kTrDiVZjBWGV+FHMKO6D5v
n2iLnQdoIgoddbahCnQstLqbSlxfvsOz297omcJKHIYYMTy7fRktBo32rR5Lwph0BvgqZbUOxegp
ucZ0pZ2vETDHR0oRaok3HSfToTNI9aS6GqzoIojcZECKARAwZPS2cweGaXBwldABgN4des5Gxepe
ZorSfQ/vHwx4HEme7klElLb+TBK6MfI97CHWbiy3DOoHKGKbZBWY6Ffd5NGdCyaQDha4eBojTgq8
J77nWE0LegkfvXigTwAS/GHIlijwBIcT5bZHHwowJPDK6KMCFvT5dBN18A6T3qH0gobyBK/0a/YV
2E6iUwDF8c7FTx7Pyy1Trs4uTxwxs8+5ttYi2OdWij49GVIePesfEb4OPMqw9f5oBawYMWz6IuJb
m9vPgxFITtCDVhejv4Eytqru6YdpxS7h38nZCRquQf2EaBZrz6WAdTV1hs1A4cilZd+lEHtnbZo6
IeBUCX6MOFXB69GJOcHaGizdoDWN4+20ZKroB3Uocw2rqBvXjFSfnvcuhOs7U992ZsyU50GA+PpE
pRxDDhu8DTZmXPFHuxwmRRxhlyvuoAJY+pc9q++M1f95nAP0D2mnCz++WXo4ojzA6rmKOpQFIHMv
ezTg1Yu+VP+tRcqhi0XkUSc9ucKG1VjFI2pCWW6Ysh9ZbNtbZXxHBBdLAfbfWgoWvwd8kj0tRFBB
4xBQAKBEs4aG2cXd9uyuP+YBUl1veVhj63hfkBbxx/YcKBbRcw2PBwp22F37DHiHFSGWo7gV7lVp
mo+noGsxwH6zfwWuTpYSaOZfKhx0pB8Rj1wHA7sy2YrGyICAb+E/LYMYFy0GklwOUu5Kl7upnlde
/So0AKSYLIslo3rBLFc3lZz2mcia9R+GZNgIo2/3FE6oq5p/6MwvZssr5pvSklpTut5OiAtr3QRv
dxu6757ySXV5kW4/SOl7pt2ULaiz2HLepcjoslNH4zsGgbos89lbe41bJkDDQosva1x/3Pj+MlG+
dg7TqVrMdGzUDw26azZzh4WGfT39YXPVpI1579vywX8NYdlLEpBbRMef6aboG4szCjPewS1v5fmZ
iGZT0icHR5jvuyFc0Gcm37QWMyXKrDhwMiNgUGluYCfaTe5MIv4J+71PmRO/5mgbJV2z/Xhbb6so
cdVLCZgvgxG1WCiy3WE1vhKKZfYnXAlINxivA2n9nUAaHXBnxCb9USPbvvp02WQ3Jd2lq7qT2dmC
Ba67dfmXLI3Q87UMUZBgCh/0N6j5IFAlbV4XMciOQsSVfsPgBhe2WzQPvIgM7gwAwmdiG4mo/ho2
sZRfZ7GxbZr2ezS4GD90le5JDibljlrPwEbllpgrpH4q+VRQYIMsl4eXubD2k6S+bjIALVku9qLS
FmADtS4lJB4LD2c5PGnrtSM6C6eFRy4zijsNmASb2Z9hCaExE/pq3tiXli+8/C/kKOL79qoNCkz8
AmMhlp0K7q3uCDPtEg/NTp3eMFNuqmjVh4antl9krAxUiEdG8BrNXE9CYL8rjJKZsB7uKjuz3zih
nuOm5oVmccZa8aI515oApzJ3Xc2+3+geMSUGcOht7RRXoYmEWK10SIEv2UJKJNDGxWpSzvSZ8NtX
8cjhac8hlD5bseOdO0NjcKBUOyWGVZMeDXeLg/aMzNaGp3cBxcIRqmytjPITeySLSmgB6UH7STPu
pkrdbCvz2chnDv7q6vqANMuZSeN4lD338V6tV0Z+svuIFf0IBSPuJC+qQCWc20ZvLcdy4xlIqYw6
b/IgVSjb7rw4g5IC+N2Y5Wex11Hm11FzdxI7v0ILEwv03Sc7LnBfetcS9cFqD0p5ultZ9/Dvo4Ex
poFE68w87G0UxpioLmQL7YDy931rgX/UXpTuLWJu/l+jm7RxRJSF2t0whbRVBW3RPiRc3icuB3hR
VyJYhYnrABhmRmaFWpBB74mYEqYEJjfFZatsl0+FhtRv2fLCSe5LkuGWy9Qzv9oLNQGDEOR0QP23
6mL2HPFcczP3gGKhbt1NWDJ443AOJQz9XWLEQbqBp87EA9Dh3vr9aJQvDZZSrU+ep+ZOrdeZ6hYy
elz9zSUf+qaik92Etw/hQjhLcATlgXwqh1m3beLOTS76/Y1XLFlupd9vD3WofuKhKFReeURWU47g
An5o6/T9iFnde6ACoaz5RJYOler9S6tfsUh/SRDXYsd+Joxw3GXdaKD4H+xv3CpvUDMztgrxsh5S
fjIVd59g7yePwfnxbpszibjxwJZlXZjOv4+omEGrutBbuK6mE2KtBW3GFmIBTIK//OwwAAxXOYtf
9xRMD3GFOLB//6PLIdn42yYqEPFuN+gjPOtGavpyAL7wFnxWWVbPvytRe5jdLHGk70u4RyB9/z+p
DqmGTvZclHl+nUrLRuqXLhPxOlBQ2JqEIo6mYkhzGzq9FShQubA/ofLf8atfNrehbZmDTuMPBMhs
hp6Tle62W7jFhef7ItmA3SOPY7GRXAOWZEQquz5b4zoW5QqS6fSAcO3I2RUbqlEutaqjzi3MHIoU
4YhkXyNXHCuNVL01YVh8ZPB5jCW9fMMWvBjfyDkNbBQVI7RbmbMikRVZVRMHN0bJfH+tMAtgj7cm
WMeRCWwIDJ41VuOBu9eJuxUioBUo8s2GHDp1G5UKxmBUTsEsLsWYEekIef6OoEoiQLRvipKjnVwx
K6BRl1729wF8nBwow9SFh+w97cHvAbXWVPWr15j+qNCSI1hVY7fg3lfYVFFCpE3ktYROxpqL+oDZ
ej0m7aIWsdTggka18RiTJt+19nhQyYJHTKPFeMqPo2dKReiibDVFLnayQp26R0ZTZHetjCeau+uf
HzUH782SdR0DoPdEFIefbGnxGYkle/ig27RzeG33Ommvj8e4Gqy0Dvw5tppJTKP60fPbRVPziODM
v6BY7kAk4TW0R/bnazvlaoufxT937r3CHHGza10HNo87CwOa22cq5zhHji9JeSPaCrQ2KO+sOUC6
W7rCBDjvn26ncQ7FCrpYb65pOhtmbtRV3OmMlCj+PDTQhmtav0RArP9ticnFEQlyQz9tr+dPDzBZ
eUzPwrtA+okkpjSCjiG1m/mES5FCUbGizjMyc68iMOyHTWU5pBtXNwgO+XDYM2wipJPIjIRTOIgC
94GBcyvNACi9QnZeHD1m6Mlg/axfRJ/BTALaob+CdyCASv+2wilWQ67xVRsgAxTNVIdgbShIvf6o
Zr9lAGU4AfyJSjN2VmRX9t1SVjPMk68RmJpi9/3Xcrw3lPErAy/6yzUJgzZGdQBxzhd7wHcf4wE5
PW2/y03sh8Q5aU1TzSPgbfcV6tFeeZFZuYlCLCErvXiPeHJs3LKCbVg7ybEtktlK685d64Lc/ivO
8y8Tqqt/9SYRkygf4Mat1Lt+lilWbNupJhe92kcXMWL4wNdCzcWYTredvYM8t3BX8oPnU3TSnDEG
HsKhd2LmIFuwMqXX0LCw4pNemZYNJz30xoze7vh0Ld17jrtPio6m4i/kn5vUjVuZHUu7Ur7ATvM5
Df0gWX4JoR05t5WWX1s96eX8sNfjVblxEtJtbEOHj7I+iyZDn3cD5Wlji0jEXi8uHzDzqtB5Cf0q
+jDjGXlkl7VfJkXNqLVs3TWmV6ME40OKHy+tQkKqglqN01ELTlkKhsrQoEgNVI0nPSdabwteRwoO
cK2TKsDFy/ug7UrVZhamxn+0bl2ZqkYHhOLA6qBlSUILvlHESDu+Yzu87G0CpZThP9QQFNEEmvka
TPgpom6cMDosRxn+MVKZD8Picem+uS+PEf0v/caLBAybPlhtwHKQxw5QVqCQ8WVPi0oejWSJgNuY
v5ngjVTndXg+v+1EpxsphGyuis47VoYam+bQdkX06Gy81NJ7Ug7CX259jSE34+tfWiPR3YRRG/eL
TBBtPBR4ibWEBNah1GTLT1VhChr63uz6RSmKdZrTRaqlfLOLqEwp0Y2nkTDGWrIFO4x5TBPgF2Fl
Ro1ckUpUSATdFqQbMRc+5zBtf4Ncmoyk/sznLehWX8G2J8LSyJA2Kx7ixDLYSDvISQ/nfBopPWZ4
1ZA9j27kqYJbvmmP/9UwE7GAkYbn/W6UWXRwJke43ym6aIl72tf4MZua//FPBpGo7TPF/G3DeBbc
zuTJzXbl4T6AfK8geFKr1+eXOgALB4hRNbesDwfGSYVQLEKwDE86hYDW5BCqSfU6QHRScf8l6qi7
0HsMTi/Et6zBlIr8uGQ0BEjVk55G+XbdqPMpL01YQzihIaF/gYPLdIpH9DisZD58rjU1NijWGjbL
FIb5slVpD70ii8Poq5dzccmv94NpvclyutOwS8k9/gIMylaGWS6KZKHWX41WN4/X6aPT79qiTXQg
k5i+51jyqvpca85bJdlUiUIxIwcJhIWPFgVhSmRGS4CnTkN2nw7MvWEwHIZitnwJ9N/jzflXa558
JuoL7xgXaZ5Mnu96HkN+Ws2uEmuFKV09ZUAkouxUYeUyPQf0TmIOwIdU8lqq4IL3QAE4FYoCpqvw
4H+GOTlFNwSYZEHrDyXMgomoLZ3h1GlS+hSv7sdjTyFC5zp4RVk/JFkkihFNTA12e7/YIYY0EVmA
MPIPr35s3U22ap1Lk5ghpCErv0YhBdfiSDZE15OlG4O2RmQtHRHKXPjuHnhUpySKei24mqV9zMyG
rhhugrkt4on9/AU6O1DJaEUeQcnUi0pWX8kTT5FRwU0DkwI0FDzdvdh77IM5VSa2SDehGZb4JVxs
vs7ZdgdUx7wO496GdEHOiZx19YEwZ/7Md4czZhOI9Fz4qSULarTh9kL9DxjvRpTe6gnsJSNGQLCJ
7AQ+VncnKrXFaKUNVNBGbia2ETaGM/Z33vBntESrNX10kVcl1osecTarrxeHk9U00B05qnvAuhpZ
Ya3K7gDpVnlbTyrof+ICSnqdI50c5NSU8TUl4QYvDjXtglHvSHXVPYfi4gdcMz1/lahHjp6n+EXi
HaiGcbtiGnPYLTL4Ln44AK+z+LBb0CkLf2/v2K68UGwz5K7gGHA92AVUCfmaBOhVlyeAFR7ehBBP
3VQSvqyPE5HBrVuoCdjJhw7Dqmn9jIlgUUbM8TOwwoDxgP2YyfpCwa6SXqY7z+52dxEO2MUJXu/h
APzM/gd6Dx8wBnc+IXGIyDCQYZnz++PL13k5Er3nXWPNxBBeeRcT/odC2xY2sTg30EPAzPHLTNzd
SKdOm2co6oANCIcNqpS4dwnbUk0qbwrXsGSSEW+KN13NHyeIlRqBgk1Oycy4myTbp9ZT5xB1K34z
/ecMDQg09NmocBWSUWiw7MUHsiOKrcG76/A5RHpm71uouQ7VHrBZWH1La4ePiPSjlD4N1Wj+Uxiz
SizCWJhjQ+sTk1+oAZOSI5Lxbc1GFAK6H6lEFpeOA6FaXEtzMKi8LFhgLAjOZPoXjwUFmimLKcQN
0Xbtgw0daRvEzFk+lMIr/POoG+K8R92Thl8WnPtWCs9GBy7J+lo1tZqlpL7GIq3fNyxQykbIl+EE
TPquD8g+GTo3oaJSZLZoSJSCUhbXnw0iYSUaKoDauv8CJ7vw+ltxyxr6uRnB9XwryQ7D3CUt3a20
YpKSxIlIeS5Cj2x1KNjpjvxYqO/VDBpvDtRsLnHwvjs4nFjhL+esNqugB8ZlFhK7G4OpjPKkuStO
QXi+WYw0Qpgt1cyP91G4VZaht4bzKwsxY5nQz7WIATEtvfASESjOf9r8DjCFRu8qSNSTegYLSpoK
ikoNyDckE/WAkA+A1KO31ol8QqfaaBpQTr+8T4HJLw3vHdbLX5RpGJmVXSoP35Fcp8IsEM9FnS59
ivscR/b6KLCjtUGfusiwX1cMk+EEb39JaYUnBb678dpuaKfl8lPEOJSehsBK+RqBxEidn+u9tHVz
vMipNCFutjAzPgUg5zxGXRwerOATeWUldBJFDMb5UvAFP8ACzpJqH48VoFXnArMJNkeddhK5jd4Z
i1pq0Mx1L5DnloxIpn4K7EYFCjh22p9Y5GxScbNi9PeBeKVnecjtfvBsY83DKraXIiEm0cSkiidi
TE4ZqIOTu14Y07N06g0t6eQs5/G7WmS6crlgcegEN/CTO2AI8FuLF3gzCGd+97c+TSQvQS+Q3Mph
rp+6fSOq+TARWciDP1S1FWHLTmv5ns9V5qeAH3iHhcUgBCxdfh7OfrbAoLGf3lZLNDlbQQ8ka1RF
LzPuR9TNsEiorDsKowv/VhWeyomCH3BjH1RXms0123giAxfhgi86Hhcx5vKQjwXzVZ5a9kOzox09
UlW7rBuo5rsfhPCjI3eVWGllf4MpJMeJ7Fu85vUaeBAkjWGnDIubnloC8YTTjNWoeExA68J6Mbh3
/gGSPw2ICePIaFliA35LPtqFjK/s2gHsmJtofq/XjCAOGnx56k2lFuUVYBMoAGv2V7d5MaNBZNrL
HRYhQuKe16wrtAG1aHDOlmr0ebv9Tgd3CUwxULoyhlBFL5XxeUauqKWohV6A03VKFaM4iCwpRPjK
6MD4vyI80ncuqtYo/7109Zlgwa57NgqpQ0DMUogWJM0U5cwDyu3mq4PamUXqHnjIO3q0DFqB4g0X
0EsQKTPUYhdUHLjOH7kaght7Fa7M94sMX/UTLpNVxjb0ULsCHXnI2dwYMIiQgjsS5vupDnRE8Amh
8PJFxVHW/uJHTZdzrVxE8hcUr9JQYATxUETnbDTPi9kyV/vhaLq+oVpZhTZ5LqtlNIdfh3uJ1gNw
YDUufQJpbr23niBEWbcO7k/17d7/nSYqvR3IuJ21Elk1BQg+2O33M6+sGBbUPGG1Ur4pt2FkqlVg
2Exs2zIY3Gw1vEfjeZuiV14rw4/fpP66x4HJR513wb8UmL5MR0xqqmcrEDwj/UIq84kuY8E3HMrA
hU+s1okx+bzTpLyJFMFRdm7HbziDjmW1CWNqLYRgAYA3SKBoCMg1d+Exs+/T6MYPfxGd5854LurZ
swgTj16/lyDmbzE5W4s/QmsrtefovdfBjrC5egEOVkoV0SKgiNrBJu1FPa0wIGbh9svci/S2rZyE
PPcPW7BvJrcQnZYorDdPePCo1ndIZWMq7TDZImKTDvXnNb08ms+hG2mT6TBHH9O19Hzur09iYMmS
1tYvsjlbVWkHNESryaTnvOF8uW6CSkb04KSTzt/914Ye4B9FNEeD0rQLUcrRvSETjN96lenVj1Wt
0t3emlZ0S22HOW3xCPTLPtrJDqUtFOWGipKgShhVoVR5Feo6XdQTb3ML4Ms8RvMM3ctj5zyzXCIV
ERx1KwP4CS9jPbmforaYubAVD/flVZws1yn3SPlI7ZbkUm7uG75j9IPYdSC3sqW6zjCqys54y7pp
uLA2xRSfuBns3WNhU5G2Y3ukCO2Y75lF8O8ly8++AoivirfC2cMgYS844eirZzN8pjHIT1MNrqvl
U8bydfrcjLB1yFASRWPeZDB0wyTgN/8GCMNGnj6/luTTOAjqBX3Mjm7O/NmJDEbgysDM8D/OBMPM
DevWtbEprb37iQ94miIynjzlSprz9CaRGMrPqv/4FsOltAKAkaApO8ZMBUFTfhe1cS1SZ9xrIDic
U874mXbAZtoCXZI4AfoTPgUER4fD9YcZNKjQARHlVUvYCdZwhGmIt1c/2xuDmoNajWScMpO69/fh
JIMweJb86fUgRZzVyLFcq+RaoMhlGmF+FpA4wKLluaN3fdlgtOmQd0iKph+NvvdQVjDT0KftbHV8
YZQIPd6LM3Qk3m3bUoPLNY8Hrf/uRBGgm9KCesBsdOZaBLAV4T6iTUoGCAoUQMeGY3vL3wseCve5
jHFkJO4IJdNHheDOVa93ik98aAizlDegrR7YOIqy/oV7QU25sbMDFIGP9rX/vwWv5nRjeiEgrsCy
xeFObg05oKhMmGRtpKjFDd08F4P47V5NX/zhl3TKc8Qn27SHcKSsf6ew+78CKNl0tKA/Q7XHLIlx
nbHP3UMXKLxJS6uk1eKVMMl8jiP6hw1Bm8jnUUpyqomz96f0H9S0L85221QXlYJpKFP5+3wBIahu
IMLX4DoOVDrXS0SWa+GUcNuMhJmlKi49yVpoXAIIJFKCYi9HE+VqAyS26AKE55FY4y/7AbUpT6AY
GjY+A4OPQKunLhjJGYUm4/PEew+DznvGjbrNSPciiwJfSRcKT+ryxBh0a5BVgWH31QozYkDBfV3m
/5SXRGDngoGr0eJdgu4Ui8RJhI161pYMKxYuPeRf9R5L/XzZuPq8uRz6BEkEM4ufosDVDhHczPmS
qrvpffAaIZUHX/c5kGNgkZ+ZqSRKqkklr6Jb1dOOjJMVq7qz7wCAQ1QQB6eutLichxiFMvBCWb6A
YigZY2mHXd2nGKKkPOfQrH6YR7kFNypwJK+m1oQPJt3pZbBhoC8G/WkcNHGmMEhV870b3bmu9QFU
yVMbAInDtr1DVzB3j1NRppcyqhk/3t556TbI7u3myU1guYIq+H3BRlsGM+AZgVtejxW1ILErZBwE
d25A3aXOinBhPbUf6CSUgtYPOUzfbEsdYIq00Pmz5Wpwf8VqnGU+wXyh2NNV8B/qysCebayz9yFU
t/SBYWygbkEDkfi8HZLGGhQ7QKYzwcLKnlhuw/89RKFTY6Rruscvb9DKdkie840oXPXHZx6JCDfI
KGuUzZfHgZWFPXcJx0gbNszgUL++6F4y0Tm+vAAyQmuutoo3sFZg8+J1ULOy8eyL80o6HlNJa0iI
brLSemtRABK7Oxbxh53zBdomXSvR9A45/MOnvck3vVaohISoglrZr0HdGtrDwgctYfg/uyMsEoHP
Jhs3kulkrjdfFSdYK6kfXzHnZsxv5BT2uC4fhbhvjv7KZQ+anW4VLGHhCxlF3rIfaqO6l0ydj+kL
zJlZw1b8G6XVAbXMv2zfOGkzBbZNZosFHlqA+LxvNJhDAqn8u7B66jNethR7ZtrmyBpo4wuZYs9n
QeezQ27CykMS9N5sB+xLLuX0a8QZfnNbjqPiDAQImUhQHexUJ+69aQBfAYaoT7Dpzcwco4ShxJxr
cc90hEKt36oyeuh6v0cwGdnaUCrdZc9p1WgHjo6Rxo5VhwCJVR4u6WZR2NGZllwIIVMpOtfoneVP
6DBTbIyaNiCwiuaKZu2bSJI9pnShg0rc/rqu2NTAt1SkXnmfX6AKNgBDicSntaw+KxrH1ieh2SX0
09tn7oG1iDxYrCo3P9tKnWqw7boErBPYN/zgwLXld6z/Ja8EMN/e9iOgxVSwm6SlaPqcQQe5zol+
L4KmqPZYTbtkZo9B4cNAk3LmWLach28CK5uIpo/D2N8u7wtbkPfyeNHng80IYrWwM8gJRn5ejol1
mAltb2AIH7+QDJvkkoQEge8WjYL2/HzdAbrd+BKHcXadh2M/Ib8WlZwtSh5l/HQWDMTQTZ0f3WAC
lbafoAgTWqjzWRqxSmaLcPLY/rxceuO6zOb6qL4tB1DQ5q5coCdorxAeHXytTXncghTJowOnrnlE
NFfJal5L5Ah/zVa6Wm2JjnIUwdzoc9PEDgWcDbyioDDYd9Q2fnjapmgyAJ/siZhq0EqMrUn8lI9s
2DlXOpn+MsOZ+HYh7OUNrWB5rUSE/3uGCQ0bdl/eBO8fzylHLWwow9jm14O7Q7zEK2Rx+SPIfxB2
bLwCMS+e+5Kdl+01NopOVpwnI2/XsswXiMmQvvGm1O6Z8Vbpm8ytOnkxhP3OvP5CP0G+m+BkKc7P
9evaphewBrMAAWBxrbWyKtRAAmZBgIurK18dHXsa09Acf2nwwKbyQSqYOyYDxqmMYK6K2HkNX50i
5tjAIoWP8t/oP/JvtxbCwEJ0RhoTwRQg6sUrBklTcfpa/dQaaLjiH6nd2vj55p5OJ/igJ7BEoYyD
dFHg6u+4XR2hEeKgi77Ar8kSraHO/SknlUGv0Xn0UJyjzmsK4POEXeWngp4KjmCFdWVShgZ/ntrB
djF3NtWy0i4e4YfV+S39mfKIDNHEnC9Yuvryf5eoOnqN+Dr9U8xwv4rEy5jPZ/SvH4CRnRfuNh43
FTEnCrp2lmRWN23n4HhOt9+pybIMojtkKqZobMLguyGagYPfqTiL0aGak1pR6zCAm4+5u3vWDHV8
NCS9fa6caZ8jnQHOBgH6OsSJZ1kWQRCtmJOaPDH3kIltXVvcdZt5Si67f5fKk1JVvpwt25v7Or/F
aGerUQJkYQU49AdNnovbq3hUH0lyOEbLJl3NMBdl0ANjMr1JCH2PoniW8qKyAuppe+dZwGiTlPhB
DjY/G4rhnIGEYUlmJXVKZaM3TUcGmuFgRSlpeWj0MKfwhu6mqRuF7ANLW0RCZE9f6xNkX012AHzt
sEjz9TQW1Uidxu1YtX8C76eJwjfJVrazLfLcwE+cz7YDIY1LLWogD2zc703Eawzv2psNTyQpXb/P
eom4CDOnrg74q/lbjOHz25UFxZqwGWcE7y5C8UlvtqX9fKJWMv9rc1/jvrvABcuyJ3hIPjsdVWiX
H7X9gWdsu6t9NQI14hhDqiSmRQwDvGmfCqpBvjNocdWTQO3gtWUizx8Qrro4QUxrAOBRyiMmr+/G
4QsTLmHstTOEnte2xGCkz2hmQfkazdOqfB4geU2onSQmdugKqXAkqP74SplfNtNr/DuzzQoBDHuC
kBcCnM+blgg//gmB4Jjjuc7yXIUKZEFftMa9YojdDRPwMMYdeR/4vOD1zZ0uXyS0aQKjuGMaEKqB
VrUmMLZ4Gqv66nM1iaBIdFSj4Z+RMw6bH/NfssQsz/hblA3ijUDlmsfCos4iAsZzDeEc6iEkUm3k
aP0T7bF0HSGIYcdVTwHNDtUQCBPkcIse04Rw2Ya/YP29fkcXi8zlwMH0OCICzWZRY2VI4eNH7gQ9
Sh6GCqn6XStZihyt8lAs1XLBq/5tRlaqOKvJt0LXJJXMGXPyLkknZpKCWeKM7jv9iR44XRGPw0M5
3sgSKS8HmGbbtO4ZufpCrUA+mbC109VxfeM9smWh984qX1NU/62zOpB/z+IEX3C+tn9QNiAzj+ER
aC25MZmLHp5755ewys/NEosvDvGGbA7kFXh48xhv1DG0o/sPu4UpNLAnVeqt95oxT/Xkd/dQXs23
Yuy9loat/Inob5sEwsr207q3CnC685qNWRnA3ZJsy+z5QOSERQeNy2zwg5iWRHR75SH4HRlGzf3p
6GT1gDREYNlRJjNSksRMlpQdBkXHUcHkT6CyTgD/iI60ziEahFfduxPPO7B/pq2sa19L7u/UvE1c
fY/VUJ7WeyLuCeJCJ0cUTZpLpqLMTUtaXOe346/CnmUpUi7aMSRZLuHpXFbG1vJc0GhMnYxxyWpE
5AwJ4Dd1dLjie/WAs+6ymB5DKE4sCKEySsTIpCbEQyYTCJueZ4DlU+HtU75ql4vTYsSfPxq8hD4h
saV/xEHX57uwrTDs/fprB6JJDUNdRM9F8eSC0XFaPl08ptRCmfPey6F4Qtvaaj6VNK4FGxIOlrtB
qHvN19zXaTJi1rHZ2Fa32xEVdYVnCIfmZUOa6WrAagKLpsCC2Dr9nRFIzf/lldrOC3UpD28sC3uC
RoKqB4ik7eSd39rMypZhIi8DoDQxktXKNF+9arMtXLOX/WE0PUV8T1Rw7mlD5rukvQ0F1MTJFOuO
qMK/hBRMwK8t3UPw9hlLt615f1SKdCWNTtUyLFIV4AlBn/05OjkwV6t1EWrDcfWU2LUBPUnK9jvm
BJHOHBs1Mvq/A8vTV/xCYIhEhx7bfrNNv96ZhDzHk6oVtD83gKwGvkEs+yrgFwBL1dT+dH/mhQcg
AP1vJMzhqGsIxnJJWHsVx4gfrbTmj4TeEGwKPhDRpF4HN0TI5FcxZD9uUJnRSDELIdHPRg+k0XYH
Y8V08JoMs7tY11CQdu272hRurXKUpsdBLbse/YujlBL/mORkrvpfvwa2LKj3nfgcDiyz5ONM+zGN
ZbJEyaVQrYBGNsmMEJrxUnA1/WBFr78VzW7OrWG27TL9N2HLt8k/DPBWT2z+giFmQd7tmtogqiph
TKvTx7PBnWy7vbiTvReAy9orY37A95Hql5lYIeIY2+8BboJvXqMpjAb7UKcqyvrCM/JecBa5GvDS
F2BxlMiiv0uIjaY5Azolaf4T8Uiukt/KLKU/LiMP0ykxCWHo57YYJ6yCO2Gki3YUNEMPzVOh+eSx
oOrieyjh7t+nV5O1y//2l1UT7Q9E3z3JnhQW3zSYZiXtLo40/mY3ZrbAaYxg9vtpXUOL9isKYvXg
cfd05F5srOBJ2jrdZ/e344l7AqxVpCVB546KQFS5w5I8xx8dkjiU4pu0WYPLNSMWUQ4MenHiGdKZ
xMszhDtQjrKNqmMWLM0+UU1aS3au02/kxRrPyeyFvnJio1+lVV5VrSacGNcze04Ev6s4RWMVc4p1
8VqO3WFwTEFGt2M7a67Q/o9+UJg8DDC64BVPR9/TkdtuQkrR6aFy2M1VEwpE0B3pd44JabHsnE/X
l85MxuzkRJ4lJ6y0HL94Hzn+Bv2Pa9ZBWVR+JyLrNZe/EyTxKwlSsIxwLfXZpwxgLMSsCNuXhjkt
MbjQK+pIxMZUm2gjtzmBLOvKyUIc4qCD8mZpeC2SOIUJl/CM0FyXnJ/C6OMrglLEGTAQIWP8GDBh
BdN+tah7R/kDXUj+Enkuq4lkRRQXZhy0k1rc2ReSnrEavG5y+7Wnk3tadXA9nGI6EtErn0K3J31K
Wa6P4HhurM1R3BT8RVVsZb0DmLSNOs8B1xNapE3/1ytvdvyO7H3/w+6TtEhEDoRe/KLX8j8soxDH
sWByRdJiKskEyRPJdMZTGcqy0O4RYXP2Tw+CHE9pauXtEAwYpcy0X4PSgW59kCfxi6FDhqz70r/E
R8Y2D+Cse80UTy4+G2IOzV1Fiu21uct3jq/MWTT2beDfMXI/30y7CvIX9c4znIq5EPYJetvUw14i
I9ZwqFmGxsXCLMLwDdQHcnLyffx7CgIJB5pAKlG4MFJhqiDXbDywWUVfSWZPVdbmh6a2HpMoKz4E
fSoJaEvcxzDZMInjhNaMzjN4rdGWYa85VF+MZKngdxs4kH6gfmFI6VEprZQJodBRWuwDcgOHGVNj
nh0T3AZtly5XwlS1wQn35q0r6x/0h4huwbN5I2nqojeXXdwSnbi1BSZ90QvH6Nc1F/6uHz6IlWxd
Gqxmn10Fpx5HRXb1Qnj1cpiHxL+qrqZexxPoh7biqLl15jVJ1Y/3FKLlf991LvG1Xk3RTxljTgXt
7MHm0spV9fvxJjFb4A+3SIbpDrlJF7BCiOSeyDAwmVa/5dXau+ye1wAejMT4weawKJJq92XsomLv
cP1F4fVVzD2kwuF3BJz+DfsIT+lHsd0nQJGO/FDLkmhfktdVMjSWO/U6b3Pq3ItDa3g9mM2j1qYg
7q56ODkCSaIgmByfTynuRZ/jXt6syvvCRSnxs/HE/SIG6ekof4NTsdS9exa/bfk4wsnSH16VsVMf
8B9eo/OeZMIbDbv8oiRBjaPbHwnds1QWEjti4c1qzLaiuKSz0hl+OW1Jd1B35s8TvNBf5A8Elo5k
4nISRxk9fMSfplXMQoEWGRVb97qkGfMlgC76cdUC0cWblyK0J/TvjVseCmsxbnH3fzNNuEOdN4y1
S1RUYTyDmz48sIZErxodJ3zCvpBAOyXBbapwmBzo4z0GX4BDS3/ySPfGXItQfqCjT9I28btUHV4w
2j0GpIpGhB3MfPfKBBTNQ3tEqMfeTNGcoelu3qIyOE3yHcJvlKVfalbR+L03KuOUTpaWPj0aWkT3
++v9+OEbAgt9rF3X2qrd6pqILYwynDLGxVyhTKPBPckX41CMpE6xrsaXcv6ddMaNmMUHMmotIaOv
8sYStdt+FhDZS79f92sgOkU7O625x1/p2F42QAixgM3LpqZJ7dpvW7kEkVEYKzqFBVW3lDMJHBYJ
QjM0lWbPlKDob597uVgKVdH5rFXEYt9WbFCG7bOZGPik9IOgrCpeBIjiSjMkbxzKTKjD6zeOHkRQ
J+K6zYFjW43u0U8k4FlAxED7SbVezr5Vc4zbU3m9WyL83pq1du98Ex2P6f+Z6f/C2TAbkIn8tV3u
ALVdU996XISEprQhco3mnAzndm0jTtvwh+TIDDav17HIr7vdHyOOLz/DaxP+sDZWc8ETHaIMptt3
geKVEwCYfAl2Z7B2KdRXVbcGX5lzPK/v1mpz2dapn0qkEOZChRJ1znXH2y4siiBD0lZB5Vo08rRl
xrgyRiOUXuOyM23qFSpYOokqz2ZzKIXpfvDp+vYmUPYIhnYwcIpkGufq/mXNAdIUtoSs0OBjqdFQ
cGPF/DUiFrn8XMARPbwt8ZNpVJm1YARDYgkQwPT5ChpijiUSsCLvBx3B7EEnVMg9j0HN897ai/S8
Hf4l1vN+nN1aiBKFnHG+rWkPTTWiH6xOxk2NlGn9KB3pm91ysrIvsqMPl/PTAoUY4OZBYrlsu651
RTO8x8OqzT3gx1tZuaV8hspERPP4P0a0lCcDDKRm32p8HSzQeDS67P5wjo6ARrilbirMvJAY6W4/
GdT6VcfrEkpA3umu3JjTXq75/91Q19JjIV2uA2IPzZuF68Rxxi4nJgU/NbhaSmATL3S2xjeGbroL
x4Ayyv43mvCoosE8mp9XUeRiHfrqG8QUDkipJKftZaBLRGgnxKroiGnQBOuamFeKAS4qKWPJCWj/
21YVwP9KcupHPUi9+v5Q7d+rKxKe/UAkZgJHVWCR6Tlo4sNWWTFgtTErWXjlJ4g6uhC1l6KuMkvK
KgXeLs9PMqO1ZmOwd51iUpe85AgI01l7d0dNVuYvPnq9OgUAh0oLC25G8m5P0Pen0avYf5dmmbap
2MlfLSD7LrKKPAHbUUPf/ii6GIdMZbta8N+eR82SIZPkye458qSKVF/99yzVLhhhskBARz2zKeOP
wzR91W05zXZgTNl46lP/obfBW33cLQ2L1VPYQttBftLFvVIjeNu282zj3N+3cdc+e+Kcd1kIC5A0
4Y/VQiGjL4GYCKT7Em4JcbvrlCTiV24gJxIljsTmiO8FL8AQmgWH60WR6cgvbfAUnQrmk28G2nS3
CtJAGA65TCfFd4jDsgReZuL1OXct0QTxVIjlT3JvgBSo7qlZYkbF0udVDgPw09pjhvwUL/mEdBOM
WLqSZQ4NolbIsZ/ZC5KFPaFM4HBuB4bmZwXwmWXtnqyUg1glOmrDgMRHd3gX718PMRIXPZagLf8o
Q0VK65hCOf+u1YYh4JbTGlNvvKd2iT0w2TPr5NSKP1Fnm92Hgu30Wgj3ehx5eml6AVFUQc9luU6R
0U6d2uFMR04zyWFwledNDGvFryzL1XZSU+wUjyHqjUNQ3bC0sNa3wR+wpLk0mAspxkijjyLXMN9c
6z9B3UOPjdul1S2MhtPPOJMnQ4Y9Ux5r+JCJMb01JT/7QEcaPty1hjceTdZv/HEk9oMUJoYeXNRr
r86tfqZJPeVVXoo7zMwoWBjyeeDLS4YSndGVwPmrqSKVcW1sTsjgkxOcdvl4MzmdMxdVLdGQYJPh
Bv7wFvzVkC7MpXn1VIS5n0LBuwz5IOaKuSMJUd6Cia1dxAKt4PVCJqRqmlWoFxbBis3IvCE0K7YS
eErhkl8oWb7xgWCs3eKj2YMYyYVdp7ZEC2XznomT/+lZcxJBDVc5kSFMysoBM3TaOre31algGCqs
UhJAm0KHuEW8PorLfTMUip7EXZU6IiPI5I15i3YtC5IjCGaMrAVPq8kxhczJT92wv1g8gSyUMU1B
tjRVxM1P+bZxauSfCHQ2EeGVVxfOl+wWaW6orDRFetCQgWJjiaHeR+3H9ht/ZEZ+nAshe0je+QFF
+OBMtjfj4/Ul4LASzeSzVYUEn55wR1HoeFKWIC2EQmVypBVBtortVnf0CW8SkV+K2e+ow0E86U/j
wl4PmDlmQjyz9tyVtw70rLcWosw+NVQR/osfmiYiGXjn/D4XJe7QrIDHJpTBDPIgUMaPJVYM3Tyv
GH+/D+s2lkyeLXdqWUXkkzHN2NfngW1qsE3I8MuhkZZgbPMuIvVE62m6cZcJhaGjTcKMFFsoe0t5
0z8qlWikr6V/vdAIeUSqE8SlSblkwwP+PxK+HepL9+SBmCAjUNUcDKipoieRcyLA4gAVnE0CjVxS
W5vY1llF/W5WL8lfUvCXTTL1XiTOueGlC84JPv6WTWyhPVPj5sVeeN0h24mGUUSrcA2k089vxlah
KN8knYYiLHH5rZMFmdXAGCvA7J1Usyu7LGu2rnUFByRKDsFOF/TTEGglhYbNtW8Wr2FHVVEpFqll
G3xUFwR+MRQKKJoFt97M9WNhc0mp2PNdOoAnZM9275WHNUn0nG9TvtuOxS1g0DIhcHtRAW/KDF9y
Mk64eAYlFH6GCqnWDarumfeIqxt22p3eUdF3bohm2lfC1Iz7klg96nSfWvC5LRPEoVitW45GXLx2
NvHaAsVzOeuhRJTuVw+KAtKEkdCUJNnhGxRASZjowWnR1FCRtUuEgeOutouv2BMW8LSC89pubp2k
VTF4XgI6Osc1XWpS8Y2Fz4jW4t8wLqxRhMl0ZZ/pONZlTzWyRxklQAUlm5HS/CJFzOaz0IiRJzBw
qpiOnFzdPJ4jxVnfMTwle5dmlsAYsYnME87hFqeGBbhgfOjYvJdqxGaRgDBOBveWaP+5C/n41YEh
hclg3Ud1YlrHgJQG4RwdkrWyjIir3eGXkBnN8+jcI615adz30YsDL3P4ADgpz/cTzqE6Ad8BPLYX
e6wbPVguhMbcR3mIuy4EAF4wQx5c0gJ6FKl/ynw1h2LzpQtG1K9sAdR0jVzdatppxHj7V08a8hEn
4aFyHHCB/Ma1vK5+HjfJ0DBwIE878jX1Gd3ova+FsU/v86Wenv7XLV7nHbcOT3TthS2Fm3E9r45x
iUlosQt42pGpwcIEbHpQnmrCngwFsTNl0avHY7+0Z4pbrWM3kIc1JmDE4lve8RQ7KE2bZAxsvdnu
8wboBcbDqXtMjZQKmI3Ug4uUPXmk6L+KohMACtXV0wqKqFUGSELJz7+1H2t6EjvQAhFb2C8bBnOK
9Hh30i2N1ieTM8MM9zbB7Mv1J2cmnLpQVAoE8pJNyMZW9d+YlhKXDlRfB1rLM+xk9thOd5UHohHB
Avcgr5AmPIFiIzW6z4yZRG7fhGYw1Xz048/30zRHjcyjBu0uRT9Bw2gWo9VXUy51bb4mEAk/BTkK
wKvuzEwNfSqKlAMObDB/vtJEjEH9ZCTwFp9cKJX1jhirxwwZanXDNpppp5pr9iZGwvk8jbwq4vFD
KY79RKzHxgV6ZwkJTx5oNDUy0kQZ7KArC5mr9Iw/mIcYqkkp7/hYk1cLRlxA0Rb/K5O6xLXqugpX
gBM24zLGpohHDLP9Slpn91WeiTvhKHW61mis00fc8iNkDbWutdq8QY+5NoIlEeEjaYjm0BcL03hI
T6ahlnV3F7VWLAzLD4MYlYDvC3SE7aLN7Jv4FZGZM5GroXUm/XGOV4BZeyTNwxz4dxIwEAH+4zc3
9kK37ngRvvKsfYXLhq75PWJXUaHyZuZOzYTVbZEELsLd4LRkwrxSdBTrXmUO5DvZ2DKdICGzfQDC
d/iR2lQLfOWAdeZ6D7keqBuCiQoLgLHJs3V5nf654e0guNSSQvepzk8idNNe61Wu8+djQknhvzk4
rSccpNrkIU0inO9Ey5ej+YGG+/OwodudFywuouj/i2/P78B2LLYP9/UGoTtR04bnCGVuybOboUYi
w5XEPnVcSqoZj3tUEPmMxiTJtq8YiwmR/uHbFOCSSWj3veXIPX3Ku7svHbE6YpTqPzxVrDHOYHcu
uzYonB5MtX+NwNP8DWP5QU3fuclTquU/70nGSla0TSspHq/FtFprzuvqCt4yWpD26qdpI4QG1g/Y
tkqu2BUoZfo2nRBLJnacV7zGO4BII2il+8SY7SE3lM5h1j9g/qw9/wT5seisb5LhiDaXRX/6hbcD
IBlVjjDXDWJtJ8daw3cLD/hBjFViF/EN7T/M4J3Wr0Ei7XwrppyoPwsm6j2ziXENU4XIVPtpwWgF
oJRGtsPkirDbyS8aCb+KkzWy/2M5KH/C1xTFOd19eWISs/4WGZsljTlbcBzvNMXioNJmSJdSJhSt
HMOCjWrcsgRL6/1By4gDT6v0eOgigFwYjKGtKSnXlO4bUL1RyUnpBTMePg/ItNB85jJdH4deYyFG
+H94iWQGzvdsoG+wfTvgLrIP00mEO7seGtvl8AzkBYh8RqaWDjrxycZi0wC5s7fp67m8qVqS1ciq
y5Lnrr+W5mJBc3cMML04sYJDuu0O09S8uwQg4Vm4fKeP9oLER6ujGNgzeCWmkXo/uCexHC5mlwGl
GRMAh57tS+jTKW63XRuoJCUWJ6CJVKhXvyTrN3ZxamZ+yzStXlQ2n2CULQ0+3FYb8Vt3ppWy/uD8
/G78DWZD+ZzIdFFlY2+Va0JztjLUeSackKUgVOvLwxTwkqDHdo+KDqK2K7hDLnIRNDseCwvOuVtS
9NbJ5BKR8sEAXhky9VEKpuQl6mZV0qszcYWDgE5QABXS1a/v7l6SOF5hHqO6FJUDeXipYuwr9hit
6A1VeOquLW2rd939nDxN73Lq9aYHUrcC3P37XQ9lmr4ReP909RC0K3r2f3sOtUZEbt+vbdKZavoT
N7rKFDPcpRMluEPjKBiB+AiM5r878Z51lfXzh+2kECylBFQJTkJ6+WPU5nTiypXKp4WPTn3/gdCj
I0AytR9NtEupU13286ms9c4q2W70CM+yJjJBKMNeIxBlD7WRTzRQ4ylFR+s0CoaDX9YN3iqOJQ1O
OH3Zo2j4dXZnrp1AVjLFuZoA4C1RUTxdCiYga5joXZTXE/csz9ASnfxYo40VRR92IT0/n2DXcYJF
Hk+fIb9UXsqM657q/sn7uFcQDAt/1nFUlGVXY8q2vYqq77UeqzQ5rqMfY8eZ5N2oMPRWEshqH/tX
Mt1FwIcrlhGeIvA98ZRw4H9c2ep/gLRAeNv6tM8hlLeAPiVbDCRWK1Pj0lQmgwn+B5F/0rCBgQVR
9r8t5O9NAPBWpVtHJTSpLilGlQytpaL3IWuMNr7rjFvDmbE20kGQgkuaX25AtVCult23p92P+EfK
mYYDiOMSTDKVA6LQohnC+j7qJiBs+Zwbh9OkzK6Bph2Fcl5BeWe5gI36YET58hNCo4FMHGsgw0XV
x/xRHHeUXHEDm0lEh7OzvuhjKs6qxEJmn6cf0WoLX4kqfji8n2JRXxDKcAoIrLVrhgvy32JTu5u9
1EONMlzdR2HUV/EDyUJixKUxuQN6ne4QfQgbrTEpJI2jUCYm63652DlFYioblV+uQcc4c1rLV4Se
2auQ8bdyXMwDyCSqo+MZM1r/VwLuKGF/yNjDOGA6AK6yK4DY/Teaqce44mE3bb1mGfVqCNYARbkX
Kj5yv1o3XeMk7T3LZSPjwK4AWatbjwr9ABP+uMlIGZFGfl+gg6vk7aG7xFwfD6TdRa3OtFDPE2bj
ITi45julCzDLdZT6CRj5sMM9RbySAlcMb0ffehyiThCRC2kQtFTyt4kvT5VyFMcJilPkxMXDzvul
lspvr2yKW3HktkC4qHfgoefBDYpp3Wy7+Uv6WgDIJHr5veritR5OxM1x7wQvY1zgGSwOO3hLTEij
cee+rcXRDfyBvIw+Ib5AocgkIRRWSLNvPMGIb6Ek8fdgraBaTIoImxi3o6vjY2PAkhRkU1AKUd2F
bD+lXwYx+c59brGiFcIJM90Bd3nRbzSC1tGnbWaI5gsysUQ37H+30a/7/0EQ9NMMLS7RgrW6UIrK
KAiY55JkD2YzCPq3GhYpHK5tPSeQQlWzgEeQOLCWc8NOd7gauT20A98FD4ZhdPuVV8MtFQyQxjLm
pNKKeUhLVsJOq44qojRQMpnECksPGwL8qUhWagtAGUXMitfrahhGSgEucLLqzi74RdXppHi02hf9
/oI+q1XIlHiwNKXYwGotHjE+a/Ipc5FFJuqj32bGjHciq+RG824dLIdc/FBApAnHmupzl0WgvPbl
s/lqXWefBMIsLs3+1Rgw1ughoTIos70+pS+hg9G153RAl+1DDWOg2eNKZpWOpdqmXu7+Xcwu1dxv
R3Py/M/ycMj3LnjHusifbwKUwE8sBwYt/+yKd2pxoOc6MG92rPWipBM6AhhczPF2IV4kwyxu1vCV
NsGEKRZSNbwe8d9IgIBnz7t04kGj03hAyoVwarQU1iEJQiP5jqXQxwTQOBU1j2P6Tp3QL6Cx0gb0
cS/8PT7PrjavA3GV6+i+rMndtgVo/DV+1OMUMnaL+U2Cdf8KBYw0GTSkNiHpdxu5RXzme/+sZgz4
dRoO3Wt9klZzRjUASZ1nh7Douy2h6cftDCNhvSROop4Ety6x8Lk6to0hHnsdf31LwHIMXpX5TKEf
EyfwSyBeLcqb1KX1leV3r0FxhvZE95mNRF4I6YI6wgUg2tVCSyz46Ji5JSwZRcdYc/8aZjRT+MPN
I/aePj6a0CxJWQ/ffnnp7dt3zyGjD5yVhDvEwCPTINirfys4Y6GC39K3iorL2hON1NbkDVpyRW0T
ePjP5v5D1Gm5NaI62hbQFNMk2VrQg3ffnjly3O/KTzsJrWM91YQLEhKqHBWUb4f/sgnDzgeU5pgU
O5v6rv8Z2gH+ZWa9UNs/GzQM0oNH4ZzCivw671mznG6ioN2GEL5YteXxr/L3abwJFRKnTif5VwvW
5LyrxiCiQyafF0tGNQikW+2KCHGbMHkHE1GyYvA8BrSPmAS48ugmnH47H77c/T//GrzpfEeD68yW
LieLl832kliANVyDRsjlTuGaV9Z3gwB9eyF3tbiC4JrD8DopJcC7NbxX7o5Gt5H92Xg/4tCGm0YX
L8SRl8py+ZKxWO5oKlJBrscQJ22y6AQcswWUaL1HwGZ4PFEEpkKEcxes6B+AXV5wAKc7MIfQ1zND
r4oo1toJtj0VLx+176QWQjsVg3rcCWJ0XHE4gaLlk0GcqVfYrnQ5CXJBE2f5qWvHNGiUDL0IErwT
klFAeHPheyILM9PqHA6EV3DGB6f+T+iaBjZeGRnGCgMa4VMLBrpMILE0lgXs33fWow6DZFFrNuV2
bjpy2XBFJ9auxRNWLfrcyYGCZcnmYyHJom5Da8NcGi6sKWEcd8RWS3ZwTeeBpBdNzhWJJifx7Q3G
bFkSBbM7d4spd+fzWIw5wMsS4WPgXvkgjf581DnUFCyUSHGgLXPTzsAUdx09jcoujfyh4AiEpsaC
wo3zRTXErveeG/6vpAH2who5JcvI1CEMHDdlSbhFZJ4rLUd9oKE5JP7Hh8L/KsWGmXi5e/KQ+FEG
PRwwA8ju8XxVUQIgrxLwDwMLb4lVUa9X+ueym1teHSHpD0nGvNWzX8xQfdOj1uVFSmlihJhMHVci
6P0LJllF+m8XRqtdahXNr7RcaabOjiiUedl7zHUNWYoOJ/BTD/hLM59FO3e6MCot8D/TGCaKk9x7
ceiCyQZmoSoYfRW+TGnoJfTRnvdmjZSycnbfp8l0q5CPjw3e8lmK9Xe+QANgI5xG6ry3/yozq+VR
Jpfhpbr/Fa6BwPJyesMp0klP4sjFTt6KJZ//lLj7hq2STZzj3QYa2TGkDUgHbbqgCfH/6IQGOCFN
IGZa1P+dYPA1TJXVtROTq9xKhbo6WEqzC1ewI8NOgeedx9B8poyZnRtyeqSr8tpQjuSnjo1CtLAs
zab1CT9AkezezMYjmA95D3mfPNxWJwbKVYCZu88ri4ZkiL8AhryB5vewq3fxsjeeOv9egCTsqRam
rxmKueJOM6/8ME0qXfp1N4aOfpso/ylwaJySZGrvzQiHY77rwytjGlxtlS0bjheZ/C8qqEFRttG2
IGiWFVbqx2WyUegNGkNJaBcIFjKVW7aPAmCPeqUw/X0lDbRxkTGOvlpc8M7Oe4cUT/1z1w+sbkCA
Ebr8FeUamSmBl96I3opdBCnt4EZYLkzbYyxLk1h+SHsWhyJwz66q8ExGmqF0Q3FUlx185XnS7bTj
2wLK3n81/IuOXw+97lguguToal69eNEB57EmW7rYopoRZuyE27+S6FS7JmEM2Avh9wC/puWWs92C
Kl3CdBauj9JquIs6zI7UhCus21/+m8L1hlEjNvfXS+euw8NTEYtzt5/Mv5dT0DrU8RuZBVk6RUd8
ym+2DDjZObuDlBI7WguXi6z7z0RPt1evqkahUOUQ9dnCTxupCtZMJxrXrsz6zmfH4QpXHKsTrmC0
AHkJgSkO8xPiD2PGJkG0iikUSgcoWavG4N8BEPA/9CI/Kus2AOdk8bC6J3OB5cJaw7Q2BCav4Bce
5gMdGf/8BEPY/mEQam84PhXBo63m3dkZPhe0+mjSlClNpsg4DLSSlZABlI6v9/uhbRbbTBrM/U3w
KDTbTgcZJnFNva9hrqizqzyoxa7sP3Zadfv0X8Ic+z8JS44dCWk5D0ccCzUsvv3Aly9m54fnpgon
jzXISZNyXTCUdJuOr2uzK6hVJK8SQnU+ZrQU0UxoOuHIxFq0bFWfs8NCA87wdkc522TX8Q10xAao
qy5MBFzAPOHQDO0HdgS5RdZB4vDD8tRy44IKybrK3yzsnDIkua/hbiV/ri3xQfqzjaI49uZ37LU7
umLa2Qy0hB+SI/Mg/iX058NoB7NAp0f2R5cyJ5m2C9+tz6sqVj9g1ReC2/Utdc+Njj6a9vg5u1a5
+V3f0TB4qVXN202tRv/4VP5j56hjGENun2W0duDxMuUKKkU+jk4WAr3yQGFzkf1br0FnoDz2wO2G
9QY7N5DSlpHk/gAXQjeqJSPJ5yayFq5NFz61QzzS8nz6X50vcOJabgn5EduycnXgTM/4YDqEGP1U
qo5zj5SIW4F1mDqN48p8JFN5YwCl6+B2JR5Ncs7l48aZ9ncL+GZfXbFjE1aT22J9/d9TwtJIaZKs
Z86Yf+wPKjSr9MP16WdCnh8gsUnLT/mCh+OEeZ3Xdkheo/aRo4KQfsrL+aPWTGH9mh6w0iespC1P
1hwTwkhPH6xppxfVHF2t3WJVSUQ3d3Mf4stTHtbiGtyHQEGzdwKVXfST5rRV5c1j0NSERQDqzZ5Z
zC12jC54znhnmtpqYl97mcZxGyFT1lv29nEiJrPm8+OqwMDG804iBv2Uwg/8CwFY0EuLSgKKFR8+
gqUtW2E/UyLTCPTaBmLfCkwGfEcSG5buB0nyfwViKJv5l0yxE5/itgWPVtXTFL3VfROlG67XT5J7
xxIFYbx8+iS1jDJbtlHefkahkQ3VFQdREJr8SDMrpljsgFrfjywjg56XNEhFvJaSbBoqS2gmnzAk
CZyyghrtxmUJmtEs6wTXS0sfpD5AlSaLZul0u8zsxj1leFIdubCkAxT4RdfR97iPe1OdFef8AZI4
R1hMzygZxb/WSlCca6oeW7bvNOV74FLBxLZV8xTonTUXRdKwX1XVMLFc7LFX1NI9xXIY0+tqOgsq
4bTxwAa7b0+fel0xjSHyLI6vnDPBGaSzN/5j6aDwR1fKHJW6cAP9HtJWsV/T/7gc/pkIk/xWpcn/
KVlag11p8mtLxoFQIAHlo26KWP7BtgKiG/TXdGQ8xn2wcJyimLUxdAllC+uG1l8Nm4hGN+1YPl75
Fcstqxln8e3rDnHMuUL6I/a4EjxvKYRNotpVR5ghE+Mew7cccCLSOmOvY1JOe3gbozjTCMAF5rbR
KLLE1ZaB/5ajp7jrl5px7LMFO9cU8j7+huTFqidZfYvSt/DQ7RwK1iXt/RIivQvZnLTH1jsJS7ML
ghXjWkcZwmRwDYfUk5KXmxraRvW/B8NfUFTQ6xKQLw6Vp/rAwgPngB5d/gprTGRdGCdQqzIfRtgg
HG6TeZY77fjEwfHKsYF4V5aw1tU+ynDHxsXQ8+5bta3QsN2AqLLttaGAyaXXmsem9xkUrsm91MlP
2IYIH+6AyTuqovE9Vh53wpKQfi8tLDc6kccdEc9NvxFR3bybLwmZk/7vc15Y31HyHUTVeyGDCX4Y
tmLOomCjSVy3F8YMD1/Q3n3jSbM1YLk/tlEqUp4dE47yhKVaxk5OxLJweAT0YzubZl606THZ92iV
K/4OhA220oV1G0AbPXph6Q+ZrvVmf6Esa0YMH1dfx81S3YHgM/iAAnWoYxWm7eKpBaGgBQ1j5RCX
alIeoun5RmhMUdpnA4h0iM2KMNmP2qVVxmrCOH4X+ZQHfewRxahlvT33SHN3ON/JlOZ5GPwEftqD
o4K2GJ/nDqjg83EUpD0QOkvuIAEph+sk+QjE8o7kCb03XBgMUbvloS/ah9kWc/NJNBsch2kV+IUR
iquf30h6AMpLBB92FQrOL4+yJu/pYk3IZZw2a6b3IR16dHqRcjwBv8Fe46RN82VogJav4AU0NLwo
/BbN2iGOpM+NqbDqK2HcnjGBW+DO5BQStXA19iA4N6/j0DoE/0V4/bJljyev64LbJy7b/ZcfRpJl
eG1tB5xvgsfGVQ6YYS8X4Ua7ef+p4thfwvs+neRIYu/qzm+8FFpqBwFwjTSwwk96GlM84zEBekqL
z24DjxE9W+gvA16042JtWu1PuQIQoF1esigu8cvrrdCp4hbs6cezRePAjnOXxjXyS+tG7wwnZxcL
eR+AzSdR51jfId58xTdUmMW8mvBuuO6IoGc284cQz8ncCfZ/EOvmDmgCgsgQVnjiVehDovFE11vL
lhF7Kk/xx3tXGxKm4R6tc/KDHsv9ziBgUb4pgDk1Cc1S/yU1Cr1Ao2kEfM0enmSh8ewjNWWi3QkU
VbaXl+20Bb2E/3oNWHppuNkbjOVYaAvuBNuTig53j8ticxxuJfs+4ruX9HWjve9bgG/hj+jRW0H6
3gkluOBPuWLAcxLc74Y3AkjOGi3CRltMUabh7dzf4nnHkuQ9HTBkD+NhBVlKwfJISLt/QvuYQS0Z
hf0GSgW11cxnyKo2szaKFXA8H3I2yr/H+hGbIlEptBkVQI4JJ6OeCa0mXrAV39sPrlCHvAdSIs10
GjBRv/phglxUUAO0gZgw6+RmE4KWrzRdDrCgncaWWEXmsD/c7zOzNT9pn5ttBE0zhtRftg73var6
9JbV4kAFXzibJbsQiXY6WkRaaOe7GM9nKbzCNCyszvCOCc4Guot6BeqPeDqRB7E1GT+l7dYii+32
Ij4BeDSVSdsnGPhVakzhXVoIbpkrMcHED20SsOQxsTzPZmJU+R8x0q/H0Jdev8KUI17Pqjcj9KS8
TVI59B3BUmQR0R9vxHYiWN2dFU44rt6AglOIWPk3VZFK7JBfBGJtiFTYCeeKb1AH/7VpKPbSWHMt
A6YR6M9SZH1lI4Q6Sv1eUnxhDIiyIXMSWtNKxxn5/Kh/mLlYhwlZr/ye/8h8qbZSYzoZtgsA13Ai
RRywgHtSbKWAdtK+QTX41L4A2ZDSd+ggxLizqVrLH7WK0AyQ5bZKlp8vRwmruh9nxmi99Zluzrx+
d1QX+PyC9+FJId/lcO9o++bVzBK9BzYyA/mR7pg+wzAO+piLZ+wotKjWjjcpP77izHaqL93n84+K
kNlbpnItypxOkklk4GHQgj9pBJ+gVbn7iP59KXyWoDbW6FYIB+EsTQ/FXtDgyW8n9MzZ7z3fwHN2
AvHULZYETXJTo4egorQia4CfDR0MVEW9FzQkIou8JztNOj7zbrTmAlIzCcjWYdbZM99ZJu8BvjPO
SUt49dKdWdvT/F7SOywvNUQDvKzeaLV7iqykwWQL0wNAyw3bM3IZGzmlUPWkj79uqR2QLxqqIwL+
lzboA2d1Xp2saVTljVjBVggPLHQXuxLFJMXziPJR/8SivZDKRX/okVFKJRt4E5rq4Y58z0DsHNXQ
1ZdWNmcmcH2Rpb8vhu0t+Qy9Z3eDXks6ezpK16RRY0CCk7sM1MqwrWP3yrz9Ydry5Ka7r8A705ul
Ze2xOC194EFdS8kengZdZoyS4+24yCS34gxP0qOfaoq2w3TIhq6xG/tnvBYvB5ua7kfoQlffP0xV
W0uR+TsIxNGmR+2SKOfJNfZORH55QXQRpdWo+8vmE9JAJcJuhwU44RKsFqjHlJ/HDvshFaeVjDoq
yLpNbeJmARacdl4hOH/G96A/AePuBHpuhEPouTkpzkqOi368oQEL1DJAzEPLAMbvpudQR1SVslon
8G/3B3EKvs3idJSNDFeaXBzYsjWIwWq34RSasP1zjff7YEeYLoARtG7wqYMci0/ovUbSXVd8OPub
l94p/9Q1287spssOAPRo2YMLoNX2dGf8ccPmIuWepHkgKakvADHEwvQAqGTQCZih6lKxufjRUTjT
G39H44vmdz/ouiPzlerXYSXVDPQ5Ps8RkZt/0Yr/GB6PAEA94EGUJ1knfnAGF+4yevnE3oPaJpB6
6rNE9ajVwRYzAdbqftOd4bT6Zy2Rrs1JCWuhtKfYRUSdXi8my1e1KQXYBE/SF63mzsEgIyyUmwVi
eroIiUUt3qUEEHFVhb+OtUr4FY7tFMYnVGaP8YxP3talADndtRy7yEEUwEqyh+UraZqS0CdK/0BM
t6/Cpvrsw1E9wMYt+0CN2wrxJOafIzSsJrQvt2QClx3KkyFY77ifQCTzxQaJOw0yBbyNUVclsK0W
rSEweM9b+EwuYwj8nwYjNh0rdQt94ppVL7YaLAXsg65HIXy62+T1+KQnpzLiDuvgpWqQbrloRrdM
/5qTqOEdYHiKnJ9zldL9N+L3SRnqDx9KY8VJkJ5pRwVj89J5qp0okzR58vdYe+B68h8n7L1fFN/x
M3vZyNn1i6nMhehJrGiwnK8BmiloFNlPLzknOyfvt7BvRUgN1cozvqjtPf6CqXzXqnOpvQhgGf1H
htr7akkkiBXXhXR1x8sTGgyjqXBpyQ2oBbV/PvZiSjFzVGqNfOOh594rq6fPHLrfNMFNXg/2WA85
FXQ6RQ8aJv7f2mTSEf9IJ9RlkovefRRpb317HQlOsYOkOhiozD/53HdSJiTI09jhCOKZTELt7GKP
zFGP8kT65jFk+q4sIysv4yHLcz558fX3daub5aU2pWA2usGDSnmIAQdPDmVMSTz6yqwv2XmvY4Me
z0Fodglc+U95/D+QxYroUjEExiUmXKy/SfmI86T2zcxj5c06KhB6UNSQt4RI4umA5xw9x9KvNUke
QAUmSliO51VSa3dpqbpiIomd+7WS/VkWkUTT18/NGj5dpFGoQNvouNb2t72LR4A6l0CTtFCC7WFx
nxw5nc43bKvCEikT+ciD+cshajWcPIDkgd/ALz78vnxDrgL067rstj+r+FHTcy83y0o6CniRbD7Q
JlKKxv0G5QUh4kfnmzw7fKZUAz6UngGKVX4SiSxxomhwt1dWa6W6+Id5s31KdIKcWij0+ulN8LIz
rBEiQ0IrRYeeRePDv9RuixqRsQl5LC67fIdVVmlPRFyvwGBlGth1x26dWtl2NvClj2IUC79Dx3lC
s20x5gyp3lftUoLnQELZ7G/ljbyYprjS/JO21MyXtUqdCU1BdPV6X7A1czY96FSbLog3yx1fwidg
yP0hYMe4ZlGJaajFU3s4IUBf6w1PHc/wNq4TCVvWLum8wwXzBdoIthjNpD6keRTU99ZOmd+Ek8QS
DDoliwMz9aDodo27e2Aa75qCXELyCxt8R/EXSVKZNtyw4vCEpxUZV3EnmsD740QPz7kMHk0AjlA9
pwKyGoiBSfsUGuGGFhZUSdvTQn2V0VYMJwArh1VIZkUJZBkZcDlkWoRN37AsUIcFbLeY/YnJEvIz
Q5nLj7LVtifJ0amGDGux/bLM8xmdmAanXwTPMvutxmuYn1CalAdmRWTsjo+xvFpRl6bNbrCooeBA
v02K6gk2Rne7Dm6qSpfh9JtC5KTLx8gK18pYd9E6wwjhWYsBNubDATipDaWDJKkZW0oHYvZu9heM
LfM7M0veV+7ou5RLd46IsCKJ2J2Hvu4QYyTu3kjMoO5iiYM+Q60Mxti2hwIyKeiTKW8j/ODH8i25
OIKrQIqws3dK6jFtEpb/gcvfZvCrzmOqwVaix8xqXW4qEfcpRJKLB5fYzAZ78hOF+Tm8Ye1pfeKZ
+ywj4A+Bxf74kO1JjmLuku9q/pHP4OwvvrcxbmeFOOSg1/9kLxJW3GWF9sJRVW6dWyTZ1pIjoNDf
upuKrvFVQbAn6M2lZuZIeC8M9nDYGBcB/SziXwlgtnGbo56ySkkLOgX8ynf5KQ4fPDuTRVuVQOec
HwFWiFC3U0f/YlZFOzD6vkaZmRJ624EO9h5Cg0RDcVjPD3EQdfrUGUV1bFgxtHu+Ju+xVKbNTU/7
a/D985QUxx0ERuTU+0aB6LOBGxJhoNFJrAH1YxiQZ0ICdHVnXNbDmgea+J9/YdKmp5kYQHAntxuw
ewy6UHJUtQcHbymeWN9BdxAG29nySXXPxM1RcYYtbp/YhdrSB0Tv9QjPuJmY0t7/zuXJIwj2o1z+
Cl0NKbxRewFMi7qDPZbZ21I5BysEINQVqIw+AbOD1Nrd03Fke1YZRxREeiv9TbvTPw4xHeEqd3E4
rIhOT/HtDwo6p1/rb2tSPHeIkWcaW1DrCqkiJ6TuV4Bo1k6iRV1BI2U3u77ZoOs47LogaDRxWndO
VscgdwgM+lmW1iJP3Uu5mKeMvzwZxMeqjwgTmXs7ntsmQ+kieGwnJyCfQtOGoi2cphgn3SBaDSU6
oDpeGcbK3to5dE+GzCOvyfZlqacZM+hpgfPjOBbECVxS0MKGbxpkViUKom4XwcgAAKzA8fe0YjwQ
AO4CFBIDJYHZqukJhtC35mxeVHZzjTUXeLJE9djhjU20Qvb/IKuGuIDr0TncEBHUBQh85N9yXJH4
fZn2zASHFC0P2GnBSPl9C07clWmjoKOyS5n8veyVE3roITTfnpnh5kk/p/Z5wjeDhvzDmZsfD7yR
d1qyRFrmtvLVk97sQvXcLjQENUPZ2w+byFLF5x1LsqDrsGFsq1tdJlXbZLocOI1QifxeJiyaLxm9
DkhvD8H7Tn9GyCpbrS3tFbM0LDzs14G5agzkVAGDTU58asbtVPw2KwJcOnm1Cz4RAgak9ZyfXJTA
spJVR16gRjGZ78rwb2NFo8RIOp3wdYr+FWnduECRqBgm1aFaVYsgVnPlITKmsP9FNlzLyVJfgWCB
CFWCh5PI2qHXF0lHOdPQk+1+OnC2SIIyrUnqcOJ6gB0E6UcEjOy1SZq07Ot3wdLSIdoBlg3ZD1Oi
suPdD1j1SWL1VLXrPc8zU5g0SxgWjT241qEYdFrsN68LO+MzJjCOllnKq4bpXJ47uQAVpJPqyh8f
WWcO9ECnFtDWA4T6JpdukrusY3QLTJg7X0TFQXUXArF2cx/zom40srVDUg86ERMO4su7oEzFZ+T5
PP4W5KR1COZtvppZL6Y2SeWqPqEQM0eUcCLLPbRdYywy1lPYC2pusmFTuvuaVKeWXTroWWtisPaD
w+GtFjcca4fzm4U4Zt3CB1xKHBpPWC6u/yQxwTHsJsC6G0TpUXu0OQmyw1zu9YlBc5zqGIiuxDLD
8bwMapWPgva7oWbtFsc+09gjPdPI9wMNB9Q+4MrBuFxC0eyeCGuSDghwe+8/EaOPUiOKHWSAmYV/
XpUXJe9Pj++R4GyaF0ECL15WOj/eH0zEwgZH+rS1ErYKuUE2/uI7uqZiTYWKe9T9rIkK2Lr3gYYD
+8ejCwVHis0hMbAgwzp3QJgArgJ8un+pFte5gtD+9QG952w7c4ABLukS24D0vbczNplcWqFiryRB
XlKiO1MaRLoX5XUi3fkiSo4W8S2owFKUbIEQ8KVBNdhUqeQCRXjJZ8zd6kAC8PfYu9el4KdbWgu3
TPSX5v3XgV4J1ukh9nfsRxbCIsYKhw5Pc8qaigIkgC4WstpeQPb+5oPPCBZyCs97DzFQlZUlrq1X
0+i+cnJom2AzffQHMSE6Ad8He3u7cNOObvSsFWf+qSoRcO1vJ7I+0mFuzdYh/O66Ff2hqT5B1hzZ
OLdkG/wEOou06rkX/ozeDiSpLMr5nLULQupb77+lN0aXMnLkktBT4ij8ILHAsTrso41SsR9+WGHr
jdgZROVB9rNkB43seYh/9QYyzIN9MrWNEdxHA2LcQ/Tn59+oirNwYMxlzBSkGXa4KOwmCnp+lM4S
R7nAhW6XUAWhBltXT11lQEktFbPA00PhT3svzXBTb/1WG+E6jFuS4PexVgfMHxkZqq84Q/q7Zstg
fB7u1MDjt6fo7rdtNe8sZQkrF4mtwUY43OGi+/BcVScH9YayB9sy+7U/Uk8zrTO2X4X+ZIqUH2oZ
X95Y2XFL6J/UOy8c6muJF9zo65SwieoEQ3LA/QvWfdsld4O1YeqvtPSCcYa0aZ0XsbMfqCGeEp2J
W1QpTo+R9/qMxWRkIRrM5x8Z2yJikN90dEXBSbF2kAmq5azc7IS/tuNejfXKO+s9M0cbWpk7f7v3
6izPw+ubskEmVDjQEVS1vavn+BmWaHxsApRJ3rOxAMeSTLPZu1sINuPlOfkH5LaVglvziLSCn6jF
xIOWyCZfDWacM2EX03K5cOxg1pag76g8geL9o8i7swYobfnmB/RNYIGpAdUcjeXJemJpfkj/uX19
WYZCJBMMwK2kRfSqVNzd9Nl0pVDefcCOpH0Nm/Yyes4kh13jqVhI4BXkEZmsSLsd2EGl+CJqrYVz
7fQ9yqznRrsk8ZANwCffOkd1r531Rdi4dzvKYXB/OPzxCYtgrbcnkQpKput9Yv45YoDZ1CT4oJpn
Vk88OkUVOdmT6GYBAFJqcg1+frkkdZDNTqzyvdjBiZmOwj5Zx2aE3kQU8yz6W5pZdjZy8GnxlrVN
tsX7i1nwCWWpxqWl7XdjSu/Q0oKYjFl88AxlthCDwRfemcGFtn+0IA+Rskm2AOjQXUGGgIR/4vop
aNIOA6432s9nxCUreezvy/vyz6kGfOxxxT2xkyu/S0BGz+ubu8GjqJ4Hy5MhXcbQu/R2f9QdIalF
KLrpL9PFuunBqjzFCVRHn5DrMZtZBCCUYUMuoR7fXeGvnSFXzTgy2SJy2d9F60nV9xivE5sIzYW3
4N8Yu5aLxer1OV76NxAntDY7uv8IvT3H+1838T0Iub2Z36jF89yHhndHeawbp5/pWszYPFGTmeVS
W4NBQhIqcjDZZovpW//kJIois532novRehDPwZucjtJAENoc1y8BNieJfmX7wTDLykXru4vtRK0T
tt6lTyxAreVpAACWPhsMckMMwdxLiAQTeckVLAM59ozoBOIopnmTBtjvrOTIuaEv5+aQpjEc4UVf
qWCuA6H47fNvQKUzWlRn8ec2GCdLeiBC6feIBEkuGbWrSDp+Pu8OZqLVpeVGHcHo3OtbH03ccTEb
zVdDlkCEtNBXAJ0ns/5xpa7+BmGDgxfwpfbuYmqGzg+uoIvNrmSAhS+nXcK3mR2wLL3UW/y3Ijed
8sMndLhQG3PC1DFBRkihuhavZsFA9i0t8k5PUW7VWInAvOcWjbmIfPKtjb2vaMnoZqQTiXp9Vu1K
1fKRXJjj0vatYa4aL8zCgtxh0sckOfN1jfF9CVg6UOmMiYDv4gdlqBWm3+UigCfFx0VT7fWoCxFc
nqX0PG5+lQLfaHOvWftPYP8j8qySyQeJoZnxxM+ro/nir1E7wU1OvaP5chC/C468K/pUsxCXT9nw
6KfOl1E67bNJ+dRqgilSJMLYLfcSqcXPrG2owwAvtb/SJ8voKFk1At+KG2z8T3IxLEQIzjAR5tvp
Su7l5ifqY9jFcOnyAXl5e4Gv16LyKlGix6GLjlaEVtgdtoICuBxsiLA/1AYEVzxZ+S/OoOC7y3xX
9VCRIB21wvcxv367FWIsW4gsTuHIa+LpDRT9F/KRh3+KtMklBPqFovz0pZnijoRF2bK5QiYCf28D
JtZu2fk80T8ZprogCbwgfuCqM4Qvj2YjKVhg+iyG7ArdM9+wKlE2sV8P58BemqQKyhU6UWo1cram
ZQ0O6PZR3mD42VP8Mxo3YaWYMv1Wfjdqsw+Fneoovmp29IIfYQDLtrwobv6NDXLEOotsqXSjjm6O
PB8lxkNEGuJOsiOFJh0VSl2+xTLVv7NSLQVwEAz9hVQNxPPgq1GNOLbV09WZK9AzRtbSX0fqh7AS
G9Md6r2zZtayxAB3fUCAdU9zN3dOYUeCiaGOBc7O0KOegqmozIl9L0nHz5FZl/Q65i92+/0uZZTv
UbhryemDEREpSGTjxQ/QIX+s89llyIzqR0Vh4+aQgZcwQmOyAdswyawGv14brAMzVoykjp1cpm1b
NChSwUaoYr/3JdFbRMeGq6Z8wWzbbEKc2WfyvwedSjzlZHTQju9vaC+9LV7Oo+hOidRlF3JBxZDH
Q2FZHdL9LUcO7DBksp1Dst9YzX9oUXbxEhv9BtAgM05iTIlxmNxxPvBR0ZDxJu7GbXk073LJm2hJ
yPgPwYgTV5qc5gfDlCb9g5R8NOaxhuOiUsbvvp0X2lVoeVmxI2idIjfSCDrDw24J0Q7K2h2gkhR2
iAwRKMoK4PTkw+GX/H+FpJv+nsucwLfHaQTqvDZJk8wzKc8bluxnlC+aTLA/kLZAlyaamLsqwomG
Bgev2NZL2rdeZZjnW2j51XX/aHfcaMD4VkIcHMHLRVkmS9UTb1Va4V19I7UCHcd/LBVkVjj4WFYg
TzCC2vzxeA4ns7WazAuVsKs2TN5EKrTlRZxj7HGxPtJ5E4KltPv+tbDE8l1cQelbCpQDPV3dZnJq
xh+zjvRY/QveQ5g6OZgfhT+1C6HDeqs74u3+QLg7bYZPp+aawjiiDvpk/9u/4U7cuo2M2Ck6valS
eqbOxZENU1t3zsqGZXZFoX5Sicmfug80NSRsnAx5A083diW7e7QMcCYlIyFn57ObTpZJ3HndB/A5
QRrIZTvnnNUXGSm4jKKhKes4SenaoeARRL+TY8fl5QzgeZKWMG2x4lQe3BJBhamtJuiyE9eU0nVR
W5J7L2YdiOk6D2POa9cIkE09mwnImjGgHIZff8dHMM0SKSFpO+yQVPGW2K+3O1x2sz5nsVgngzLX
ciNagVD/f8bQxoB2L07wSxmBu6WhIO4vbA9KX0c1+xLYZ/JZ4hO5jawzf2f3EclzvSBFfNQBmEip
TtbQHafjo4LGXpT7lRsOxFxwV0KT+PbZMOCm/g4hwxg4eGowccVv8vLIJe+dl0cnBrwQnc6LDDrT
OURpY77jR1bzM9khTL7RR1VNT8kHKKfiN3R5O0fjKI3BsR0m+vTneqeuiR7KxouXHvop9EnUMyld
1aazlQ/IVb2YXMcCGEfF2M2ioGhLzi9ekB2JB320S5ZjHk1lcsOU/yOJKEA8DZ0xvtlE+DodcrQD
QzS0Lfr+S5kVcCIyD4sLsfXlfQGHpBJMxErwaeKtoHPK70P7VPttMRN9lt5zO0IEUwhQ/ISglzj0
nVZnQrSC9mbhiDDHn28eQmL2qtZGup3BFWTjZ95iyPvQTUDDWbbpCGu9006YKCKaDgRaDRYCm7Hk
VpDjtinNu4CuhMXhL3dJmmGkVFRJsRDbpHilGYJnUAdSC+BabVdkMpAmn2yON6QlU5MSkDIHpqVf
fFqvhfQWIjjBejJ7Q7lg1nRFKIrA+WHxuPuXkx/zZCAuRVxesu2XC06F+lZx291PrXpYZEoIUDdX
A4b+ncR5nBA7kv2dGK3Hx8LEYMcLw9nZ9JXdUquanCkkpq1YU075Ib30PzKxpiMJQ9WdVPwriGEZ
G9sBOdU7KB98B6sFYrNat1fzGH3qoMjxkCdrFDElhNhd5w82og0cC1NPUS7cY95KTxn4XSZtdO3L
bC+wCx2q9myXNwcpPsjuSldgGpmS5aoWwd8DlvOxEDMt5nmwkDkz5a7ULa/s6og7oL8+vC8IZddu
4JRvaHmHn6uQm5sixsl0L0I6fePoL+joEunBjqYOaRK6/Gzk7F+OvaUmYZCDwAINTD4x4PxYTHfp
XkV7HaJ3ngNl/SA202PgQ7F4oaDL1YsAkbkxXapDlDNPmgTLXEBQ6eGYAFB6rdC+cT2f+AtrQr9A
EKqhQgNAYaZNb0ZT8DC6Nf/envsNST77WcpMKvNpC/hjWLdKOP2oUYVGPCc/fmcP7TYoIzZisSf4
P1JiTCuV5XTyfJmuiF9M52+4JG4Xi0fnecsBEJ/BYRvzlCR+ZXKyNh0NFCDUKM8MUFdVinXiU0BS
r0gRd561gZT5ycwDhut4LBgmJbUqnHPLVd50dLtPqiNmh74+rmT8nFbpm7LB9yPGThvVDr858QN7
svLbQk3AN5fyyM5U1rTHB3g31zTdiZrIeTpNMWi3b3EiMdyq66Cj0ZaTkM59c5+RX1KdaMvSoUmH
xUEKVV92Dc2B+ZoiKB/167fIEJww5gSEPzOLlfZMemJfMhSbxtqUrRFh5ViKRnvYuIPjb+i4MZ6m
KRfW2BdboH+QVOoxsKXWjpkXiF3GlRcihuSX03QEEudMflGwDUUKm6Yq9N4gz4OGW0GxJz1T9ID0
smh3GSQbZKwBxhmnJiaD1Ly3tDl/2tXxczIWQqS/23rof2qzD6jL/VpbE0lF8Yt8h3X08x0IQn35
eeAgZURUXl8rKsQQvJz0xtAvcJjYUlezHS8FeB8m7uypzYQGvSIu8c0M8/eliPwYesc30YDNXK70
yqJCtflSPu2WYWV3mlQRh3Ye/7CCdXKl1zChb2hp3ION7bnbKlyqRmF+y7JP6o60hXr3FWfoFmPk
fKKPHQ+wTSCYBgbCVxuYKDkYFRPxSaNaY3VIPmZALG38rGnZx7H4QpRBmYdZ52LjvjgBu7enbkrD
7m4ASKW4zuCRIorRsKbwIFXIPFbsxGGrEf5y33vImMKx5jMnIUGUU0/31eTtCt7rTrwUlQcLWolv
fmEZ0ZLy3Isau0aG8qlyiFDXiquuW5xYwHFvVz1OwjRp6VVLwusuee96kJYHXzeM1VOY3WmIB7mc
6y3bbj4nYB9h6pmORkXMx6f85rqOG4LOtY4lD0M8jWg+iW/QaU1cNmihAnFyEZkUDxlUGF1quhW4
IQkpesR8Ck1V5XZ2Nee6oOvmtJ3JRzbboxdmpjqsr1gIthTN4n865Hd2thqJBdWgaVQMNH7K9zVz
++VpEpQxavAMakSe70qoYLrC8SIqirCCmKviv7hsZlBZrCT2lVUI8i14X+eweTrblw1be3o3dGVX
wibwr2ltuIXSzUmzCRv0I87NlZn1alcqK4VTbQ4hVLLVmbtTtSbe1CoCTUp4U2RLxhtV1CF5SfE5
qFTLZSxH/j+63CRnzeD1cz81cjh1QEP9YQvoXMU89imgB2ygXfPdHRT96e4dUzenme90/G1gXTyk
CVpuwB2gb2Jxh8HjtcqFPhxR+0hLsTeuSJMo7v4moSZQrNEsFqLpqqJDgHDUz2GXCVGWajPfg0UU
+84tFOwsuUzbFup7/RkYR0Ps2pWN6dbO5YSet8d1iI7CRGqHCe6F9uGM3+pe2xfpM0yU4L/3IMhX
jpWav8b7/ZtDGLqjtIjJ/Snj2Lm4ksQ+Mw5jldS2UhZ7BydhOplpEgEXxbI4eZWuHx7BYaAD1HsF
CUpW7hUM0LWayf4gQUOplZvAznmjvT5dr07Zc5k8UNkD36XHLs22yznkPthdC75J+bmXmn/pszNu
5DZ73AOgFco6ZF23fShpDJpeyUklgVMnNqOL2LCZ2MF0vcVrkfyHV+N8ScaQUy4uNSqxid31O23e
qAsukEOZfgdTNqPPmvRG7uCOGioWjS/WN6IpPUgGAYVnQSnwMovYffTbT6oIKf9m8QVTdaptJCuU
9F1IKN6/O0/gMxEoIgXneRjq/5i9/ETXa/to5vVIChBDs7Gt7hJTorF0JZEEsCYOc8H4bK5p1NXa
Ffq0IXWvBUrsA/OND/eqosaMS42K15gnWgVWcGvgc5h+ITT30F00t1cYBxNeVcM0qdaJGl3ckIPs
+cbWdZRgCQPsaqqsilCEOby7ks9Z8Q4l+d957MVtLdt64rOE6UduZx3jm6aJKCIbLWz3x8AxdJ9k
R/IR1R1rNfKz6pJF9VJFQU0pl1GIXoNrq/HL5Zqiz2YBjaG0whfZSeL9sm6gWNP5/gfaDugqfSlS
+CwwBjSuS4Gd6BgWNOGk84BEIZz6Tw7y2Un/RvINU/X5SiBZD+Sy4z4mUhxsACVBYeMku/uTM4oq
nj4k9621PH5oEqe2FGc8BWGFTkWYz4GvHRkKkp/9v4oOqWXA/9FCiVxVniBRiA4O/0D0SMxDWN4o
nZCLO/MoS9PzUnsOiZ7deWJ9toekLo7akInO37ryOmoggNnaJFEyC5+muQFr+pHcLu8RPF6YWiGk
L3nF6pnAMTy27CGN3Jlgd0JMkIhW2LutuHD4jP1NuCwhMq4c+/9dzcBcSxfOerBMQzDUXDK3u2M7
Ue8CMRqauiaeyJAVnDEE2vRZMC97VYtxEirbPcICmp8JD7isyhJ8wl8zwkA7VU1eBiF3mb+F+J6a
Pcmgwia2KOb7POfLVLoz/ZU6pwoM4X1dTQcWFdc9umo3j21uvUL49Cn1QDvUL5AKoP6ZMj9Zl7IP
PlZN5ux3NYez79H0PsU/gSRlcI/Kib8uka0QJiO4DIUqQvzbOgI92ZLAFIqqxbPRu15F7FNAW6Jr
WwNztvrVpE1bJJCYdTSDFI+QCkkyiR5HTr6x33/mn1bYlALf2FrJaBrWLM0OxrKV5HiQBn5g3Jic
zGzQb6aipZvtFKbYDv94WOK2WTihkgW2q/n79pzXWuJeq8Indyb5hVy83q1zaaAxNvnBpW3fMqL6
PICZHSmXa4T8b1p3tFK51Q+fZd9XuIZ+OrJp8RKcfdiM2FDqqg+Dr3T8jj9iG4Cme2dX9EbhGSEK
Aq+S+CYOtQP8fwe4qebfJToRSDI5TuxpWWa9UcoOItywV5ergqwad7QvN9oig2C9fYo1U+ColHgO
Rd00jeSRTK51W+7Vw7EFFrek1CBAFah1GCwiLuKVmYxGeJaEQiXnxdKEpOH6uNibK/Jv4+oJLhMA
0LAmdWIIjP5r5UXSAdBuKz8KBun/W4xqWaqyPwHR3WDaDYexH5Fh4n2DezmVYQju5rX1PwwQSW6n
m4roPKQlZJd8H+WZzeNzcq8cks8cD1SGgqffBDWTVkKmiklpdAaN69Fy6RAIsCWkK+fSFTUDOU+1
GERJRO9zqEz8QEHtyYpnHuVupPPf2sQbKd9i7KRvPu80izdk+/TyiP1zbTsBUvx+T4maUakrO5qJ
U5eLUZ/wI1IsSV47Vu8HfNsIcIjS6vRA8zfAda610qoCIh9dIXW80tf2OqLFKX17Dmc93LHSCtCU
oOw/MImKXvDQGi0WpR5TJjQmlBkGALEnAxcADzVLxy5oaGtPNFzJgjVgIvvAiJx+0uxjPAkzgtwO
uWhUq2WhWjHpIiV70lpjQlC0b6rXs+XOFTl2IqDs+p9g+MF8s+aJXLgkps0Uuj5T26I9Imc9YvJr
EmCKDQh4JGR0hytP5tUUtlXj9BUnSOo+gCxow5XMIx0dqjZQlerH6eiQ3RE8BHJwK+UqOUmFVNi/
yUAn3mX9UrDkty3RLEyhEvcxJm2uvIv3acR559EZ51nZ4i9wlb4e2txgMQMN+A3rrHkvRoKypp6j
+LocT3nAr7T++FhVCesy0TvflSwRD+7/NwX1UT+9LhPSNNinP6cpuVYzwkO2EQ5a/8tiE7ut3wWB
W1wvJzrru1KtFxk7zbBvZOirged3OtuFNCpjXBw0IEYWX7YDYEGy3TATRNM7dWXJlxmZXTVAsSuu
YOb+TJgTTgfRP9teBwp+sRTeWtlWI0z50um1eTqccGlU3sZ0LbWH+0O2wUfbcjxJZIff7dTX3cYz
Hx2g0hqYWBa8Zu6IGQLhhYDw5LJAHVWrPU9NdSupDNPgyMOloL1C/2BjJpUtxFz/aqpUpHvfsgZH
w1/79zmICUGiTvhLBALh2HlxB+mrcDQvNAzUpjuihc/cYFdYNK7o0wtmPaa1UoKFJyhnkYLcqhdd
Hr3jO7wgEqN7EgffXSy8kKrcOIy5oR5deBtIZgB9FeZZAsfWhddSeWVdsVlBJQGEAA89Lfm8ZGNW
NBpPJwSKYiDWomliau/LrA12GPYxcdZRp1U7B2590r2FLsP3Cfyrnq8SFGag7YgivdmwkXu8JkWC
9WqeQMUtiwi4EMF0zU9WG94HRdFfZgtYav9+V7/4NXq65IkWR6VXr1hBHwvymDZsqp4Pc8gcnTfO
YkLm9+EKNgQ9DuWCsq57zH1u7iBMQyUz3dH8cxhDRkwbtTeITor0jDpzYcfqqocSNrHB7zLbdeU0
LlWCx1Hf8nQOsiN5D7GBCqH/VcuxXb5gBFH+DfdBq7leMXM8J/DedLveFHzasSPcnJonapEDzQcS
bB8sA4a2W/h02AfGhgfqrMkoEfbSpDQhmKE96oCSjl18dxPQLkVdiTnkMuKx3Do1ahmhxk+XCkP8
AbcAZMY3w29DDIU9S7z4Aqq/WVEgGsMTdsKQIHdYlbeQfMYVkH9f4jEwFLGP/gDKrrCnp2Jq0ikv
r0ZemH5i0PpAzifuqt2Yd7XBeetORNUSq/8UM8UjZA5tI09CJ6sTSAwC6CgLy506+m7JPOE4TytR
CoSXp4c99mPx2qPhWM3+vlGe0Kv2/15f/7InnJcuEFxh/ep8P1czMOQ8IRHu315+Y+HG9/Atp436
YMP8Xjz+ZqqfohiMWcGgkcZ81ENWdbNCgMajEVG+ItC/Ce2WpOes58hpWhaD5k1bkiXq7Sinnzm9
zzgn+ImcNW1fEKI05QwmoXrmbm4K5uHrZxVh8bTNovlQfC6E71JK6cNNEmYAwZDGFCmjpTO2xRSr
58oTxqHTm3pgWfozwxt5iNTxi1s1Q9elGJVuP5QwckQwECOXQ/PI2DLGYf3NEViVtfLnBkjKVgeQ
2dHHLjFyxfjtMC+vauQ7tAnJzHgsV12SnJf28r7fUuDZXtSJIudgUrm0uugWA3j5mEwo+j0hn1uQ
10cOnxqQUHAg5urnmTKJw8A0U+6LpLSYZ2b4qFNSHZ65mi/xUx8VqSjVtiYAHbcEu0Q/GG/WzGIc
Sg4oyZciYGs3g0hGoIYEXrOCcwy3bpdSzlLOZ4YbFUaVlC4RRZK9i8lWd7jXLra0o2ywh7bW7MZI
PK91TwE5uJjGofcBMQ4My9dnbJCgzA/11Wd+2e6pwOXy4j6qX84HR9THZB6I+nqi6uBmyk4mC3yg
ALUOoVOqwFj9utNHgGHQNPmKqfwOBBw0RDUSZqlBX2t/PHOnEoxXOzKy1g3u8SMScAlN9mSKngGr
9YtDyMF2c2iTrVNBRVIkHi8P45ocxpZKP2Vh9gEoQI9BVd5quGVNKHmTUY+uV0Poq7j/6xV7aC8z
L9flc+zeoJAauf9i0PzU0U1jh4OyGaCquKi5bkFIDTlzdbL/rAPhp1MYGo8HwuoD3kENRPUJpJhl
OviU0WoxGsk/rTUZ4Y59e8gtuzBG9jEBxvRhasrLfs5EG+dDBJH+CNm9Fxvp4rLoCe2+U+CoP6ok
Lm6BFFVjIbpa+PIw9Q4NtKabVPJ/JUegpFDy6UY9TtUC7Jg4HhOB8dkpQnGnlsBXC7uKB0qQwsJO
j3hxfLsxmzr+QG5ozbFgpoL4JcAxpR1jim4c+Uy5xZWa8+LRYW61pifj824/UEARCBhBEuRaAVRP
9dc6p70bm9HbQWeiiIsVNqoYCSfgPlIJu0OTxgrtANrvrMUfAx/oul6heLanr9jDOSJFv0pnQ5Ih
JvPjIcQEtk+4YGos85VwGNt+QjqoWhwotRfGOH5zJf135jo9HrEtjP+Gb3DfA2DOMeTXKD/E1CX8
zVCfM4BdOuEu2L+YgLlH/MxArgDZH7astCijALiEEm9r7CM3TdQnSqnfccZ75QjFCpmZnyK8Xwff
4xEPjkWNI8+5Q3p/TTiItVJ6ZS5xC+0byr7LAPfi5kLMjh4mZKSGUv4LNBI/bKFfWYcrc5JwEYsh
Lp0ULt2akqDYyTKSw+u8apbPQ75dR86+g1F1YzVU5Aznx3M4KMQqzXg6RE17DzbdBB0kSnu3em9T
0K8N31mn1GGOW+F+Fgxc00piKL6s5mFZYiow1Pn1mbCGgILoCQQv1MK/IGSY+2MrZb/0avUWH0sI
5onVcJcTTo7WqWeRBJqqhv3+i8/NNpvybv9VvsZdwaKEDjCklODnJtZo6llKfXgj9WSF3viTPmX3
SsZtrfP+e3ueQJAnmAevLgT6rIovzA7yiekRXGrz0q3mERUJ/yO0LDqVKZsLywYzIiYJNzhLgZ7s
5KNXrk/9KPOYaTXhjgYcSTLS4Zhqiujo/CZWhJ9eA7u94Thw8yoLh1NFn13Va9rhB5T49vbpPF+M
cTaFvMSwYGA9hOWNX7IxUEloN8Ia9EF+eH9gBzUCpHUuQg15lP7Jj3d2PNqF1TDj65qnA8JaNZaU
Tq+UHFWf+G/oUsIqGqaiATzBwCl7HdVohWGopY4+iVVKrpsYS5BwMoalrpDX49wMOLlgFh/xrEfr
6RI6RRTf/dBT67d9iNHpKMI+qn6DGEk3ieHxKdWwEoPgUtuAt5l5qEcMQwAfa0+H6QEqLF2ks5jS
4aBRN9ih/hdA36DDrwrGf4f7QTLPcKCJCCRuxO25sVxoHZyLkGyZm1UQhH9Y3B5Sc5Lt5ueVtz1Q
bGNz4y8AJet1oqPNt4dcoTc70NjNJ0+/fHgAJFf1G6Sd6NC0CYhpvYtweR8Tgqth6DK8UmnAiWDa
0SvINH4NMPzrfpl7vEueCNiPfwyAtAbpY8+uknHvE5VIY6rEsJyp/y1BQxxfOJIV7Yx6o3MPT12f
oRLl+7xRjkUSYIlxrrJ+Dfi1RUWXellGAtThIYFiIsoIqdCWZAMz6eL0FeJwML6OLeBN/bf6Z4YE
HwH5vdd2F9CVqCY8lpU/rcRuOFyAFUuDGGamxcm8OWa6r1+PeuOE7elIBDLJPut0ZDXRrgJiO13W
9oXEL8mWfvsTdXmCsCpST6a62YYzQX11Hy1ZZmytK4S6xEIgok45IEMvMPNYrTLJEwcvxjHQ8ALi
HEnjuTo68NUF9ZYTmQR4vTn2i76vqXD5ZT6OH2K1JrlcddvQuIB354bXqkK3fcYjEr5MjqrI/anp
EuPF3ckX/iJLE3iKKzqI/wqyAQG+sloPm54VvjXsok598A2hdQ4/3WFzRvZWG5rZa8rSLrTJslv4
Y7TYbd4cQU5jU37Fh+oZkyz1VLmiEPiDviuYs3eqUa125nRck/UZh6o82cRY1CQAzhh5Zi2l76va
/RJw4Gi0pbE5mGeuHmz/iH53ZDeUPRaFT/LC2hbe4aCoU4X1EYvvzQ+D0hf6pZ05yOpz491aN1rl
fjQCv4G5Yn1yNyn/1VntW7IxFtsZidM1FzW8uMOzErmQt9afRk/Qp3mnM0oE3Ndk2slhcrBrNtqD
ehDSVcTAbYnfrFmQNnW3wfva7XukfDGdggc1DaOhYRofgjjO3oEpzZiJ+mWdHeaFlgbo1gQIkF5j
Eaud4+o2+9GqfHpM9397qWiqbXRNmehhvoGF2grAF2QrFIJgpOP8i/jWqrKoOwvD2n8SV8RfdHAd
T/QQLEtET6e9dyVH3TdaEHIkAWFxO/APB4FNTf5rfEIB6YHyxDm6mRFSqZTvhrJU1S6DO2gHvT8Q
qG2oFk79HaNC/35wg3eeHd4ICOc+lSymePqTWQCXwQLBUL0yNAMkc9Rz27NqiA01MGIWQWQWEtvU
GSsqDrYbA0KGnARMBV5CEHl2Cf7y0KDk9N1RNXmbTOi7PoyYJ/PPfSXvaVm583L3KPFkYPMI5YAX
zdD9BHBl3hfJsUU+VLWVZ8Z2/S3/9QBmWWqyLvWY/DPOUmXi03d1+lgXpDRWnsQQlh/X7ihEHFiN
PAkN4YPMmHg6pn10U52jOp2Pp5IoOfxUVh5lZXEc5NF808xGsQMd9n4bW5V4ETSb3aewOvCO7cYF
4hfQ9dNd0vG7cSam2fYjnH0t4OoLvW8RPbLCWsNJij0MVYxT05hicBFx6UnBIhFC/E+SSmLsuGgJ
91M0ZH1hG4hvYd8bP1KY+hLR+VlPrbWIu9dq4NCMnWHrcGaV1bNFIddCsPdiQG4blvTvzc/IWgDL
0E08cCf28Fqwi9LhuEACT8eHZVOsmb1QwlsAI8apkLZ89rsRglZcLsI0X/x1l9r8hk06DLzEabPy
ZId3guBZffdq373uHRuEnx5xzrx3xLf+g+hI3LBiKnwrcrVz1yHZuRtat6mWFN4rXNLVnnhXGjnf
j4jEakYANdQDCzLhYVbRKv/BEak9d9R3s9QMgRO8MCZydZ3iq/tt1aFv9HtYSe0QctaotWthcq8L
NrhFlfk0pl3SyoACTB02Flq4sJ7cjWYMsYxyjF0kCJwjDf606IK/UN6/5v25UtfuotP00EJVOhhr
hbo2gPIemRG+p9mfu8oPLX9xs6RCwDyKKZIJIALgLYiuIDS5FLsXaRAAPp8Z5uoCOKGbq/y78WHu
rn5ypvB4Yp/bxJPsFGKsUTToUUHRYJMr+x+FwoshYWzB2daIxXZH5RPdO9B2gdW4KmcTjTBvRQmn
Z6k7FCf8L8chcGddb4e4cdTMDlhN8Jikgq3No2EN1tyuOSByuKM5TclK+kxmaVgF9nXsh9Wlc3ys
C+dSKAtlHjqmb3+zKQY+myo6dY3suoTj2OPJBj7/D0gzhXpZIRFhDAMpeqQj+wVMrzJcfDwrq009
mAH/Vgw8kwPk4G7Ml5ufFLS+qXmaeQX71jtYJcJ0Fv1axBr7u/QYaXfIBkxTA738DNxXO4CN8d0G
EXkcONk74Dyn/DCzYmzz9Qq8lVdPKJ/1chis4E1bCfHphOBDoK/ldQtZIX7vliCnUk7OVCK2dLK5
GT49v03ZhOdscDugx1pyl6XYy0DtfP2kfrwNGdmpm7kYiZfjciQv2t19wHzzKfiWj9FcWePiEFbR
wWxodxvHMrgOrIrpDgKQKjFATAuJy4sQhV/jv5BkNflSuqWkUd9u69WelpfVWIiFrjNA0NWPMON6
faDXISFtIF9tvEbrg4qckQ8Ny0N6WxVmY6P29R1SZkSEarEucjppkIpYfsilciKibJXRrKfn+M9O
i7YpuYQ9qnfbnYZazKybC1ltFo9PstV4wIYTK9ZSGdxSeYQulFAx5omJGCaqNythjTzgGcMaxyFX
EadzEa7wncd7pjXd5tJoX8Fg7bB/OT8LScIwQW7aQ3WNQOZ1z67D+NN+TjuAo7u/PtDxoGoBiurK
OdeSACINHnI3ZVj4LO3Y+4sVnIIFbNs5u6aw3hOKsxjVdTVbMS98NIs0Rg35ZBCWPTiUUKXWAdbW
+tv26gEs+4WrHimoeFEWtaaKB/5D/JvPqIpFub1uOlHFKQrntxjamxypRXOwAIQMU5YUHqlKgySj
RXOppLhE56RKIZUpT8TJEUcWZwrOLmDMRRZrYdoGX4HjBfz0z9q0Y1MnkP5DPqSxBdKlzbzY5jBQ
Lc/v2YFav/tqicoh3xgUVjp9H04HpTwhsH0zUbBCJJ7iA4vw0ovW2IJhQTarTnstPKySwY9VJfyl
Nvy1fNjsEafJ4cCXGfF8SWFD3quOLtuOiw9cYFGPS7FsonMUw1HtELaBSvLxQGHHmSw7pvMqwpoY
sv9RtP4gUNICPTib8tM3xGGqmTciwRGqmGcGVsX7v9d4Fh/Dy148HS/hLG3lZ1UIRdbATncGZ9tZ
a8Ap6T8u3pIB2mVaq7jYhwbhAYj1f4YWHp3pubAVuOFlbyqAo/EVXAIvtjLJGXPiEH732hJ6SiwS
VfbymGafcB39SXPXhBGMY6GrB4gHahT3l7dYYYIN3KkKwIbWwfBqfGBY/tf5ENI9/JuP2v/uX778
4lqvE05K2vc/Dl2iONHEgRlbkX/q/9IOqkWzwLefzZ3EjkUrpCD3/KMJdfcEjS0/QUj67+WLlIri
It7cRQEntoG2UocvjX5XYt/tKQ5p3C6+k5KmgnDHzaIgR4Nu3iStPnWOv39DXENCNzF7mHd89ZCT
e9c8JXlcmUFL3+EUBM06BIIWkkCSYv6AbhyZpngkVJ+rfzNgMJ+ejkn346Ba7vstAsZkcBTsDAwo
4ely3n10hTHzyzuxNaDDdUt2ZrT0YgXBvKcvFLjFRL3bYb2xfEVlN7sK3OkTB0h2UbqRBdEsnpMp
FGRnPzhq5YX+9JsjdO9qxWDhW52SwwG460qvry8iceNM1btgMZndbYw/oFWViwG9IeOYj2kPw5CP
G9WR7ZGTHNZfv5PniZ7OTcwBac/tBMN6kudeI5tEaNWjtvjW0nIu7pAVJ1HKXzWCHdDmqkNFKa5H
Q1PKEl3xdfD1j4TpGtKMnb5fdJ4z2uAyZ26PulcMgrPD0npyvvuqG7BbE8EZU2WGOcv/DoNX6ZZK
9adIfaNRFqS6oPGI3a2WXiILohoerOdmhT0ypkbDHC7vo0/hH4xT/2F8mO/rKJ0nmclUhhzvtonT
ALEOkg9B+03m12uhWw3JIQDwPnLho4AzK1jbj/+GtsxaL96k1CckX2o2bejEpCnErSYIOzWLXxxh
t9hfdJPjzvNxJITthy62XMjn/K1oX5D9dofvTXL7Vb+9occmmKiKNJY0jw3eNceSo89GoSEFa2lx
Cppkwiz4lsXgADJkBEJmoRHAYtjOdsYin5Sgzym4QGj4n6WeMxyIIKeJ9LWe0G4ChUK9Z1dKgKN5
bbcC1k3nfUbXGN1wL9o4OBgLZEBppTubeThPp35qO4GRNOVRkenHQJsLRulO2HuOlKwV38Y2teqZ
FV6P+NToH3ImQEFBotHLgIfEYcewJhMaVXL7eWRlyrGVQYqKuMoHOyHwyMp8qp/tpFTcSPi//ztD
K7GG3T3DBm5NzwPkciig5AmAtffvHUHZFNM2o1yZOJmtwkFFhxUVZypB3APsxolitqLO4HAp5mvT
bWZmB5rnrBpp+h6Mo7YyVa08l8f+QwCBOHFfMO2LT6X1j95dlH3o3UwYqOx1F6n5z9taNIyj7s9Y
qSdr5xOknbcylaBzl1DcNg17LbM3kSuaoi1I1KVpBRH68XB1kYDlNBCZX33VqtagBUPj5ZH6ucrQ
I4B09feHB8QdbbVsGZwmyndDARqgWp1s+i5w+9WMs0KFCxhSzpUDwKfEUDWJspa2cKYPQ/2aIN0p
TC/vqTbQ4oP4uDuBIpKLK6gNTslANEcdaJEFR6YfS82V/u1udZ/SRH6nQ99CuKUTQ122sysf9rKU
YQBELbxcGjQrYMQfR3hZV2PTeVOHjqwojUGqrDRZ5Q2XJIIVTHAiViiPvwv7X0csH9afa8Owvijq
OuggSFyhTW50nnF46zWbPI3CDs+kXUfsTSTH49yWSNjJtcwz/ZKsUQsR0fwFdnGocH1W5RRIz0f0
ZWX+1yj/CLmSOND2LnP9MTQC9t9puVfR65DMYRHIzvyJihuYq4C05rl0tWYkF+kJRIQHofYgubPm
cIRTazXz7cEJBV5mqtbKN4gKunUqbhvBXyRG13Sue4cmvYbFZzNle0cwgMr6TAoVbFb3u71uRaho
inThnjBJE8qsGZ0dokEgDfSoBn2Wmv103d6w4m9/1BPqqXtrVWAIWitL7PqsIQaGXzimRbBLZrXy
UJNw9/Wh6jr8YUz1M+ahpjOC11hlDAbpvDVP1rDX13ck61oLw0K53emSgsTRynrF43hlVGj1daJD
UkQW2LggnM69amRDlWDTGDkAOUd09rYAV7PqBKFUN6ZSJxFD0TVYPzxyyFQ1oYiFrPVz/4D1SbdU
iMSSD6XKSKqLjRYVlb2VbiW4Wl412QkovS84XkyOgjFl73LgOW1lYxsLzHBOyShTPP+iBEV+xbab
+68gL8uhHWTCUhA00pfcr711uI5LmhJWGXuFWj4b7IMBFaF96XZ+nx6SAJayvae0xqHd/+03LFX8
wvelAO8FilS40SIVXUzEg6MV4YEFMeU2cxlA/1GB0e/3kRiaONeT4D9xINPhTPTyJlynVT17dpGr
Uy6sl7FNaDYRDrDwMA+x/CqcXdTydyuWdUkX98TtmqHyRthjjz85kaYisffJJkhwK+GQndd4gPjU
hW6RhNQrJAVXdO25V/EAfQRLqeJeoNn5cbNB+MDKBHEbH63crbWeHaU9Ay9IQtfeMng5LsCqKuNU
GiioaI3BW9/sbK/3XZ57qLcWemgHydN/vUA3Q6b65CkAmUEbZY1ZwKL8moaoi3GIgOR4sFFKo+Gh
TlCZg5pySvQfuBJ2+KtLOxh8Pt7y8ZoAh/f4PQo5eRFhxKFeFrPx5IGQmvXLwA9BF3yUia3n72I5
/63vEhWhn3XirxgXPwSpH1oVhtd+BVAhMmV9I1bnui1P4iAGyjq7PEcz4KGdzW8o8UQp/fHVfsZA
U8tyfnCnqOIxcgRl9sVKPPC5Qj5mfbGcl2tMbxvKrXTmru1AWpNHam1XpB/mK9D9yoFTfyCNaVz4
r9hc+9UxeZS2s5jN9R+Gro0/lRhjxutA8n2OcmP8HaPYCdTrFw80cN+yr9E/nNNUA9TadFeq2cmM
C4H5kyUnzAEOqhagGy7R0E9Y3CeeUz62XkpfvVAiFx0AE3PcVvpW5+eYMulcJCesvPafzLmbGvZE
7h41fwuD4e53iyaOcz3Vdy9TA4SwgD6Xxhf3y3v0v3ocK9n4uRA/uQwLTB1ptEL3YlWvVbqF/YAO
i+AeeFb7ugJznWozxKgrrEvbHCorNzErl61cSKjHT8Q6UTF+6zpxzczHUJo6BL5DB4vlSgGSzd0c
DrUKrmvbR4ZD3lwlYFRLu8qeqsFvpre3vAbV38JBm+BTUKJ+Yjk61tEHttpCw2OTMqiDsjKXOtc9
mZdL034O38JmbeJb8zWUKn5HRitzVB5o5wl4W2mZ6XimEF49uW8TXSws9Vlg2jw8vhhB5vxiSq+t
er4pWryaEaY1j6M629y8Pz05qwnL/Zl2GZ7tAhG4FIG6dj7f95v49xjtXiWzbf9Keu5e3GC3UxTi
uamCAzH07i115KtUMbyIEzMU0XTagXtAUooCzbvOolNMyFxkYdtms9PVVGfuQnBxnwvftP1E6Ap/
q4tEmtj7MDB7QyzgwPTPTwpx/dz0tynsx7171O/yMxhZysLNfRKjZ+M2z9j9cQa7ZIcJKD0Kzvep
8PVd96Hg4GNuSGXbi+W6rUxUD4n4I5+D2peZk24rizJ0CHWeIfRI+R1RtvsQxNgiKbD2oa5xNWU3
6GBWOhUSm/UryQq7NKT/v/pud2tUEC1hLDFh6K12+NL9QrX5aDHbYkUQwaGNEniD8FziWOVyXJ1T
6rYRDSOfXwwEhiKsq6qT9oChNvfKtryYyoOeWDsz/pvcFDKTPSPd9o6QWRlXQ95cxdx95i0X4DRM
8Nn9aDLG6WnZfjObplkKMfITiKwVy/XRGSum01DL0sRk2AbgEY+g82b/2LBojfus3T8QcnSwFKWk
7oMDvHusmbdVeqhwOM8R43DeSJnesEV7vzaupGRVw5/sbEZKnAngKBTf3GOFiA5MEaz2fjv9iBoE
/o9z1ryM2J7bwqpebShyO8OdFmmNx2mLBoFeKAXszQgWlk111GjD0ceYGDr4Oc/wvtnt/zZjYU/L
uP7ZOK9KVpW4BBinnAgusVfnyCVR4Ttb+gWsCixeEVAacwt+nfRrz9gsbuGDIByCaZmc+ZVobvWh
gbt6r2LynZzIzXUbAkbVZYqPno8uuxJNeClCRJkw663TiUUtIj4YUDp8UMbtib2stCVD+DZSGFg6
NnpZ8xsxuXFJCUt0z5B7AAQ5l7G8lkzIziVkvnP+T/5C/llyAlQH1c/0q/2DNBM6CKKGVjrdIzG7
N4A/wlVqWVqpBA0Oycyp6yrKbM4itwu4q2WRMPKyNx2iEAoqztLhFLYyf6ukv2ry+eUi4lkfpKv3
4ylzuOaeZK9E7j4JR4g74odqwgWlAeHE4taZkMwqD0ItRP6fZbfC3uqAvvlwGS4aGzsNHiW3d4Ft
qY9Z3IKEdGsncAOgwJyF+BnFYL/KWq8iupCtzHkTtNjz0H1q+jq4NRWNalGRI6l5IsAG+BJdj/D/
l/DzGtka4G6NWovmBY4Zb7wQtZsJ6yV0aG+qvECCTXWA/i//DKeS4fIGMlmysQmtgXozbFpYsWb2
5AtR4r8I8zGrkyr6kM+gfUcjfic9ljpmnOlyiA+nVMamnIou3vw318e21oYzL2KBRPZZE41mlV6U
QTnKrbr+sqHou0vc5PLM7uebCFBKaqKMuYV6vpSrnbXkKqPXxxvVjgU5yPz80Z4lNSeKJi14lpVl
cbWV3GzRcPCgZDSQinbxWv5UD/7aVFSgAA34ZnbkigVsuryRUqWqoiTfkkS64ihCIY8zRsxnk9Bx
UTdsuwtEkfsKt+CgIzJ/HKk0PIwCdA7PGp50jyvOXzluy/gd7PA1bn7/H0cVtYZopbeEFtopRCs9
xKm2K0wV4cWmlx917cFr+BSjWtSf+cjtUhou4m45yDfGsgxfOz1ouCd+mCyO+QWI2MpF9msXRSXq
UI01tqk9XynX/u835XP8JzfosUVbcC9pdi8Kgn6+jnjNph9shvS8a29YeW6R/UK/fUoK8IVxe1ue
HZpbwLghd8KmlKhD/6sfx6hK6uN9DIDdcGtXlTFmBYXMdFgk9AMZzFoRNCUEIxwgTREPf3J+gWV4
JWj6Ti8LJ9XnsZb7fvMMiJU6itssgME+L0xcs9hhFGykJWJXKxZ2iCjIYitIKETE/xkpjs/kCr5Y
U/0+HnXwwieXVyIiCB5eN2rOCeNgwmhsIdrhv6uCeWSTrblFY9zdDAhU6Hh718hmlKgf34skXiwC
tbU6EM1Lp7mLTEiRTxMD5xVsVgKaVl8quDqQgpd4mMVLd70wVtawbKk/tW5crivS7z2MhQTDheLJ
w5ScMHmWOIJqHQKucM6FloJh1GdbJr9uo8tYFJ7ycj+76MT4H8hF/jppx2iNjPZnkavLkejvebnN
6nxxZC92hQ28behMrguh0KhJjfMZhhgbGF0oNxu9cJjJMchua3bR7TEPxv4PwQmldY77YAkd0Ljk
ZS84P3E2pLnpfSQurEYV8xAQY74t1tzwyywZjR9L7p28hsEpnmjeXocOr7uaf4Jn7Uc/jeyeCLxW
rzgH4bVbQrbuo1j7ZGSQTKvefgoQody9cef1duraIRTp2MM87LW71QkUdrrk8dISMS0IVTMGDkt9
OUXyRJSTBW2Htsi/NlO28mIXkxKI06LA7RBKEqYj9QBaqQdI4dY7ChIpjpKtfzZF7arEmIGHbEYd
nJ0hn6erh+SYDEl4xHjvX82wPvMpII7XT32rBv2qIOO0osZG9b6K7qbuBnRflgJQoBf+57xz+FuV
Tu53+NYg6CNGPXqfDtB/GlNkvYBudOWlGnHHvlt5s3EgQ93wiHKQU3leLD+2G/xOsaQBpDC5PAqH
sk+eKH3enpMgkEZftdR3PekgiwvOknCqmEnhnkK/J5HH2QRG6hZd285eE4xpzedLJNK4MXg1BGJ3
o0VvgnC8iZfQYxig01sJfrl8UctDLHEtg4XGG48SgjGkz6IhRGXqXyOBp9t+tANm/9Lq8Ug+0y1r
VnetG1hIS2zI4MgYjZIoqX7TEsF90+1OsbeldMwGgenKIxsV/ljfDYF4PPiOKPrQ7Ncfd5rzrcB5
wPsKDTR5bXiiAl41i+ATw2icByfAMGF5OuMtZPuDDuXn58uDNIUNjktQqBJUX21VBurzsk10a4yJ
xWCQ4VWJWDnJ8QciCntPrkweiE0jCW03NLx0FbHZotl4pLhSds7s11rKHWVkvzBI7Vc8jXpI+Ieq
brlXlwsb13vomE1rgPr7X2e7jVsCJcvq+GNWkUwmjuOo1Uuo0M/DuvHbaGqqBnSy+XbCziLa8HWG
uTH9fmU+kwRNw5X+Zrzy3rUjqwDsCHmN5HFUY4jNv7+a87YXbPMCSR16Ig754Y7tujshpva14zMb
riOCm3xoYZVmehoZd01q5A4mqpdvvmpg5JyWLneOzJ0HT+/xKJ3GJ8bnOCtvNZ8WKKDz8P2TJQUm
4y5psyeev+Yn14al3bBBEoUpPSVHUKGqiF5bJChmAiE6nhumx2021gxrAKN5xcdPZxbBkYNkUtqF
DgGxEsjxCI5hHDlDcr0oiZMusTgsDTCMLvLT200YJbbQRmNYjeojE6lXjT6pEoSbcFyBlfXy/mLG
n57GLa4NXPTxtDgMN+z+0QX7aumDlPW+DHFPvygc+j3UYb0OuZCkZLchTy2O+cihpcRy3F86p7/M
dxSzEiagu8fpe9dy0THo9tU2Z0S1Bh6OQGt4nEr5KR/UsJrU0Y7bmbopOvuMMpTrGgxHkE6adwMV
7fAra/2oHB7FC8mZhLJQM7itciT+BauWuU4lFF9nP+xcXAbAIZ2q3WNAt4mdPqDQ9Iudq3kOmFW1
oQg0EuZC7frF0PtmczgBnXzKHMje3w1xQGdb+Wd7idDU6+Ho6n5CwF8IHLhqZdjyLrSpjp8UWgkx
/2sb/DcWZZfLhNnHLcZCGMrbO5YbrIGwrcoGTyAYXR8lhKol2Cix8EamWfrX67MVqNVqopm/z7Rd
k/ndQ8krfPSfnlWOplR+EceWr7kwtwB9EepvayVCVLV/UQ03eCxURRtukwzr9TUrT2F0Nk34MpH9
nHxSXQzHM4PFz0S+h9aO3Eh9XW2ojF00OvLuRnDCZbJU7vuU3leGPf9E1Ii+8WQYAXSR0sOJYop4
DmA7JYkk6ZsEwPDgUsYvGvTjO5C00a9ga8U9SWdwXeTw9JCQdQD9ruInPKr/a3MXLmQlvgyg3B0Q
VXU96JuySjkHor51pLQonC/TUo2nrBIIYpNLNLV7EPZJEKktqcJSnYOKJq/INyiTHxCSPWdAVl+l
r6WXsQ2L2ZmbF4/7WpSPiWur19rMrqSnpMAaWe5darb8OdgfHGHolfydVtEWoxKvIp9dZlL5/tDD
ni22Z29iluzyo5gEY6IAo01O7QrjtA+X3Yl64YaNBCTEiMd3zExjC3Hgn3C/oUT81ydU8WYhk10x
K/CuD7ssZhm2dDTwyboxX0/lIKkFS5pJgKNcio78xPPm7nqpXjGKQZTBZhFLoWPWukuZ3Hy6zl28
RTtlgZkW7giJJyNJR4zjTaVN/78JtjmJjAwtc4hWYKsoJWXO1SMyOdxBJwUJVjmWMIPgoEjkYJuL
HKpQFsu1MHenPVvryYLeohHy2L2sJtsZXm4zX8C9q6hTwF0LwigsDUvF5qy4Gcz6DH7xX2K2wXI+
FGJOlRP2OyYs6hXV261VqV/RhkbgYSFMxBdDJOwNosycft84oslzOvmcF9UN5J5Ri505udwYqr4H
5zANUcDiyAeq5h5Z3hmTS6YCPDYx3AO1wt9wHU5f3nNQQIvJepTQC6Nxfn/SOQSDM3/vrbOfirFh
37mAavuZwl+d2uWXK3nykIB1uJbW9ye3wW/GjLyI9+paQHbmoS7by5znaKpxnGVPr9iXVFgJMzDg
7IlP1tSXU8XSMZZYlXa5dX6eet+PIWgPJ2uAscfRL1MudxoF9SNL8cEx1qWLkaeZutHr8TqPJy23
Pl1uVZrBnz3B8wft8dradKozgD+KUnwUQvxW/NKhJilY9yMByc20kjSbe1UEtOnCCZkG3+mOqZIp
tIm7hVSVkLWDp3T2MIdHzqt18mJNpiDI/CtjAWCJgnV068OuG/25AgTXNdN77/qxNG9LXYGDHHDw
fDvR0GKEUftIAgcc/gqBeR4/quTh0SDuYFh7SUGp5AkMGmVSaR9M84DAnW3tGudPO55EgoQKyWew
wplg3EuprPtZ4vNCY0H9uaSfEC0wibjoiSbk6UmH73EmTTv3RD+8LZsdn/BR6SoXwYg1rfSgoFGN
L+J9Mn/LywsZvGIpNxVpCSoJpkc3OG3VNz08bxUTVmtjtT6WzbRkpM23h5mDPWW7MJAJmJqSoFsn
alBR36rkvQPNA3TdnZOnobMITkoMNOLB0SSs+w1lHDdit/SCdspwMa8e0LNlNcjW9mzo7owTkSnl
Msf0BISimozpHxLojeM3QWH0LN+C4fwoC9rmC6+GdXCbTIaiDP7M8pw+UZIAbTkv77GJQaiikphL
10Kj7yur5vll6Co3huBo8w0TrYdl/9t6NmCg4GsMXYSVb7eLY72qrg1JcvK4zwTjzco1HmFuEkSU
mkCZMyT2094OCcubXWilM1n3QYNI+Kg0R+NOoZSrkQA5u9y0OH6xcLFb6kxUkn1scVjpkywjhv+U
jXlQ7R9/2OSYwJISNBFKIsRpLGF7hRjRNw6+XLX/ChiLwGPy5ETKUeFnKpnyeLIN2HX2HOfdGjtv
BYh0wPrhbwIv560dCHkNjbuVWoeC9U49BuSD3ThGGyaG9l8IsKSYGOhYcqTYqwsz+I20HO00h4Ia
veOTY+YPshOks/PyIcj6AuSWkos/LAuF0MV+K8YBSJTKIT5qNYaIjxopGyZZY3HmMArRlTpEu5aa
pGoHSlweyK5bzW47TDH3TlB3ubrykvfd/UwXTP5br4Ji/4ZCkVVOQVAT8fn9cGkN/Ixrfyei8bYR
E+DpGaqb1WhQpaxS+LNQZQV9l6nKuiVIZYOEn1KdVybWoclssgH53mTkSs9hCYlrXf6RnDkG5tVg
gtH6h7hK6Rjxr8a0nH1Lx8S1aHPo79T5Sv9RvShPdIjsS4tHyF61uGm9H1JyPbD15jjIHRAUAoOm
O0+oXodrGPj8lijLZjyHHn/zaYDDUd8zg5RA7KbOnlDDhGv+wZEW10yXicgaaMjubqtK3drpXwmF
W/4N+B4nJCTCHE3YY88cSc9iVrYhJ+KGm4gxyR/bA3Zff8iV5YbFfG85RB5aUZlBqNkYWm1k9ChK
ndAno1V27YNWDYVWDqxuX7JxL3NccPf0WOzUsR0wx4McYFfmfvhr0Ha9RBoYRJax1VeSOBPdjHwu
77GjUndDzn/QyotSsUvxmFnxg3v9301YhaHSkxcP5blZLNVUczaV2KdWh07qa/4PLOJU36WNXpN5
U81zqCFp3EvcnxeChIninaOvKS+hMw2COhNs9FIe6t7vkO4pFtSzIV0TJhTExzzK1uBfyrPOvgFc
jRWgrwuLrZM14g6CXJ5VhvUlMJXoA0x4Yc8V+SOahn+vDU0i3b30UfRZLVqGr6aAIXBbxpnA3TZG
84AKmPdCPuZrO54ypy8JIuEh9IUe0/+H9SYDyRCGAWMsJoSytfsIi4J9NXMQ/aFGuRFzZLxKIJLv
fD8cauI1vxL2XqWDDUWYi7p400blJUPmfGZstqGXXgwLzCh351gYgwCcBtxTSZahuMHF8zeoy9EI
ilktxwBIEB6bF6KIcluXstsEU2UN7EkgmcgTN/unGzwEAmrpWWu5NsARCRK+ENOkKp60QKQQb+Nd
pLDYp5rqw9QfOnbs3GnAXyaiqVfSuWinPimhL8qQp42OeUJbPDBFVSaWEya4kV7aJ7Y9NfgZDWks
tmJp6/k3weGyjUFafLZA8Hl8JAiA4fEKyEuIGYdnw9TlP10/0hoNCKrWbypMjudZTFVRaCy4TAlM
6lDTNpCjEFQfEHeEvDIPQc3AQkw64u2GKOf3NzCTAtCxbpOWu3JHFYReT1DZAIW45SlcYyO0nyzB
OvcLWh1UlZys5QXmK9rJfVhuk1IK3TMfedZnSSQ/kG7ZEdTgtBmdWZbB49aQ3j94PTekhRp6uBcn
l4uokFsZPJf+lzygjqQKyHIs4ky+97qxxuZ+os/iqtW2Fo4H4dHYWC4WUSwfxMZ3g7Gz9yykse4D
mzbLHe6jOlqBML0WTDn5Okc0EEARpmXMOyY7uXBaBMvY+peR25fgXmFcp1jDk9pZA1Iwc/ScYVbj
hJYGOepg+g8Snum7BvJD7N0y+KQZ/GfMquu4iUVhqMdAUstx7kFzokhY2FpUoI0xCKNUo+MYNP0P
DcMEHorOOHMc/UoftVFi4kUE7vCidArYuRAbmYpiGJ/CrJYTWKCoR92Na3l+KTw450JMlWQqxqoR
D/uXsgWIxnKecQYRzwDDht1PCy8FG65M/ayG9rrl/Q13zCagLRnBQvCRZWUk+39tijCi7wp9Izo8
aR9nCcw7QIxjNeiMoTHBy9DlgYc68iC1aYvUEScCtG8R+6aLA4q83WJODFnV9wFBoxOOhW68YqPK
NjmavrkJ+XZ3QobJrZ+BcIY4CGqaVSONP7dQnlA9397WQOJ16vUgmiXhLbYHVD4dX98Db5t9/opt
ctWv2ePiI38m4nZ6D6aoho0RSae78sZMjK/yFq2lCJ8LGkA3sgns9tPdCT8y5OrC11cVl6LycVeJ
1+pgRMD/xjQEMiTW6aR1fH1w8Dk4HmReOax6RJ6rinDq7lH4j++FoNEg9dj4fIlV6S750GZmEPSB
iiMmp5jJeJHpCJUOwTcxiRJFFaxTefaFEIe5IV37P2CGoPyZ/Ex9m6iSSeLEXik5DsVx1CcG4aMI
lXXmqfXI3x3PkOc9l1RgIRgw73A2Cx3lAJnHXFu5OdMPipnzwOvk5GFDCRrrbLOqOHhH5l2Z5Yx9
Yho5MSMWbECHqon5AGja2tbqDsHJCB2o0wlCNvGRvqHKssgnWfMKokeMsziZAm5kABirMGeJESVI
jPubOv+r/+Te8jKTrZb8AX27VD6Q8X1G+usKm8Ow9B/+YIFI6VYWbl8WICGgdI77O5mJ0V3Q/jYL
+RHoRD06I1vYoyF+g8wtR/u4xXak8vcY9faWJwpOi9Q/NYv0FXuHTJ+aKiM+EgqhQJCZstG49ntu
O/RdEKPBp4kd/NTl+Rfx8eTl4AoMJoqgB6Gw8oA5+rQoHQCoWSbLpYtnxO6LbzNse8qQ3/q18SqI
kHlPausgSToOezsTyWgNwyR/+xPVzeAe50jkKHQSNGRaRl2AlShedo6uletgKRDaZjT9esw8mtat
GwqcE60ZqjLUmNw/tWzYOmjd7/Nb5NQhLPPCdAxAjQ8a7qGybI153Bcsp20vEyKE3CWFQ0zqTG0O
18ocoqUKIoYggqz2KMNGo4sW7KjGfnolvNiVK/CxfgebkUHe4tqe7nqRU6bhe9rpLc37Q5TGtxZb
wHnQdwsGiOx2laxE8WAwEkXG4Qf7MDyE9pLYjd63jjXFQG0bTjp9MQhrQkl/gP3GA2oPGknKUlFo
SNi0x341+r/GzXdoNtWsQgR1Zz/sTFpjYE8JaLOodplAmPYO839ROaOcEMNyIdTg/FTlW5SWX5sm
xogQUizOU5uVm63wAJYZfA/4LtHwJ+6SsG3s+uQBFxbufE7/MbOYldoK5RAmNrPWZM5ACEVFv2Nn
ecsqvAKQIBHCiQ0UY9BqsZMUYQz9+chz6oD2up0Rd+a4kBkpSqyIDJDiKgsbIUr1dlFirVMtw20t
8OFrwm6cTXdQ4ReMiW87ByIJ/nWT7qEf9PUcyySHdluj0JbEs75O6TX9XOUUQUQuJNh/PXXh/CZP
l2Ev1IymaOf6cJhXmNqiPoeIJvt+y4pkSiemgGPTY5nL1+ORTrJCwQIu1qVEQqYt0Hv0cSaaHzLY
Q8WaPMrdtetFHud3IyKflLsCsa7zDSJY6/PNL6/AeyiuwQOEvNDqJMAsa6ijBM5rXgujt/b0Xub0
noxKriXFw9NDuTely6RQrygbWMq0nOTJDHQPQhf4E6h5xCMqAMXfC0mQpskSpRtVanBvlZBxBq78
9VhYCR43ox5rQinrSdBEkyBW43ks8HLTcIokQUr1E26y1vos++56vVy9dRUDbXcns+MM7uXlgc3p
z6smSLIUpF/MhYWTKjcp7DarhQut/KSEBUhXpV9PrAQWrLbRkc73iLaFWPb9EDdWr7QGxisjQ9y8
nh24JMwIwFe+FgpniEfRzDIPMKBKc1I1Ldkil6FFRQA+99AyOzJp0pgAw2iqtBliAZozeqfjK5u7
1tY0iyjqVgaRcfBu7bAZJAQKj6LI8ZTUxKo154if5AtS2MuWuTigHV1axw7RuY8fsvSZ4zWFiYnN
GH3W8g3Xd/6G9BKxA8nMWZ/ui2+92TrhUZ/d0voOXWa/IxvyKwBIpO81vfesZ98hMo4UpEstTHEB
rDpY/I7kC/5Y1/J0ALE2N7/w5oEQS81P3Nc1D9JCJJlV+vJb0soACg3QqZqD6wxKeidkSOarXuJ4
LlA0OUSOxhSpzzbeuG45x8JsUTNuoaIZcySB7ohIbd+p2XWZdO4MVPtugacLoD+wTj2mCI0Lal/a
3fX5c6ixSRNwHmXfvm3swOYfzSLcwC2SeD3ZBS6qe7DCigrtQqc7OZoD/ZrkOMYPftV6zetCqmlY
3e8xP/AV9z58Ul0cXcHME+dtUE8nUehjSYH5iRPGSQc+iPUkINIH/AnBIzVbLKeXuszX8aHIQph4
m3f9uqhYmghBqEVzHNkC8OzeDl8+0yLFOPd9wI3g/yOwuk6w4B0PUnpGEa3k+F1X4cjsWpHaJZhj
wfBI61TTddKMZvdt1jb8eS9qzR5DIjr+9DCz2UAndnXzsc07TwvanP8ZfIjKK0L8ZDsAVmq0VCF1
7zegZYO8wWBFBsrPPfCYODUzdbTSkmiTGKEUOKLtbGfOV4HGpCPcGWx6WI5fMm7ijNbJIW2GfPxL
/4kdsIzYmABFIRGYxmSiWq4GVc75s7egLnBMUokLN5r2hPaXkUTQ6y7ShEOcUpblVPIoYj2+4CC/
/HjH/lw0nbGk8ofBN0RSMSwmyzeY7qCwV4s/igphZwfpw1S2JYFbKN+5nSYcLKA5C7jhi5G8kYzx
UqIM5WLjldRg/uq44iQmbe/JfAwrtlVpc2wqJUMDTR+rrPVv3dORM/caloUcsSal68Z4JrE09Wtc
R1Huq8VOMLNMgK6PbinongzvVz7PwqPsh9HL6qvEJMvsjoTsD0d8z6eN0X349Vp44qG9OdiP/5VC
CkrSN3G5329kVLAMPzfHJfnYhJ8htM51DcvQmkndSi+IPnvy4MNWgRmNR2z5rorIUhbmEzKUpRfU
HzDkmN209W+9XKzm2/JoBJ3eaUWncVoaoYTJ+jbVRK+RYisOgYN8Bc40YWLRyEo4JIqy2VAIj9po
fWWAcco9BFJN3YRrwxEKZ+e8nhoDVud0oc8yj+gm/KNpAsk5J0IGt4v1fVJVpDJ9nOGmZPLSMzsZ
UYxKi5xQejiiFny8nWwJpwF30RAzuHEiTANrAxQDntpOuKH6HvE7DHYdw5a8eiNFl4Mrurf4CqOa
lAGbvWtxJmYO9sJFUQ5dzSmsrIIOnn967sgZzZ51URDEhPoOgQWr8fnjywQiS+de87u1bsxBxA3q
hAvpyHtWt2vfytYQWCAj9RYBTbnCKHMfYDopmrRiAuKl3/3HytUzv0RjcfPTSsi7UcCSHwVCT0Y/
lU2AioFcv4y7BmWd6Nlzzwkl+w2b8C4RYF8YB4I7kJgwisNnmx5ui1glqGMS24NXCL/H5V0xh1wX
YlkykalThMSD9qbhu0p0nZrvvlwiTC33V2+pmSsoKLMWJ03BAHhDjd2jIFa2APegNAZbWium+On/
4o+ECFMIY5seE8tnWb91HXB87AnQ+jeQ/j+H1oleVppDdavNr9K8o5RTMrr72azgYW/JB63m2H/A
VjD+Lygm7dXmL/Ad6X5dRCtJByqSEaf2zxJpz3poxnKYEQ70QyVSfPJ3VdRPsng4pWM9pkGu8BIa
UnhH5l3hnbm4rQ4Q/sybQt7ovcZO0eSUH/ZsD2BB7hhS+/StzZh1BVUhJlBayeMJQnCorT5c91Xc
GVC3mqUOZkKWQArpHV+zeCd1CLYqJRvdHWR78Si3510wdYGoCk+6OQYSHlo0+XEZdJMNJBBPPzoo
H+TbY1JxOcmF5kNP4RvqazeCIE27tOhF8wAVZbvd+qFfBaEuv6pMJ0BdbEeLsopR8RiB5pEr9VTX
+bNndlT0lste9Iwfk14a9hstGgj4W5c0GtSXfPQKEdPjTip+sDHjilyNgPnNQA7ddNrBuKJ01Uz+
IYrddoqudH/eoxTrI80djGgP077smvUxrgPcXw6bHh2xr/D6hR6uJW6FqN4GA/eciL24YwxLVyYK
psnpzXESIXMzJq6Ef5s7x+YWDoojn1k0okUOd5ZvFEILBMvqmqAHQmIiM0ybL18MpwGyMY2PULOq
yTekHZ1PUqvYXrZzu3qiuWIkhHphxMmwPDAmAEJN3SgAQNWM8iYaOwuJEbzCW9Vrd912YblvneVk
nnqNK2kxeGFeizrIm8iK3HIHiOwjYWqmK1PAGhqlOtOssqPfdHoAU9KHD+piy2hg6YokbguvkNZ3
RO9aJJVtdmh8yEg2kNRaEARrWIKx2zrbBRgSxF7vLXB5mcwxQOLNQVCPm0po1/zBt0AlCjv1eu2A
x/kMoutP0f5Nh22o3uEccdROwCR3zZVOSyNSqrSpt3vDsCbr5s9N8UqlrnP5hFVw9YYcVCnpZ19W
mYnjtEdxNqZIy3OP0+al39YLS2zinAhOA34k2cgUho9YBLfRc9G8LAciigDd6S7c3d6GJw5WIcyL
pcnPlvw3A91ffe5HGmZwWEkeKtRYTSxFh49nBj8C74HxrFWtEADFR33Dl9ItV8W6tOauhjjl2oD+
2Bkkt58rpSHj3FPkjeqvup1Oy5erPYVQoN80E35kXWz4LsitRu6o5hif0Y6qeH0jqQPNNfajG8e9
7ORfcTS07rSI+pq8dMVyZl5bPpadMs+4hhbTOoPRH99+kO64ya21u2bopleMxYk7RQXqXeNWuvUd
BWRBNoKp9pKNe5hydFRHC8LC0u8mReJKK/GYmba781/I2fLpeXV+qQD/zrZVEaKi+2BlC5qGJat/
DYaYywzvGZCpspiPu/o9AhW4Rbn7aPsUeMtwtRucFgKErjV67P6BZmKYNvVsMzzeaJZF8WQcOzEo
OBgKt46wAuO+crmyvi9AhuyHZiVd5WitapNvaL9/GvHVwj9I5zwdwNU+ZE92noUUKQmL9H8uLTzW
poIhiGKD2tcN+QUVK5ViLvbbIw44N9K9wk80L5O91k7phztuADKujIork6hSLaQXPXMsfBBxxmFQ
WqxpGaKro0a5MwYJ+q5sDtLmnHXE5t4rYsaB/L0kKWBS/79qmAR3omtt4l04boMtX+UfuvmSk8p5
uksuMy8Rz1ta1B5cD/Vh6JSPoYNnhpAx0QuiRn4dJJ+ylM5WYrXOQpA6KpiNrxMmp4+pT8RcKXMV
kznLUAkp6x1pbBOdQOV10Xkpu5DZUXJQRawXZO59yqgonumx96T2t1QfNeO8+HGs9ohUEjk8lF0j
Fb0VkW79KzY4/y5Tmg3/KLhCrlCK1TEYP8CclknuE9E7laKIJ/Iug/sOEJA/SDmnQ13nfeh/hXrp
jR0NFHbTJqRBbSLR1cyzoVvY28CiaUsBFDIRp9A3AXyQCZGuh0iaRoonenmG/V8snqaCSWKA+2Mg
zzrPRPFLkzIgIUigczr9BQCbdx4jDofYwqGpGj916atl8OKymWZYLhg2YfoPdAFqJ9ix3GHuVSM9
bBZgjWPRanTLoLL9zMPy82XYXimzB10mjKUTmMjGJbanVh+Zsg1J6guJpAvXhdUmAnVDvZpDPgja
eaAIHgt5l+vGSXUKfJtZt+nDzGZCqw7+5PTV6Qq82wufUU17mQq1nNbZVcqCvJryEHRH/UxJAjY4
OIIIYzAG3MAZXB7W7lYkUdW4ycW3axYRyLk/D1HY+MYm6WXTDUlOrXLkTX4PgOM0WAb6VhszmMgs
A7TLr/kvfrzQrzhyARaLwYjx0/5TpLcj8emE6U9NicgfNqyeCXBhbBb63kKsOV00uke5sj0NGxY8
kfze+t7uJfXcdO7B3KJtt3wlDoDfRgAvzlO+Hk0wTiYbzTyeRWDzZRs3LGj6d5nuJPiAzre7xaKu
r9AZsEUzkQ0wG4V6o70un9uO8RB13ck/4kJQIN3zIq5e1PNmgmY9JXPF0jQzb+OOQsmJXzYbvlmg
IkSERUFVzTrvo2U3tePxU9ebHr8vCIF3nySk0yVHlAFMXVMjkhtRGwhzuWjpcYwzATU9UtsXAR6b
bZJn1q3yNE6FsjIpYTCYsiqa0RLCOeJZPuuB+RB/SaDJVaJfPGQxJbsEe9eKz8mcdDIWi7ZvDO8j
p6MV/GPay9yWwdoebCy34LeuLz5R6cXhZz7pHA/hBdUpG9KXa6Bgv1kg8FvMVQ/ux9qz2P7/MyR7
GNAPE+/4nKPZbHUcSNkFokpUGbDMpApVg5sUCgEr9DfGh4CM3IP6iUxxFPI/ayBFH5wbsJIsB0Pr
wRf1Ntz0x7auKoRrzBQyAx8c10p5XOjNoY38iv/+LQ0sp2wqVB6zr2/Zif9i0HXLCXmx1RF2LlX0
S3ZB8/m0ZJcMppYiwBluTzeBFGHII5YPVMOZanQP5KK/5J8BHv1WTgd0DVwo9tKW0BaO47oKuE8Z
lU4hJXBEbAbQQir/Ev8ajPKkojkMoZQ6X1q3wBrJaj6xWid4Ju6wfHBitp7voPRUtw8CEMmwKY35
2DAycwwQEW4lNlMvvRqrZJ5a/Uw4Rys9V8cLFacxkg0DPxJ5DuQdg9zd0TbqJVZO+VSZnJutlLuf
hLFiql2eWkbS1/e8y3+p4uL7zm4AFbVlGf17QIV+RH2yuAUHjwJm2DSWopGj04nkLIBD3Nku0br2
Z3BIt/5UaBjEDo4F9SAYxVY/S6PwoLEjQpYLDhj1yLe+WuUSC8mymSE/ADRB1PC9EdMT+csHqbfz
GN+YnANbMvqet0YRmT3ePh7x5OsrXksjR59oPgY8r/JDbiwscNOwWcEzp+pBvacRK0mP46Z/f7O0
oxHsWf88G3xp5C9dAB/ZBEmN7B+OmcSp1S31LzYotFKNuDd3uCaVTIinyKIeSMBXxyfS8plz/P/O
OCb3xoYe9oyPml75lxliJd6qDeh5LpQ56CPGnuW+MUqKgqmxr//f6OafXOrXon9T58hecYUYdfKD
t2C9ESWqxX1CbfeJHP4pL1NeqM7PLmD1xG48Oh1QltUIwZMGh84giT3ld9lG0nhjgEVrCOeCZwMm
fkpRmYs6jpawOfJUIFj85Yj32S4v1sC3VfxWTFnGDn98hgxZxCcnSO4GKUgxEMw/kP72OT7nJ9Wx
G6i9WF2RYSFileA4cmm9ANTJf6iIU9kx9jwi94JSbZ4fskVPv2LMmWC1c//nQswXONTYoHGkIc8P
6QMPC/NHZhe9uC3FoOH/83FdtaFECLxlMucw44MFyFbFgow+/0MiW7KzUmDEHNXk3HgZy2+tSzSw
pMIUNZNw05c0teRqtNRpgo6mwPBFJRf6btWsz+QgDzY84oQbNHZ6ektOqoTmdGQyEYamdZE5O3d1
8Ve0ELGPZBkqkDbWcjTXDf23qdkB++pBy751IZuz8tFETn+cj5p/6QSZFbELTIPRtt2SCayPiQnA
JzfGS19brt1FIqrXFc6lPUf4vrteOfdZ/qowGWJZdg43cd+oWw4q0bZ0TrKtR/yxooE7d+ryIRr6
qGbw8MPSt9cjz6P9ljBEwKngUDlmZRBCC5pvNWstVzw84eqQuB5g1VqRJy221xaWZkOiWR4+kpLl
yoqT69Ph7FWDBta4xuH/lxY3c56HGrsIVKKtCdIYqDZyOUEOMbeECnKCloH8iEIuck5GjD0Jlvwi
N2Nm3be9din3dJHfWIXuVbkd+YIQN+Or1rarUkeUorPLGrbSggc03DjcEWWNWOLX69oreKqfjl6L
swItItXk5me3SXqfdifN57+GC0fb/9HkiqubYqFnq2JdGSr2qZAqHP4GJKMY3o9k0+yQ8s2hn81I
U/PHn2clSZIn7qmqo2bYp4CJOAuZTa4ydAkxhlQs53Y8RkkDEP079lIheAh3qMNgTCK/GtPQPjlL
7sNo+OY8x+dHzmD8iUuHVfOR/dF1MWg/3xBVfhRbqku1fyQZPjLMDooaB40kiVc8jMKzr2xvhG6S
KKYLJr7egUsqaGNAaPshc7ej/VpPYY3A4EYhk5wJEvzd8LnGjpC6K90+xNLq486Ap4PBynMbpxKq
aITFdn/IXoOU4fXacz42nEljjk/+LtnyvpRk6lbqWZGkb9v9G96ROi085/25VjDcwzQtpILQp70b
80a12vA0M1YMSuGYrZMG34vRqDB6nC7A0bJlp1Lu6M08Vak17CZUHQA1m+wM3NNLHBj46mO0ZPNV
fJnMbllgcmlUYQzbRr126n7xujmcvJGhXAnowVUyGrsoi8cExdrDikV1OPqW+PDIEeW2Uud86qDy
9hSt0Wyd4wYF/6fI2S2RCXx7UQHNhVCdKBVnwrrfBOm07sDwFY+9d972zyAUn5PoWL/AHbTcBWfa
Yab+h5IuUeZNzxRVPdNNbgK9q+USZNwGTErGuzTK7Oc2DJ5l3lZeZKH4T/YnlhhAf/0BzwvRGcMS
hm0okAWV1rsNuB2CjZFIeQpW8DjRokxb9fKURgmadHYnbO2tj3obIqXJ4MUqdOHbXT1zgv/aw5HG
IDfq2N7u75o3yoTSOM8BV5fKh2oogVXzPKnYHKdbnJe+52aJ8oA7m9Ps+NV647E1myMqF+ZF9S1E
rVhqK+jOQxNj+me2D79YhKzzbUeoAu+9DA2/yFea6D50aoOmgTK5D47LbCFDebJxvUoMZTaBdx6u
AhjcM13lpJMU+6q/DuBMbL1npFXwTKCuYvsOUZs/tZ48pWxLbizSEba82ceHzu1bh0lsXOXUD4oT
rY5BowkmPA0haNGBLrjePS71Rf1uKbt08V0Q5Sq50oU1fU7fxJdbDWUc7ztFti5qL2PkMDlavgMj
sZOuO7t20Vw+Plq/oohHz9QUQlXluo+OITsGrrTgGFoK4xj6vFfa7IqeQ98L2CauxXlz6ey+mQ5R
gXOoUXabd+FglVq5kfYYLBWNZPF2GKFCKabH8BKdKmt+mw7zo5MrwPhhka83WogdhV+nGE7aw72Y
D8AZWasgJVY3v4c71WHom1MX2aJtmT4PtG9shvIU9RLei316fWu6qPuQ6aisOYA1YfOilZ7SopII
QekVWO0XEUg5AHU2VCgz4SiX3o2eKH9oJFiBUYNl0DTIjwTyVydwTRg8aC1+0IOAOSoo0pKp63fA
pzE0JKT1U8AZq5mRUwMxkAzxKARhnqCzzRvfel/CAMxzWp5m5lU9I6FIUjQ3hpsrbw6Hif3NqYkJ
R6dx3eOItZXAshb50vWjWucC3WMVHJLYD23Ct3zNumY3YBvaHqNlBGPccpYY04XRtv4/AwaODPz4
fVgpAR08kSgoGsIZX5e/zA/7GCvBPAjrXV0rSmRyPZHJe85nV2DZbrlzXTtqXYUwdZdoypgp2jy7
UW9wpN9LP4Y11EddtsxuFCkoPEM039SwDSjCC3rC+LUbDa0HlvE6TtLlOR16iX/jTE+A3JM9DqCA
DbMowdUVY8Wq6oRq+aH5bUifTRUGD3fZYdt7xRQcoDjCfg56wYcLadtmAzFO1U70upZJvQ6wgh0N
te3aJOPoV+FkNGS2HV673it6nK63wZm18t6HpHEZWmZFH00lKgQq6uK/IygmTMSYc7/oQZmIlW7K
75gG2me75CMOAuxpLPmIamrf1L2iv/AOVoi0Nt9tlOhaBxGg4VO/lgUYc+cSu0FVjx8PX0jQRIwS
uG7w4RorTvuRAI5LVYIamWvr23Igbr47yu7i2JxvOWSDEW7/1qm99f1eZuyPeiKCchZUMp65+a1W
5Te0jSzj0HSaC31yMnuemLZ2UUrd2xDQMO2x3f/ijnxicsqwUbtu/4feMObt/zOf6STWM5HUuwL4
A5EElP5gCBD35t8/KLtoV83vuuI0W/PIbqlvsNEa1kavanFQWL3X+T5oUoo09yeKnO8jcYGWtdRE
k8TlbvxyYOIAZMxXmZIXJoVgrKaMu/lfwixY++FdY4V4sGMcXS8qd5CW2iuTRSy6EYTU2X/lHm2d
hTZr0L/u6GVANidwWt41trDv2NAVnanumkpLrycO7tr7+GhzlL6q8/7oJohOynP5t/yRgjrGRTcD
Uibry2HhwV1MVieSUAVuOFL69jc5kGj9vBtatQ3Lmmj9CuHSfX/FFa+mDy/G9L5/fFQ547XIgp5m
7Q/AJKE4yo6bcaw3beSz6rbYPXOfsG5OnS6MiBU0azM0JTOFcsoFPk1Y81VuePA0s2todBuq8pm5
PtZhCFzGn1IUzYaLs7zL9FM9C2WlguHaiR40omMHy1auJTR1sA9F73/vC4sle1NDO04KIIjEfXyY
7jaPk/RQQ07o+EAfsW6oKAefMPoVbvE8zROm1+W4I64hYXpqZ1P2QK1Bg2xsZ+lLhncO34ffs0vV
I7BHf/m469BIRPAMLAUdJKdFOc4dK7vyXZT50XuHd6g4Mw6WPObMTtD/nUfMNiYQK/2B0ofxMuyF
My9Ot9xx9nxrjYh9T2VoRs2kX5Rj4MdHvmvchVDyqAn5fzIi+qrAISok5wc0zZBj2AXyRvJiW0QD
9tGz7DqoxZyhge6JiAc1IpicBT8pA0aJHi/mBv5PxUCP8YVgCijIeheneD/mj2hRvuE49aayyx82
KgmQ//9dqjSxgzyITXBMasQLEVX6gP6JbA1hLujSqFJVHHtpV+G2h6AktA8onaWXvUpBAhHgwqKF
5iJq7w3nCmTqm2VVBKrV2iar6QXudrZfkpS5XohsXn6RaOZGSi2D4c9mkJ8pbK6SkOW1wE+Gmhd3
xiocVoUO3nvzqNc40kSJRjM/nD5blvD60oEi37tsUq0tZPatrCgo4JDHvpzckOHkpnvTrRO4o6uN
Pb4g44GkD16iKQoukFR7x/K6LdgLOaNYhxf7myqKiXzCjVAxABm5DH0iY56WMCRRgL47XgFJAi++
EWDdnK6+eqMyxpeLe07Q702qUjO+ykbtuIbzADxMIWoi2hpReBEwM3w99ZWHSyitFWBofJ+YZ6c+
bDGcOfhb62gSh7mEHuSUwd7MJ9gziQlTUXGT2FeQgvi2B8nla9bb3ZWVTR0ZK+bM6Gfk1RIXN9tS
F96rtCM5s+TAbQaQ3PfgtnJfrFxUIik+m8QmXcf/z+KpBNpEOr1RxSfFOfJYCSdS3b4pgjseZYb9
c/drW+fhAqvs0lzJBXFu/KXKEna0ZCBI5ltracHxyBZbSSRnL6q6O0/vZGAmLsP0kOyWgEQ+FQUC
9xtUM8Yajsr8VMoUFfLgvAORMKmyuPKPEsGX/PsvnjBiPInAtJu3cJj2NWoOhOvKzJpW21WTAZ0F
LN1Ja4P/N++GJ4LaW1re3yipAqdM4h7VhoYd0Q4y1H2WRZZ8wHi3Xy5Uyh9AzDVD/sphXV/R5aJQ
XfEH3NzSt2AvS/qAYgT/hxAHciYWknsRc6pJhOUgAbslCG53r7nvk9Jp+3zxMgICcZweLGjigUWs
benCSsWi0JRi6LWgJEu9ziF5hmbJ2EG797vHoMpEcaEv9R3Vqi6Ee39zBX7NW2u6SVJJLF2xHXVq
YhPfo0YTi3a0hQmvHv1e6Id/6eJRBIvR19AoQ60spb/NJ5hlq3xJb+jNcyLhDzcY37aC/XHtgLWN
fsJ3ByOAkyib3au5v9plq01CdHhZFtVq7A13smUm9083+mISY9ka26m4r4XlNfbmRrAYQULNXDJu
ADas1GA3v+g0+hk2Z4C29lxyLkXTjFKhdZ6c1dLSq5ICOo+LY2snkQP4Z6QqH9ylAAllLXQgFGpy
jyg/ZfjL32tXmeugdFrRgTB8+ZPsC0Qa1A0PJtrzY5floierpCVrv0D95v4xy4/cuvrRpkSZk8Nv
nzE8+NrY6nd833x4PKEBRXWif0uVR8MgmjaHS7XGE7zGZil6bb76qEk1krXUhkvpMIoINDEDjnbj
94DE/10Unigo7W1wPJtqD6sNpnRfdM6BoEr6a8YNISihkmPkyIjdxF0uWdmciN7Xle2tMyEbiwMG
dx+vYnYBVMJtaKe8kzYj+OYPHFRJe8n7eAggea4Pr91F5Oi/wfkiDbHlNXm/hwEbgCK7Rto8BY7J
QO3lqUce4qm5Rrwj6jxW2Oif2RPStLcwyXNZnxjKI7s5G5anbFByJyrq9PPOeZ2nHQM9sCat0tAY
YXzLueWHeAjxzjQJsw2ft3U1OXrkuEGKAqoM4BFBETrcxgGzO3ibbgHO3JHVTUqydUvwZQ1FAr0E
ER13SIjxD22Jlh/uYPAUj5ccHbWmj7tk7D93Spv2hwOZzFITPHGbR+e9OnMoWcELDrKoLgNlgvme
aJZNIEtUxpwzaplL2S7hNCqNyNGmkxON1yYs+BVaujle/B3n8lPgz9+vI5KjPNnCYrOxYHGgKcN4
lJZ2WoFDJ9COarUelKwK68YIqi1L09ECjnH2OecSxg2WBRYmrfS7H8EKee7hnl8GbDBWfdiN4ohG
iU9Lajm2N3MoAfqsIVR4XkXAexXSCeQOdyl62k3O4N8l857FFUidvb/z9SGf2WYOoU97YUCwacKz
UM299N2rEnoOGJkai6bPi66gm8q+Mg5q5Nh2KBpzpiwMm0NE6/q/3QTSZPuxtsaiNED/HsA2Tliv
aSvUXEPpimD4TS6QByWtajpBE4waFyMqT8YgW5EgVzpjQgyQbkq8Gzl8R3oj/6Oe4Vdby2wa1WtW
bqNlaTj3z5xa0Sx0rD6gMvPtVXjaoZy80MA+Zuea9akUk0m0RPBC4dV//kagAmGOAizPKrNvxFE4
GPmc/fBvGlLYf6LQIkev245AGbyHiL7Dago5oq1MdOvvhmtCUGmUY0z+H4iSQw1X2bXT4aEI8ZbA
3JJjQdW2mZi2/XFCoJtz9NHrNlrQ6BtQlYa1VY1DKFnIm6yumewFmUh08cp9HvES5JTnJWeLtsl+
Tav8hrfiyp3kyTArjLYanPtS8BnH3Z+r/E8g/Q1zK1I+DVF+ouxQBAdQm5Eluzu2997YZzoZHAJE
sESnli+cTKxBedcPfOF+iq8L1ls8VqaI333zPhonBA+22zvxoMIBCrTtB6UhNHUYNSmwjevhPdrD
5Ia4YYwkEY9lKwnB6O5FevLieXKZTvJGCglyXGQ7xi4oQA/2u+L1DDMSXPGEodkpR9hYigBpUXZT
BJgx1sDyHM8wBbY6DS1n3HHUf0Rw79epO8CPBWMyzNiprUBT+wro2SAVB9F706MwIftEkHZZeaoF
NPiYtsa1KRoJE7YGs1jr4BLcvtfUMn1HFJjaCoTEZaFGLOugTxmwHk0JiNT+WjhJJQq3Shhh8G2y
ocAnPM7D6KiHkLRIiEKsBWwlaoYFhhNtR9OzSxp09BSrQ6u/wCAY4q/O5gwhqA3loz+q5Ms9T6gA
vHX1rVyd/xvDe0nRQsByYIzEmbX2xeScUAKCFjNl80P+JQPCc/5YA6E3wUgF0K2oQHcNtM+YOcQS
pxmjTgYIoPfC1y4U7uggxUIOo7JVDM3RG8mN+Eca3NXiu0z5V7nCFtmJNwQJbYJV+vciIm6GfU00
uwpNaEug7+TWKV3r3bI5rYMsrFqzWllr0M1Y0SYfmTGqthX5/LzWPf/xCAmDWKeklZpCRlE+Qrmg
AFvNdG1EjQZPVq9jt3kE52REKPMZFl0X13My7iW0WN+yji4xH0oG9spZb1EZRfPDzfLCYP0WFjOK
XHD2RYDlBdyRsLw8oP9ucRZ2bRloUJC+E0VGfUMXrJqQ6dgKyQeBkjTAI8fqfIl1MdxAziNL6uIh
95gwufAGLn2BzdYho3J6lYXdWWczSKOgKCCowPpJkcXpWM0WnGoyxaFuM9ZqHVq0NOSBYInFq14z
LsWj3lWAkdb5O7nwTkB+LF5IliJIZOuYE+5QZNgCJOaxghrEWN8X4nQCauZpFhn0YlfLT1tORwek
i4O+tXtyEq5Y64f/FjsO5tAcfoWxobPKyUpiqtCMqKRMyi327hl6bwPNukUAc0+n3kVJ+HurEizC
SWytSh4e3EFF7c8S5DcfVFxoCRe8fKOkA3bBKeReVU7qFmXyXJO75k9g2YjWKu6XCSCc+5HRz4ay
HAXT/6EZWCIei2MEdOQDwuX5hGoMOD8MJ6Uix2axOcmq/CqpWseepsAJEdieN9NXbD79IKUMgVMX
UaWeZJqy0orajSmD1X009R9UCSHL0kCfDFC42i7ZvxDPQF6B+ZDiAooTovoOl6kJL2M5Vmy0aAtz
hQLz4i+JxW9T9aC2j1q9qxDvdlb0fOo67SSZ5/Dn8T1uHHTAFinD8qT1F6wliMYl2NIl9QFZbU4k
h49PMCZORNXe5N93em+KzpqKlbFy9r96Bx57SQ3gpwr0QdlTio1aN1umTKvvaDSIi8T1iHg1zCSI
0V+0a96QqE6obB4Kl0YbWnVjSVEojuZJEmLsJN5Rx03bOlIrkDi/ITCmgqAwcMCeED8iVvUjpg+6
SCG0cNvFSKME8Cypb/sYdWVUonq20FkHEwh3UFUHnu/Xst2ylM4PdjsiMFJLxCmKd2LwMfqzh1LU
EUlvQqku/+yUgHyN65pT/DKJQ1rVzWDSZlkZwxhpsYlpo50Lf9hhM2khVi3Z0uZnpxdTWldS0fGx
cB6XUvTc613PBZdbLZ4+qDzhtoS5CxAy4RW9aXMaS124NFN1zbwYLC3yHMANQDwR/+RhXMw+vBCm
Q2QBWuHPONTyjhTRpSaxnxjo6wlMnMAImDoajHgoaK4qWGFbDMbcVXH8hFK8VboEJIjSQn/bQ82g
uUh387LxGk4XWUz2PiB3g/INpAgD0U/FYbAa65hhYrqJUwB9/LTdOuNfSqNEu3Ol411Qf6UPCaZm
hr/W2QX/ywcWmY462bl0Nh9hdGdJzSuhPI+/wSo1ukB5UZz8x64DdOal6R2r4cTVUqQFCzJUVYgK
WTV912hhvC4Uq7BX2irFHRsPDa+tmxJRNLY3v1Qs+rprAifA8/GSZqJB4bzcntpHQutpPqWFgy1L
XllIb5040lYnh5AIXQKoMCOnIL/4H1mRVC0QizgvKP8kTPKe42Jz4HPpQt+ijJHTVx7MAn8W8bNv
2H7iLUgBPz43UJu1Ja/eNrsyMh43eqooM39O7bTITUNRtWcI2pcE0QEvTKYvSNaKpri/3SJJQa40
mXHc3vEhnqUqSH0DC1iPvutPQsC6VZ6wTgHhmFdS9RkUr2IDD/RezR9r1gEUGxyTKOFDQpv6gBDp
BUO7ZDTpqdd08UYj/un2CswF4OvTFLanttoW2Zgsd5jIGs398sX8iXpHtM/lnuW95a8Sa/m8mkGQ
m0kE8k8xhM5kEwZpduSGswK+UzOFo6jAAQp28UjiTPGLXL5sLFTH0S2LFDB1J9Bp0AVtUimYdrdc
M6lHRuccRew4IHJ7WKnuZfNCdsH5/vAG3PmRDAGG7eBOWqg/NGf0f2yw3Zs+yPi7tOuBYNuRpGFp
+PIo/v/bNDByKqg9UsCKLqwPoWir7mSo+WD3507un5W5BY1YEnFhiuMfXjG473UxBmXQJ04JRXuc
1VAQ8YZyrBMpO8Mm5yg/U1em6Xsy0Cs08wAhTozZRolEbPehhK9higyPw/OCWkizQA9P7GU3eXfV
lyWqJQY6Y0e/ItmbhHeY8+NySltVCqYwDwOCEt2IW1/eD65+3H2akGqSplShyF0nZf2GkDdAXRGT
ph0H9BlYtPrReUVqjfCKtZhUQ4MTZz3VFdfvvwW9fgXbB+vSkkITRKnxfIDpSYTp/QBaHo8nQ62e
vMhxnwkzoAuXD/A8PVRa0t/WidfveAOvZ8St+2MWrWzJNcAolQ+zm8QdOfqukws/Db5GwUfbv5Bj
81KYPybDFw5Bh+zyz88VlMKXUlfWPazM0hrymr5M/H6bua4+8a+/4EgNoi+21wz7JLG8WPE9q1cW
SvepfFWQWTxWGMdId0n6bEc0AprxE9Iu9AkgsGRcdbKK3eISGTC4Gg+RvMnbgGHBqxmDHDLrle0c
E7u3mf0SYuh08NxYPG6tu3qrAWP+c1AJ1B0+Sx4LZChxvN5pnNWRClUYYZqTmawXgVcja6htfre9
dA++OL5+Awh7xBsnAQCL/g3PlJgzl7jNCTKoJ/4OhKzIuBT9UttTtjrAot50rdUh0LLe44UIIv8G
j+vV6TEOkO7GNcWIfM0mFLKCIXCZJ3eKeuwFFKtcQ78Cw4gmdB9OZ1Bg0Yi4hSXQpyYefPUDAfLh
XuL4L/9GI7TWnRdBmYIcB0fEqFfN2Wf9DbzbXnPWcXssT36w5F8qDNb3Y0jHsg65Gq8Ke7MXpEom
A0R3pKUryG0VkCejmQAE055DXn8PW2nSHACwcHSBNfsP6ey3hXVzEm/XzOjDsJ9of5t0/jYPTWBM
2v6ggLPIo5Ueb/uEgO8BmOk2wU3DCDN+AZeu37DOGXH1Kj95vU3e4vtZhjD/JoX8plqCSOy9vcFx
6bU7MKNwaJMRZe6bRk+yOLKEiK5k2ulwv0Rb5CsKpXBRm1WZmPc8OGvCs9lNDHnKqgR3gEFjmlM1
v/LUCQW1wWV+LRZyq/M99HE/d82SZcGIK3C/Qz9xtPYHWyyBbzbyrmfBcXoFBaY3cNqw2wEPqI90
+JJXjY34txunQz/W8RxT+tYVIuFpMw5a7fUvKjily1yi77yr8SDyj4FUf3/IO3izjfpIn2DbAhE6
PqUm8T7+jS4G0TKA+muR5J/tXTtINHo/ClXbf/Eqj47/Mn9Jbt8ecFVuCxWMGuvqtnrzIuA1lXJd
HinilfU2DI2lj1w64Y70YQpDfPKHJdpYJw90F3ewS/w5QcAMfXvw+viQ+wYZZkI/ZgaXaiU/a9HA
7Inku1ZNNmxAs0112m5d9iTXKU94ClEWxYRGORgnkRsnaSUMDbR2VdgCrGGPh0L9BenmkwMT5a6x
hNh5OTMxCKOQxjEJGEAvURxnGOSmWCHlxYBfAcAERQb7W3Q0eF6xHnpqfB1svl6tfod87QBInW5c
lVKtGJa4/E8rtZCO5vfCqT08k2u3/rjMwv628UJu0e6WE3mc8x6dt96VtTasX07rCgIVnUam9gqQ
Z9/5pjhSwEnaCoNJgJUfQdSBknFVtnct3w2uyScPRl32LwAOJoj783oJQGUk8xSRFfNM7x7WmNxN
tadB53xy5++a96+yv9WdVxO3kr42LShTFsJEXmWwG9vMFG2IYI7EEje1iuuzwfd8r3zKUgDUBr/O
1G+80POYRykoiyOF7xnShqV3UOMr16HtAOIZHQGXTBSMb97rz8vdILOZ3aH7YSxq8kGYb3hrs9Bh
81igzLkuGtlldRZjGpQfyZZl7zkzoHynRLP7TCeKWvfz0qTkRu2WFH8GfnZdmYsLXHvsGN+096Bi
UxZTYk1T6URiq50mQp7kVo8UWoy8RICJI1gzUQDmf1NrTp/KtybwJFBsyvFBlpRmOM3mCb0BvPwU
m1mrzSIfbiDwIIUhCkvFTDwgVRLjqeaPHyFn+3ypTfJ2MB0GmrvKOEdRxQnzvfVC/Xb1Xt0Yo3py
OAeWsP3Izna6TcJv9rtYcEWHKAMnNXUmNxNOsPCSbTirejpyV1hR9oVkWVpjcuyTvM5feVnGLohw
TQSm6CXQsTEDuhBXXvE43QRQJBgJrQT5nbz2eLhZpL3A9qRv70k7VkypgZGfVnNynSRp2e0YtvtP
wccD/LRA3okpTEcgIOxnkJPOzzvkuxQZtdbH1v5cbi7N5w0hIO3ru2ZzfumcZRTPo48be2y7DakP
W1VR3hjJ0T9cho3j6bgldXbunN+DIejszvWzXCk4TAqtcdtffzPoddwy0xuePUo076kHpFGPm+tP
1XfUUqJj8tgmqomZYDaLZckEEggvl4EOSOJ+Gv2uqB3hqYP6Jl/XJVfnM4z6GPk52gHAMXFQCyRv
MjoshAZrNmI397KsZMCprAYMKNzzzaMn1N3PGRFP5yH0WiLsH3pzQOgy08v3N5FEovknRSbdT1lh
EWP6GCn2ENqCj8k/Lp/cSdC5VXkLXCVe3tQXt4JKM8KcJdOX5Fk32E2lAmKgAqV6gy7qL2KZXagp
zVtQVt5trsUZZ/af7C/tdbmjqngCCWOPdAzB35sWhkIu9VJ0tZqOOReVMLkVQIXCRJXDMTwbrMo1
7wCACw6wOZLMgo0sB3AEJihcVSab6Wlhr5E8MZ78R2bQ0BE6jdsDHPzWbRfKv9/TCAKDiGDk1o79
1X92s4UtWgIaGPQLA6rjOsRx2YYOgnZwKgNopVvb7Ygi1gsGc3RigRDSmtxsqypzA2S1j4+9xEsq
aq9dlDSOe9sQHgSv+o3VnA3YWvlx1ZghLz1M/Y+hAAit0+LurObneeqfS9WMkGSQ9PyhWhWa6Qkq
8zyBVKvmFUZ7+hcALs89X4Y+QkkXDHI6ycwmYr3VC84MjNrVIY3MTTZBAokyhlE9q+eZ5SlWuJ8S
DJA6NeTLPe7AJHT1Q9KLpvO3TZKvfije4cG6KzLfguFIImkgdp//a3C/2B5nbvh6+T6VqC8cdlJb
y9di2A5H4xBDQQqt6xvTdMdhBUq0GOVlcCQ9ZT4TCVFJaZLRRVVUD1O+arAafdUv+K3nyblB3FDI
abZug4LW7TLyF8EMePXPWcubmtumIW684yjPyjzS3AXnwilAVaZDocvljNxRyOA00RD+bDJXxfR4
cV0QHYa8rDypOgiCq4PGGlurNz7PC9jVzHYK4/q+dYnnPn9Mu+Ig0kI2wAwhGtCoUrsfPt60jDXi
9beLtDZGxJm+IkAaveGPkUtociOg5+G8akQhwUsvHJOgNwmrv6uKH8ciSsJfK730fkqbsF9JTG9y
HjUJOH41oRpa7tus1lFvMxDd2pfXF7k9rG+y9hBTsTC04v2cjOepRAfVkN9ynJ+FbrGyXmTEO1kh
18fC8un8iFWz706cKiCIcYcWCPnqAV9xgfedRuFjKhTyGLUKY4/cibEGXaLSvA3YPQQ0b9ulBMUT
r0Al3KgBCE6JPS+cqN4Yq1MJfZyZIM3s+9deU8ZTnP5arFOSDpjhHQuqCpivSBYzGFEtP83dPmwT
NAed+l8eugUP6FjDDZbxWK02WAmiMNf2DoGhyL6PelqCfrt+f+a8CPyfqQU/b54mhZ45U6vJvjux
vIJ1PpexCYXYEMmt175y2zsDfMh2jyoJnyAcLNnrSGaZ1M/ZBbF8jylGwexud1+bbEauqP9tMyt4
/YcT259m/IGCi9l0A5ywQpqsZlYq2HanQPZn3W12ZW2oKs3S2Z5FB53s8OIrZs67V4ZZ951r0yip
a+ZdAU8PhJhKw9OejQ/MWfqOI1qLJ1GybK5cp05P4FvMymETo5hYh3EE/pnwoBTMd7MerKfYfaTr
pGOwEicQTrrgOrKKXjrGNSv1XqGYSGl3xFlabR7qZxCrA80Qucf5IqN5RtFxxjdvFWu1CQLUd2qR
izaFdm8RX4BH7gs6ZYZ7J5lTwYFD7TA1B4sM7IU+efyM3eLfPHIX8wS43xMmI7n3hI3yCc0oLZAX
esCy5IxY6zQUqhNUQ/0m1g1zDFz9gH62buH5aKP1TwDsn2gQ8+PueTHkPklc3Bx6TaUasFbPtxsy
FfQvIzru/WecUwUnUqEZC+d//z7Yskq75broTUwROEon5PAXBP8K0gnxxVWPsUPiXE7DiER/Nuz1
OF2MIs4/BhsmHZd+ygiUTj6lWuXE+WwR+cWHzX+kHcmVWEyNNP+sbIUa1t6j8oL7tDaJfFhcHiC7
b9+wGIj28QXhtSTobMDdUslvVCPNtEKNIBBDywy0eDTOVUncnYO7LpN2FYu7eenNDSdjTLQBafNB
NeDY2+L3l9stanegskb276+nnXSn+m/J5XC7MizN4GKUV6Q8rcn16LqfgXeJzEG0LOkT7Yw8/L5H
2DKI0zskPtqc1KKTuUw1ukzJ0I2BVWms4pCwadoIS53qGwr/qqm5oLmHYLGF45FG3NPwfCEFbyIY
u+j4zq3KComQZn2Yflpu5LphP7RJjBtPCnUPT38cpvqQG9d6I2fF5PgK4zxlinX9ZynvvblA6Ohj
YZx9WNOqzpRxZ90QbUIsTOHgOdXmodp9w+phnAEtx4DcgzWLeSyRS8rPCM8J5MJKuAEe+49aRdef
vhxgdPr3ppwpQ3DIX0KAGVff9QTkZ9d8YWDG2kj/qWv1h0UpiE1vY9tn/elG6E5anlL10ti6/s28
sdWwYnwl2gK33MOj1oOr76rMtn3XtbUr5n7P2quARJrCYQIHOIxFZnuWR35o+MEb5I0y5Z0mIKg/
MCO9k/8u6ufcFpMX1BOD8lH+S74QO40CFAGtRWh3uItuIuH8EEQEuLZ4SFe7fjNpFa8CE+JR4SGd
Fnz4OKvPC5MSZk1UiccA+tE0ocq61OXIGIx1UFFUarruqHKvDqKOQNZkzzh9PqkvmdslN2ge2yMk
ojkiMh5jbN9EZLjjqj11xPOy6MeNjVzoKBO9PJyFkox5BI1sDubVKBbXbb5zsbHvYa66cXhhw3fI
oXWVt8aZKvmqo6qzOFPf4M3otvWEBmV/ikrGe1AQyny0WcvS6/GGi3JYYdA9wORpEW7Lyvk1pgCN
jcaU4iPFXWhVHfjrHasbsFQfheOCO8x7ArvLOFaTYtiSB50sFdLpg7F8ZUAoiFopnXJE5Z30IK5J
e968HKKVs/ygZYpsWSDpR7dtgXjzKOSJGPxfrTx6grKvWalmkWxvd/V8Lc+O4wLO1DIXkfMS/v0Y
mmD3OvDX8DoHq32e23jbmPRXKtWpvdDBltp6xhgzf3l0nXYC78L4ETy1FHiXgpzCY8GBpfWXSGMF
/xLZBLMWugpdktpZlvD8OlfT+7GR4qGz0ooOxwJgCc8aC7s6TV42d/6eSVhXvheT3k8aAeLb9THK
KFKG6Ri4JQdWQ1gzRvmY+a/0kDUijv2sHjFvDUO5phIEUihN/9vgklMM21RSyFTLxVrK6M9RmHoJ
TMqOKfgRWnGb67Z4UIS9XdunB5fPmnm5tcDv7AQNPIneVGIE2lmkn6rKr2/+/bv4lk00k4C+8leS
WzCs6twCKCIpGne3EtJoVrKnciGnzrTng7E4w5k+jKXtHtLdwTXLYpkq86QCWNICT04b8nt4/OjR
31WkkWUjTkbmT1FsxPgCF5XjtHChqlHvSt7Nv6mgQLbWDoT4VoiTXILFOzN++QtEQhF6shA8B2+E
0a9trEW+YciJFvDgkjih9DtpAmQNoE/oh7bgwaCP88EghL5JLYUWwipghy3kSZ1ap303Hc+I3pIM
TBXpCRiN2t+WNDU1axp6YFbFbmTBCzNWiuADAJg0mzWbChVRU63126TqvVDIgPVqC6cun7kKEm7U
QeB7oF01ZjHUC3mQVJxjSmKGojh6v9klxDYGBz2gCob3zUIPIwBcPzOyRA9/PJcYdMVvrTCs//he
zKI6pQ2kxEj78riEGafl/7SZZ7A+/XzyYLADiQYFfBeAfE+aj4jwD/z1cslQUDjktgiSkfRHNc0u
yT6UlK7rFLXF8KnhKRuuIAMwWsLmJ4SvhtTrHITIMl3rM6lDgjQ/Iu1hiSKca5QunD6mymD4gMDn
mV2S5dqMtuIXHBiqeRcAm2zsNCAoecV5fbOX+a08E5sAr2EFLtfRF/gkGBFgOySTmXmDdwX2aiVz
IRJTNSdYLhAft381WKmiaUTIFc8uJFJJ+Tr51JMdh8K8KExlVr2cE3cjAPWRgl6JmOt1NGicoKhI
06XSISch7anzIh2obg43HExrf774feOVaXEppW/W6xJzHwT8MJXNiiO7kXe/1M6NQyxvvv1GoyXK
t81XZnG5El2lgDCAZ76WdBA769sfQ2GOgCpPOLAk5oVinE6NPaRMvZY7b7pmip6yGixN5i8+Sg3X
ZRyYHlfVSonXMS2As8cd0HvAWhMvEwhr0+ESi9LYBvfIDm35ISBpZmOcInQkYBj9qM61hUPrzxlH
tP3bveaURG85uGiqNdelDzQOoG/EPHjYzFiqpF5eR9QFv6L73g7cIt/FzpIjH70jEKBI0vUSGRQc
rx+7dlg+YDtF6OQx33ACF/caNhGV5Q1cI0rPdEBK6MiLxKiblZL3Ssz7K0uHpGbZScKmCoB4nX8p
OuJ6IKxk7ShuEDjRj0uOVxAUxV/MqLEHhcC4kE9J8J74Bto6na8hyN68VkbbvGLJppig49d1jxpg
z4inxOv2Hz9S4bv4lXH8T8cT6Eo2tEA5HtTextVHhdfGlqLyNLOY1YoiCHuNV9Ph9wZsZcKb56lP
VUDuLlmokjmKqbE7Ta1OLYlxpIkOyyVWUa1DRiZgExOqpvs1A/BojDFxb5B0kcIoxjvhJfC6hnTa
AGqFc2ozAw8vU3w35a6UCI0SnRvfQniJXWe+75tueTNn1mmFp6b9W2SCwvg3FJl2SGa4Axx231H6
0mcUyEfdmWPqekYzRT+IunQmAgQ3Jf/df/ctWoSLtroDWua3RItr7Umrw4bDmAvCrGlgHAG7Ewhx
Z49CfSzMC8es2lmgPB70qIPf+BJKG/syY0RPO+yRp/a9zS3aWfYKjllVOkvMOmsiZU3alaTC4hgr
WdELLbI1pGQ2ewIMhDpzVGjpe2UwzJe60lR364P9GUGOW19o4ETGUfZM7boDoLcnfkuprKP2rHUC
74n+N1lXUSp0I0OxablJtLcSQ2I5Q+Tgr4nsNh6uREMnrZLwHCNVYAPACQn56X5wXjKKUuDPc2Wc
DcfegFRQi6bN6aNbXgkpdw89qMkd+/ZZ9Wg1KXw3IoCzEXC2VMZB40Hu4CiqsiRtMGGRt8xqyLr9
h1wezIC+8v9MKccU7SJ7t4Nwo1BNTlbXrkPL1fe9GNwXeaAKDSp6UT7oPGhyGfCpPPScpwiMxrox
tQrfX0H6KMd1kijvudaVLuf+aCg4l+AmNRvUtd7E95wgnOIR0gAdaOWgtjTSbievM2txlIdp32nt
brJkMDWPia6jVtiGuxYt1PSlvmigheQNnqNSlHOzzS8svKuzq27UnlxrkU/LLG91Sw1WwCtPZSU4
NmOJKDCECiyY52rLpMzlnAFgcn5J6ATdGFc3kbchekNIyWgK5fWdV0t5ZNdP69ki/LHRP/eJA5//
nBs55YW5zp3RR1/Tl1NKuSvIq0+RM+ajyjINf8G3N8LYrVEeNTqmp0KSFwXzj8ffejblwtnkEz8a
p3WAxZPQpJdwNBCgn7k/Z0aWJjaWyAhm1wIlSZQgzvcc2nGRxb/BuzFEvyeN79yGvRQc2YXu6tq0
afFlNpbYEwJjnJR1aLeULvk0dT+UEhpOP1FjEoSkai6LOuk+lYsxkIWRZVLBhk2mPa5NKHAU/1iw
6y4GVMaKGNSDJ4JVUfx/lwQXOmIj4CRFFUe12n/sOQleKPJTUIJQQJOpIkj/XG7qzwXo65utfr31
4HACU8hw7A7fSddDnLE+CEOtMY415AVzA3Un8xOlQ9Mv0RM7b0mlpVmwB97FKe0UJImL/4ugRbwv
3wD+tKPhc+yg/7mnV9xbzYaH+dw4k3UThTqeFHsPg+nNR3U8mJptLFkiRzEB25UIvddA6n5dNA3y
GR0AOkr0Y8syxuIBChrsSVKLJxOCGijjmZbYqN2Pat//FxLbNVv6P8MhiAukNmbnM/SD8CbzeSe8
/PMsLIj3K2Mcpo4OrUaGJWrlC+H+vVSKd3O33SUF3l5Dxi3GyZ6ru+Ky6x4QLm29yvreMNN/efpL
OD7+ptRPJkhoJDQIBQjrM/dYddwapwM1g5EaM9hV3F6VBcRGRA4Y4y/bJYdYrVWVNSq/s/gDj+xT
kwHfzGQcnvQAg2ukJWsPnY+atIXPmq53/YxgJWxIV4y37H/ot3eCXvsT9m7r5H15cwnujNNuHWE4
McRLbMr4vCI+09nzLUtvOEgLagMW+UFv4CPa361e9H7VUhdCQOAVEMVpRW9JaN9pM+ix9Km8WGx7
wslYs7mifDn5CKChQrydCbJ70y4JzF4ejbMIEclFpW9z4kjMsw1Ze92JL5mM42pedPvDNPe0LWzK
7c5emdVy/JuYwPl27n0iANBFu8LFB7AHvYEvkPJi+cEh4BeO78OGn7HlYZY5bcinEjpZXKf35a1J
936t0p+er9TouJ+UqV54Gsm6bfW8hORqNcPe74JjU/Rr/TcwRg2UHblNBrsVSMeKyV7Ra4L8PhEt
E8wMvtxp4FoVczLzWN3v8/lU46rnwz4U1uTkeuLsMuTG3wcaCbYOGImXde/j5OSLXaHELl9AQeOI
+/yUFUyitwwhhdJCqrUCNZQbqL73qL9ecGex9fzi1nKoo9IECho9pQ1wDPT/tduYLFzMgOkri1ng
Tudg8j8XyNUTQdMD5X/pkULYqbFcUReeFUTB0TGQeoiiJh976rNJDu2LUqRE0MhehfTDzJ2KmmW7
Jmg6Ymu0Up9YXQ2ZzBdjzBCVmdaQLfl4KRLhdRwS15YWIhICPpjEbHAtIELDqse2euB+X0jVmvcD
Voqp0m+uOGrtfPNV5iP7eOLqeliQ6R5jF+Oi5nlUCjvGSSDtzr/QlgUK3scyPJR7fj1+YTxdawF2
c3Lzyq4RuPXiCAr6NjbkcWb6rUNq0V8Bn+rJQzk77pHnUkb3eGWjr/V1QXxhx/GhMWaK0GqyvwLy
ylRG0VoqYUzw8z+6O/N86IjHdnndbZL733eypkSccAja3z0IDCNZtNbzZWSqx/z9p+mru6BX/vT3
5L9ySR+d1ZYPdauiQFRRfITpHbuvDZFO77N9SDSjMLL/nOywRbILr6EoUcCwVObetBhWno46bPfJ
bjS2UxwNCh9KNE30aljrUdXjkoZUlpxRbdyiQvS9KZVb5Ao12OnjU3MO7NxEZsk6amRct7VbXzEf
WLUcMr66EPCMFUSWkLcOAlBH2aiMiMNFco5ZWILflSZuuU3WL6udAbz5VBcQwRCY/AODJRyMTH9k
tuswDACEhXsCWP0uExszPnOCltpzl+J9OF4Y3a0g6HsTOgJOjMYPAQz5MznP+F4aroBoGAVHc1e2
Sk6ZWCZQGgNPL3sTH/8+2I0QGYpNSdDzWCh1XHX6N1pGhM804E1fL6DH8UeTSw7LbDDeidRc6AYH
3trlRUPHduu5ntT2+2Dk2E5MnvEAowKsnFDyIPYTNqEqV+9VAJwDndgKjx/S23iq78VIg8mLfR/F
UibqMRTnhcAGIyj8Kr2QptdPH1Nuv2EwCv7nAVgB3we4oLFjpxBG1OH61RUD76tS/6+FpdTGyonK
J8QgBG49aiBNju/cmNhVBffD6kKv3cufF/eOnOgOoiF3LQZhhqOSXYVDG2Irc2hN1quA0cLvSFEn
fK2GZZxMAaaTYw4eZKiAxebbia1/7T9DDLSQ9nHCWemqyabZLiHOzJkz4FNMG2x5jnKzkai3ImEd
iboC4sGXUGSTzLhfjgCIbEvCZFWPTlevR9njzRxS6Dq9jNPBKKZrYMmOwC5fJW5VH+cwXyYaryYO
NNqfIk5PxLowmGgI0tj+ILC+hV2yaDrFnH+wHnSomRDr8bhcU+qp8k3Dwjn8it/E/iVky/dt1sPI
hBLB+VaCielhBW08gdI3ltDAGezNDJ/OVyZ8ilk4j+E5iev1H9lTLwH27LzKSyZx2JxwuEj12+8s
Z2Sn7+40b2agQx3PTSkTBFJGdNtn9W+WRMiESOzW+XL5YPn764vmfAdEo7qP9J5iiNbAq/88pUZl
tzZIar+e7RMn8rgwrK6mtJNU/2hfr1UBe5hm3S7EV1lluHXcdm6ODRmjaSi5u+d8eVHiKNZObGpo
I2OOEooEfxn6N2ApDHKYOJVX2imum0H9t27nnIBC7159pEKN3uTuI8jkq4662k62fWnHuQ0p0EaX
avAi4cdNK2ZW1Gvt59vz9q/Mt3YdTsLmGls49vP4m8iFZPaqwdlA+2AmLNWGNt+BRS7T6Y3IlmmB
d6TtI4d95nyAygU+guy/3bvAwWCALqixTDWgcUDIa4QoklDONo06hbgczlAiYmDYbJV7dqd/xFHY
9IovzvjTKRaanswf/p3yCL4X5lteC6WJCFqL/ntyaW3iVM7Rk1JDaXssDzFZa08PisUq3LqPPr9u
ha5Qg38uljfhyNtPbf912ZOE6QgmMpwxTdvJn6ZIWgENmLx0Sl0oDoRpdM+JjltYAN+RWYN8XQWr
qstiWGk+Stf1JZto7rEWv/Hveo1ru/6DgShyEM7OPCbQBAh0VKFqW9dx4p4NaUY3ZpnZa8YPdQ7r
0QRXaA/9Q28fBhlIaL7/Rbi4qHlywzMszYOR2uF1IveUNg1MFdX3I3PUrRRebuhSPNujbz9IX7ob
5qbXPBou7cUfDFyZ3MU+keI6XC2OO6K7f4SqeZAOyLP0wgxfElOjuWwNqWvwx6UaP8euvMnBDQ68
UbrXGHeunxi4ddNZHUIv24Br/6jxL0BP3SoGZcSTLggZdIOz7NdeLdFnD2WtlGEtmOs0V+HtXARt
p8MTeV5XUj+QqR2jVueZa/pkcpJLRPHaDMJl4DDYwqPs04iewWzzGGjCkf3ddj7EJ8t4oKFy7mD6
WuGcVeVTH9FW9WSMcxeDM3KUIw8WFRwX3OBKVzpoTNSKZzoWlYxJKLJhJVl91xBMmbszWk+Br2jq
yUzVQ4ogtBjyVMf7L//XZ99kPdHLmysH+VeIJRnQ3s9kskHmbg0YmNxTiQ8WVV8bBSN0qziwgDwi
nfAwWriBvF9MbGSHrRZvSmxHybg+bbhT8O45HwKhtc/UxMEK8TVVkWI7VCVpaETl/Jn/+Zw1DK5u
ObWSzeBQ+zdnsl/h3XXcyjv9QB2hWxwe5DwHDjVma9mp62uHRmjry7ujikMGDaPNNQ+QYiEh+/Kr
kE9c5RxfTo1qWx2k8+C+bcJ3DbOrFOVr8e9O6zuVseWL5YdglJhbBT/vjq3ONYsecFv6ndkb9CRC
6ksh2GkAdNRzek/nnMl2uOG9cI5bTZ9A/MZLQhgPGCi1HmUjdNbjQr+2Qf75spJkdz0ofuM79ID/
0piPP/LJw/5jSi+2OHuCko8cTsg8VU/SXyg3HbEhMlXdtjDoRd5sVLU9/MLA2HP/1tC+ZLlauIXW
ILFMkRh4n94QH/bqC0WY5DUjJ82JtqyY8X+Q+9IiAym0KGfLDMRBgYscyRXFvZDqSzv5cSdHulzU
BNjvTpFFDdFQNZxX4HkiWuYuyfhaGQ4x/zJHdFcLjADEQbz82vbq2TmojtTONLwTpX6/jHpLPSBD
xM3w6RxloOoRANvinedu3S1CmabGUQxN82xBAwYMwxp89IQI2sLup+fYTVvYz8vn/KXSXmMH7ZzU
/dw5fbhKQU5eKcpcrR/MjF/tbppQklxs7D9ODJH6Z6E3rh3UDFaVw92vvSUM9iX3f5BnGb9D9Yb5
oc2S7Jc76mHSEfeiTSQhIrEFvVyfJJsg3VdJm19NEGqo4sHitDSmwIu8faZYqvncGUMviqwJdsuR
v3vcP2pKEQcSvWEG3B1HmzwE8BCH/o16z7b3ayvgh0NOapoIuqePbDp75b8eBCjdb7Kw8jFLVDOR
GKRO/mKG3V5pX7WCTrLutjtUiE00WovGqKS1ITmATYBfMU8tGJU4q1z9nGQy/hAKf7pj0uine5G0
RpzYl4milyipwfQRcOskOkTm/Vg3wAvenkmvjU7ZavU+5kffhVQvVShaoQGkKGa6V1K6DRx58yPb
E6EVRBnrV4XtNFXqYDZrRm58pvgOCuhbNzep98ra3hPJWSheyXTxmfmGhoalWVjAkAtFN62W7f4Y
QT/L/tnPl6GcX3aLO0LhRqPyADoKey42lKi8ClmiV3fxZilcXT+C4Qq3Wk98p6sUMApLNDr7oCz/
4sNlchXVe9mn0/9ppKSXTkB786zAVBaoTK6ixEmtR3zfdSet1CL0tc5E9wFTnedehwkpLpOGg+Sf
UmKfL8+eiP5VhD4lNfHxGSXApAFMaOJuMt9dutipP5ci/opoRn2V4anPXLQlPBVdAU8Fb8Txw44y
NJHl81LMSxKhJgRZRTMoxk3fDa9kBL/DrULuGRssgOZaHmldOgkriWBs22eMbdhjRvSUeAWGkxNb
/UhhZjDYzpNWMppXoHgBx4rbnSGp7tsowomnc7scWABOB3FrjtV+T6Zu4mvG/CIgO5kIwwB8B70t
AwmRpCaoqmbzzGsPE43Qpzk1SpxrJq5z+PxHVUV+yZQGpd/UZy+IAW4j8ObLeVZ4YNYFXbPV9iNp
AuwortsqRb6BzWy2yjl9y7+fip/EJ76M4MSFcu2D35+gAleIBIM7t7JOoqtGNy+QKdpEyFc8uuZ0
TCFhwsSYkV613zLQyk+LtyOxmCGwNbJenu1rfs4MolPiwDbbCoEbdzggU/Qm4S+KO1Ftlh8HCz6O
V6Et2T4w962b5kCtGJ3PdCo58BC66u+felnyzIu19WMlYLwoMb04pVbaWvZ7TLv/Cgui/6IwQdrr
Wz6CU0T/oeudiamuUKI3ON7uHr3XIjJsoVXrCs73FGPZ+ELUyEVjPiiZDZ9k8cODhIowkg5YYq3j
3jfhkIzLpLMFgj2IE1czy32vFZ92vGFd/4FaRmIaGr5o2g/JIqQXZTH4ZsQS/ISo+Q436gvMPq4o
LXSdpKFcpS1R2cuID8m0qJ2y3lSOm5Iwj/Z80TS6M6zWXyHiIOGeRI5D3v1OO4ivT9TxQ4G+pRBO
SRXix0Mcw14BtKjUfHd6KFaqcOL+hWlwwuoBFj96IcvwCeHsDT5sZrdL7s1qz1CMuaAicYUJ5hzd
u3fgmRq9RKIMgpFyTpsKrMz78Gyn3ZXp7pjKsAcbwkjP2Z7ZNtUXVCVoBSZ3kXyXFW9uR8fHjo/W
2i30/F7Z3/ujCl/Tu2MFuqcIrKY3ze8VLxR09CDjbN0NjmkzMglpklCLfJbbj6SofwbNSaRpt+Ax
QoF+gRoDGzCvfm8UCW0jQae3EgplD1rBDwVuw8GX5w6yuQJXwiBF5ifdmaSjflcohvIfCwxWnTuy
DKh/ttMjxsA9NgQX245RsqjBxWrOM/PH0VqLn7IrZhcLaWJHufasahgovI382voJyZPC1AGQypCq
QSRpEiDdRwJes/yfh1YtKNcWUIN2hFT46JxPJwj47VquxigOw7JGSQLV3jH4A0DPgb7Cdn5GFb6/
g6SjWvRK6rDmRmkqXPq2OxxPB0MQhJUA/9mmBKOymjqBsJzeOIhZLnfPwCcK7XsH9cPXx5JaBI4P
p5/hPITpf/9+kV0kUO3wyAUbbYd4xLsPRrgvex41aHD7uNi3lSJ9C0D24NHbiI+NzDw58CquoWU+
1/nRgegTdlNA/IjEnxvjuhT+7GjXEDFT2jP2H91Sqv9bism49yRAED9NWB2mqa5xyuqvWoKNQ4pP
wKpQyQD06LsPr+9Gf8FEdZ6JDJ3wCx9WvcYhmLvWPd7Nn4HBU6txR8gJ4ktij+7Q5fnLQIu3DGLG
sE6Q432rX3b1GrWtq2hJDPMd6QKoanlpLgXoJkdY9b1gq97dr9plgTEPsUPACzdMza1uTghI6Kgu
yjwkGQY302TTVjYD/p4SAU5CJy74VIqEkGNB7xX51KTlBlBeLdNPqcnk2yRLM1EeZnmA88YVwhMd
4EuYGyEiJxN2GkvyGKs9GzMuyJNnDG5n+hwogu/tZEbkQWIBcygbCfAH+mQ7IhhDx/bu7c1fVN3j
QAgUo01q3aTMw4wx5NCPP+UqxYCb+SjPsxUn3LOSQzVlpru1H2ZUxzVdwenund/yG1ORouKoXwKE
3opmGkh6VErMls2VT9udRDLDJgNPSFKS/emnfG6VVk3OecZiiw//idprhyuYK5QQxUOUbHWSYOdi
8v4hLnljQOs7HuRtUvHtyDdzBMZm9wms6k+ezD2gpiP9oCFTxJOF9I1yNbuAtfVO2TGRXeQyvEAs
W72RqBPSOqOPkCg1LCrMhMuL1q6NrJ0VqOws5tRLmcleVjI58ypGS8XRCDX2YNgWihXl2h9og31V
FffngAJjy/rYrwL8D4BhWH1PUoklArEpmWZwsjp0V0PXZQwUVdZe5ARDp9Y55ovW9/Uj0WY2tetP
s+OU/4qjeAh9CID6ZC+wyBPl1pSxNkr2/vA1H/03vEyrNaDF6Ltrpr5i8Lk/8a8W4A0MgumckE/5
PoqwDAS4fiE8Nm+D/f6IccG0QV8vajvEiic993FR2rKvZXl+tyIXodVpIg8OPNawAwefbpgFVzMI
F2JCQE2jU2nk/79tdoKZ2euzBB+FwxZsXbuuOris6pRMy39NGo6PR/OJt2vQpkZkxGR5wX1hqb3z
9mrspY0V2FTeRBUv+HjtsM2Ye3INMIB5QpcugpkbS3/U/6WTdUAjDZpvKO+ZW8GB/knt1SPoA0Xd
Z5viTB+oHVomBRWQFMoc4IkQYLs0pIfCh5Kqhiy6RgPBuNWwwgGjzr2kdgKH3lUcupGJ2xRnye7k
wakMw4w492nxgk64c0SiJemfw9rsO9OiT1BxLKXe9fXImxmVYNEXE+IKEvVTBtgVEEeJZjWpvwY/
PXNvmtFJZ09LCp4t0PKr32w+qJU/H9a9SHMkzlXM3JIDu7dHSwy49rpBbUuo3g55TUEq3qspQc5g
DkRLaPNw51lm3nWB0+Ikfi7gqdepdfM0zBM/rsAuUimTM7FQzuvfywt2X/+aiFfudmbztzc072kc
1rJ8OtpAYRzME/BewPepQXuL3R6irlKJN7x/+VB9VFXNJ2pxaXK0/NOgxWrhbfF/3wRdGFx9QWXp
Kacbh2biRRJO5J/WDY74GvBihC2lEZtwmnvSpvL0X4vNLXXdlG8BHCH6iK4grQlOTIWv7LJGGjYy
AE/YeDe1d6EamjeYLZxlMU+G5BNsBmq8F4VopjKXUHXZlkAoc9Ootm5Pcydlm62dioqa6JKzIwcZ
QZVzRLEI8cOhIqCsYapPeSDFbv2yq/+Bv4o2YzRJlsw2UbCifwkSOgnNQ/3IfnGE6El2na29FtML
dX/UI0sN2/shfAaEHD7pE3ZuSO2O41/9OyAMY3nyPvn7HMKgcP1fRjUy5V0tAk0JwR6U6BJ30F5E
GybzoCmTeG2Y1h69wje8K49STLbdTU/OF+7EHTX1ixSJD+KPJoK2kmL1pJZbVESg96DF2wMctPFY
fWLNCpNKYWZjkfC02Z3wnwXz+zWY8zWwnrvKTWg7JRa9K3dW9Revt/kAcgup7hTuUJIhGGd9sq3k
oXE307IBAseAQP5+UkffkA/RRJaDueokBaEr3U/0Q9pKXItLtlW6I7d/37kTFe21ygll9e6JXNr8
bPAI9HGn6xMshF2RyBsX2OaTXYjowu0H9QVx4F9YvFnFTWpe4sAFCGoMP8+TI3C90/ckdp0AVleO
hRdyw+JAsVX+0Hf4gJ8whOL9yXtr5FTueDPHChkHq8Ud/GHmoLItR/HowDCBtDXhcwQ8ZILNqHfZ
hnXW/vJ3yIc399uGsAl3ucxQE6t+WDCGoqAYjkW/0ewvzSwu6+Gn3bbYUD78f3aUk6IGE98Q0zUS
r7iu+0UTeSQuhHGVMWvFzkgrr4ROASdogCipzNqCvmWeRkI1+OhPv/9KvnljDVl6WqVamKarWTcO
HjFIyaLqgGAYgD0dIDvRR+Y66kVyQ04c4fxPH7E5JZdV+eElWxmtRUrNCnecmESGAH6uvtfSk9nm
sy5G6xhf6eBve8d2wpTewMlskmv8dEc4VBaw5y5Ce3x/TT6d5FDcGmof4r4IZYKxgErK8Z/zOLMA
furX7EjKo8g53vlT3VVm25RltcdXUEYBLeClkvgREcbSIaG4VWbUK/hR4S9yRuKcuvUor3UGXLZ0
VUbvvjN2KdI7sI2sPfgvPoTMnCC4o61Q7YZQz/Q/dxp6jRcgvbre9mpV3k7Ek3jpACpwrf8EP2Bs
CQo/nkBBL5GwtJzvUlDP+B8gP399MG3Egln+0xSwjEXrGmS3ZVyvmOeGG4eJ3bqBxQEY0q5W30DU
EuhhMl05Lx+n84uMa1NaF10mxVy1BMsK44E5YeXyRL/oeuOGrvJvF0hkjp7iY6PJLaCTmyzwAjj/
7KD3IStdtwhb9n+Ns2Ep7S3kxy1rG8R76a0BfZT9fOQJeDDhLwVUM0p/D8px06N25lxV2KDkSRHW
JMlsAt6GJ40xPvjUoQ2wXLvKGUMKfJ2GPkrXXMLVIcK7HzRNU9i7U9AJzrRWvB0p7CU8TulQqHKv
xgT7S1lJZY0xGToHisNPAwQaPpJzIosfRwMYcSCgfk4f6S8/OA0LaO3ZZHUO/+J1tgJ+kuGHGMKG
COupGNRkw14r1OVrYAMZasb4Vy5/Rz6C4740U7bg+f0RFRPx2VZgJ0d9DFebNBRIYxq06uZc6qfd
nqdv9MpLIeY/ACePufpAI3yVjrChQvu8Iteywj+teQ9WvbkNmmrBe7+irXrzfZfE50On5WBQD/K7
Si6UDNlsZFSFMfFHz2tt7EpvbOeazUazieyNqZmyTWfaTEwXmfOQgNuU2t7ps6WMrY5s6hOUJvJn
CdbDlUFu8Kxn5MDXXsF37hg2wIcPf4kX42LsaNlFHGl7740eb0SZKZ9fx0v++EHtFTY7BPvm3Fn2
EDFx7xzivuJ+Z4MZdsrQQ8HtF7ipC4+gLOHbiBIx7J2m8EBv8aNn/Vi6czD0buqhUcuheEkykAQs
FqTEqg6J7c9effTSGiBTyC4FBN8haHHsjAMAkS76fK0XCqUp9wzpu47hOBHyKrGjVHDU2atlwwv4
plNGtm71vs6wpmrfrQAA37xh7Bqu3YqoRGBB2Fx5k8rj0DgJwNNhcl8vh7lco8DEJjsyN6wKsGct
vHJyUu6YIsC7kfjzTrh8ha6to48YKIDon/mqyMqzbL3azI3G1ZOf5Dtg7zleyFqRUEKU+TRuiYhX
l5dX5H+5cbjnDtebgLnclnVWtOYjPmFb548ZOVAitNyGhB6GyRXFb1As/Bw4hwlIex+tyqpGLz8m
9bFmEpbiJ18apr4lg2YqC0v0GxR7rGbt6Ipb5eA3FV8HuyD21+T4lCIC2BJawJJeKW44nAd2jLSO
0KqT9INFHgL1LcnzacZ60+0vCch2bnX3et44qk8If1Vrky8mXPG6lgLhG7P7XgGb9sFJEJs+g9Cx
ad/DDKamdCRXq5M72v/nAUFSGjQnhNtS3B9VgqwtrV6h8XzZoQFOPvwb8R+HGxxigXcNkDtS6V0y
robIpgTHO5bC39gZuZjpSL+aNXv95y52LF/p3T3jh/BDk506cEWy8TSJ07C1TMZdQK6If031KviW
Kw+C7fGWXhvxLNrcRTsug+6Xcu6QuouC050hpLzDDbR6V9JFDKsTKNgp8nW9LrQ9ZRHRYf0ACM2M
36dRPdgkbW0P4T0ENdZzXSJkggHf6kCLD4aBNZ3uwNMnPj+A6mjh5E/j4nzxih5laS7r7qxlTOTE
TPsx5URTr2LXFwz5Q4HtM0zSgdX13namWQLQCeaGdCid3fMYhPaGvApOjA3r6ATAaE8PVVrrjo4K
GqBQqBDbRWbdFhYqM6K2CY4lP0bSh+BIsKHqfCduuKN3JAi0Dd/xHtIGAd7v7ysDgSty3r0jMKZp
AdeaHeTZ5TtrZniaf7jKTZOdBIL2esnrYImFuirxP6TMcV0JoTfQ7u3trFmMK9VDpOSg0Z1n3u6l
4jIGtWiZZBqgI3+3/ojoFBGAyXgVGhk8EvT44qre4DYu4Tq/9OfjkQR9wmduptk8TeO+Rmf2NGX7
zevwyda43ulyoeSRHhISfym42wFJ021kBm54dTzCV0eXUv5q7CEGQL+WhbsZZ6LuANmQVt2Gg8ws
4pqduFAwBTdA45lm+HVF7oN7OGbllybWvTTjMVEJJ+p/Bf93lHTUsWCuXQ5KL53qvVFQOvgOfna5
KHDxUUIygrsSpbcpu6q8mFeu9dTOWMdRGVSBAd0v1w+nit3wybDFVMa+BMfrv4SbXeBPD/KhWlas
NSSPTkOqpm/FRE+DtsScUJQrC6jex3TFVgI1diC9eONLaCBYBXtaSpE2NDZQrF+xYpHvfR/dP9xz
ImrtIW/YECOGoQHkLiOJ5CxwtXvxJ88jc1PqJX+84oiIAJ8MzSub61soxPpb4H4CmP4cNZCsepo9
sxjjX3Oz2dzJ0Gcmj2H/GiELT4unaM0jxvUpz0ro5iGy+drfOogdRZpr9/Rfd/ckbD6WL+MczrUa
n6I7+M0xYhWJFpY/mODaIgLyPhKNGPA9YeMS+NZkcMJpNPAU5281r81aVOh2zMC7t/3I+BAQDz7+
KetuFvYAW4jbQWYDgEhjp/y3TiDCjkPLZHFBuzyn1HmHuJQZ65zhK6G6W3mSfdbq/2+jME51hngu
ZNs0URvib3gqAlU6bHtL6gyvbEqzL88h/MXJvPJtiAncIlvUAlcoPjlsyL2uzl6BBUiSCBfeKtLS
6dh6IlaLwTBNKDa5JcDRo4Q8iQgpW2cwISKagKHvmcaKbmELEqMJpZiKw09r4kmSUYmb4cF97Tis
68PUMxVpI5BmslXQ7BaqGIaBJPO8QJBtbgSCPlcuBVQZ8h7df3a+hTb/KOx1poM1dNb0a6PGKcMj
d4LkYIOPp3L/lEEWA8XhkkbHbrD/571z2pRDsAQ7ir5abXnQJSKLb9iHLgohHy166UORgCIfDNe6
XJW/e8bxrD7dIblRlSY5ScP7M6//bZzPkph2TcPY5AkwqVtGMF0BGZYGHgkG4DpKxB9AZwEVHzwm
ecnUQYO8xtYzuqkjGtsr0InBnrtEB/9b+qvzEOHieMAzGmxljvPqmsw9wYTcgXo+DHIRvRmrzBpX
gnUry9PkUQLe7Ztu6mRjDW0EpwDfOYs17wN25dVkHpxoS/d1a7G76Ue2ShZXPCt7MwAoE7XLJQnY
Ri31bjFIIrak+cULf0s3LXqY003a+AhSDhe2qnpU5JPyP52SEknmYCaDX8S4XrYWC0yr0CD87I30
t/ck2XVronPSbQA3ulqS/ts6ZJHMHMLfWFXakI0TfeAkfFfrEJuxqcqIeD/1zGJr8+26rl/ADGN2
+HIPeYz/JWBqBLyG8jAXCIPhQN8A2rvlHOLR01NHcP6Nxy6jPXmGDE0cPWwbLeSCuA7wiOl4gvz8
5+E2/2EBNNxLZiVhzoXNuWQMFpd/1+pUQBTbSab+1zh7uOdloaKUTzeuj+pbv+OZHkS7nWndJ6br
CdnuBFaf3E8sl9id4p2CBXnkbJRXROTSIBtPVTps/ckZLNiuAAsUITCmUK6AiUyYJ21MVfXU6KAQ
2PnmQWbRrXyILFaFWpFhTOtzUbSHV/70aCiUdrzqTGVqa2wCy2xdv3PbxFjbBM16HKS3oQJbASnY
ZhPmNKAGtX+RENUc51KLVP/2wm0/1tt3wdAjJTEg9T94t/sMuAuWQXZEReXpmRqAXxEnRqMIT9nj
6PSYVmmkn8e1oqRb/uC4t+WdQQHqLE3vSKBJzSYEbTnbPedNaXb19LrkDIvTMzcYFKV1+L07Izid
NMa4RSPjFdCRPJSMizsVFD/q2npdCJd6Un9Y5kUlF4LGrf8L322HrY0A1/y4v+JlNgpwgdL37XJy
JCwtXb2mF0DDPK3FU0NPs5HmTWGWppb79sSYsc0ekA0gEZXTVqAKyT/6IQE66ITchJTy2vljz1gY
9rUJlCcn9cDwCCgQWo3bsGw4CyfEgz5+km6t8D5n8tRmZTXYt9taDsdhrcZ2SCWgUEJ8uONeJHuv
NS4G537wvHzBYAtfJ6n4F0oj2ks3GqJCCCvkHs6DghlTc+VW37/tH9fkZn1GfHsaWJyN/8p3/PEN
9p1rqLFFNOCmmx/lyydyOukSlUvvv3DYSiq1zlP945sT8LMPXGlpAVlcKwyR26Km1A5AboDC8IMp
0E4fVOc9EPWUXhFC4u6hwIgkQpgE6n/Y97R5gTr9ukfkMVRX6tHMAaA4KS0CSUyPbaMpJIYKcbO+
Vhw95jk4zJcgmk+5/XV8rnZ/HBS7PbGm3xzkR97Sj+vnXIvfPjOzi7WWrGUEY6oP37Kv5Z+xF8j2
gWiki5RCAxY3vsMxWhH94l2Le8omGWt+CNlzeRr6g+AqkRvOpPPqtP2XOb4hRD+PCsxWj9BAgU5b
GOWjfUHjbB2ob8T3VIv4wQULLWeaOng27JpHRzsc9bo1i+h1rscb3kgb0OAYqr2wEr/pM8fSCC/E
bKWJ/7erAm1m+XIj+TjfxpciXycVjm1mG2gDord/k8LcCsW5EYkvGmGSeDyAdB1qo5j+7DxOUifh
PlQlnlIS8edVAAglQKDzWAV6tFY2fXFrfge9lFhfVPfrFwu5Kzt/3HLnJQzwHG+lYAkEka3lDssT
yzMzbynSDZFS+HA0p5oATSJ+/dfrPxK1zt9WqWoC+o4SKRnzkHhHD2dxUvvqUgaYkyBgQsuBV3V+
VBvycnR8plBsEB6KVPpZWN5MJIOa67vSSLC6QJbNt5RWoTCQhUm7fuzWCNg2SgQ7T6I0MWDcV356
bJobU3LJtPtGMTDSClzT9rrsGAbPsqOKuN0RHBqXX6w967HXQEAZx2xyO0bKHEAyYs13Et2upiBX
1EPhv48nN7lQU3aI9PFIkKi0Lbntwrr8vvC8wVF5V/1cl/RXqeQiVtvGPpd5Vcl2JoDYTxmaKFzl
b/imhdHbVqUGjeGyy6TH0lAyGqZXO9UpZxkgFPkXcK8rIw4Pcv2JLsB+ykTJzV56nzdeqU3DQajH
XjBxCLe+OQ70RmivGWwJgYu9zIHhYM0++ArM8P7GXg0qCfj+2fcMnDhTgA5npL2yM1MgrMNthwzS
/fA+ZZ4HRxE72OjXrMY9dO0ma0i1vtbYx40LJpo5y7dox3Xt7f4uwstCKOxeelZqx/jD29/X7u/J
ALHA9PvbXEgrXVX9R1k1AsX73d+5FhCdbZeXwSPCdkpeVR3m00uiZapIF2fB4dwNsQjt0flIuMFR
3+/2CazYAzk0iZza0dFktGrnjL+7Q3TRWrgS24mEpla7Bgwn4xJK0AEGz//dTHDz8VXzGa4uEhqO
nF6evBVB7K/tn/prLcMAv7rUzAHVJ4W1tWZNLZkZoFz0kYclNYCfP99HaZCpngNOmhglRlWwFWQK
Tmjkaq9Z6S0iCq8fKuFJYQ3s0O/b1ltdmXwVaaWoq8S6Y0IClYrQ6YfwZaEr2F+DTjYVyk+hoZ+l
qESoai9p3KMqG0hX9E/SHFZl2uRmlKtm150sgonNNZJd5PxQkINEre0gi0Mc18DI5ygiYRJlTJjG
r8s88ORjXXotXSa/mEF84/JRg6flImCzUZarctYZa0kpb3d1i95d8a1IkEIjEkt4mXtArOUYhAYL
KkFKsG4p6dsWriZbewQJkwQFSEhFV4PzT+lBk6QHsqs4l4F9dvZk5QBmmFyIlgRRD5u2JkCg45Sg
hZU5kpRp3qtwmWBHyd4TTrpaDBXfJnuDyqjlFiQ/OuLHP/GzUXdjTjNE9VCVIOqOqpVa19TRAoBA
IAK2sLMt+nbTSM8boC3Zp2A3WsgIlUwqRzrVXWRer0mjDFwA/WKPd2AqjZU6NOJoHEATg1aICgLS
sfb7aiIdVomzqxyThV/VbY5X8FmIDQqotRk/QOnvwsyks2WD9sdKxz5m48ELhDXOjSHEjMcJP5wU
ik36ss8z0XBT3yBir5Bf4sIGg5dCdl4Ib3kQcA9b2JPdP9qewaTsMHetePOpB1I+TU/ETND2D71G
o5y1PHNMAt7wgd1aLPSmd4WZnTUO7znJADmDM3lgBl++SFmhgZiO0R+fu1bYLB13dMaCTnFY5hDZ
O4VzgzKHKC7lDYVcCuVIynwMNrFEcFUr2xA6Ix99pSVvxP5mRSvd9sEK0oxmjlePiLJbAQquQgRU
poWLlKZV3xh3LD36A23TsGZoIjanhXJq8f0B1i2i6e1KygTJLGDvdAciNc4hDF69VnzdZnKVNsLD
ia1NV0Sqq9gQYMeBNNjps8UGz4Mh7tNMdnWRJvl9TT8NRQVyzr30U3uvTnft2KeWtBwRK1XtykHz
EqbZ+MhoGcwcyeIhDowIsaSJGJcWC4QZ8gNryucAsyse3d/AW5u2H6gZJTfIxMsDQL6YoGhXUAqB
F5045oucpnwyIwEMgwuV8pNT/0EhRiJfpEGq0CEdfal39u0W5aTWLWjlesPml2kq9KNrkok0j+bJ
lrcozPFMT6ghvUFdEFH99ShWimjLhq1QwfIoXRZ9YGBLEHVE+IlAsi/o7gjIZnxjr+RRdibKMTzo
t/fQdUzR54wnBAUpFU71QgEas8oU2qyQfwrWVXjkXap9l4fe13IbxtHzHZm9wuvtjU9RuVTqd6Ru
zCAWrMXZz4nt4cFspqplnIoBTIvdO6LuUbKL9BKs+KJTgZeEnSTNTWpckZLg3mwiRDxIxOb8MxXA
BjO3Xuu2uCr1O3k5+xYU7Yq93/ggIDdQSycWQdvc8yJnX3tns366IDIh/qiQVw0WpHcec1gSNJwf
l8JGLMaIGBPN0qKTbBAUGIO7DYRKLWdU1v3ZmhY7EZdH8kZMbjNen8Jgq9gFlG5bCixmHXnPxVI0
yZOFKLbwSFxlIB8FHkopOZqAZitii5kHGDnpJlbe3UOGcDCBtDLM3oaNSxrHTQLXgywBy97gcQ/W
zTLWBPQBA6w1DZVi3IQt7oht5r2AFQQTM5LBTGy5jYu434zcAfQ8e136YrQqAxQyEbe8lqmiMGv1
+v/Dy+P8Rp3CY2NUBKEYpEqME1BPsO4iLLeFwq7NMEq5uFAAyTo+omefvdatTklZxPrLU4ZUHNF1
s23DpbW2JGUmGFHNXX7Sb5Oe0LgliNnR3AkPbkGXUdJVXKr72DtPLeB6fOn+8lqZ3hLMCLYU1iit
wP18T1IzKoZ5gORb7yhOVYMdWUNMsKMEC5jB8BfQcwC8KYkVfX4vAfZv7WUlSNZ4iDaWxxx45WmY
P0yErnbQDLnyOHPfXbr9iB9fDw7wEc77vTtmJTDN5SIKO680Sc4Lr97+hs2bXLH8XTxZaTikw01P
7xjHveKeDFfdUDxAgbfh5X2WskzaqZlOx+na8FwGnUTaW8ty/uVviRPBElUxgYehVjHg1peJ5Bu+
48KvwvcxvkA8xP/cWjVWBBED5e4rkbxC21dZKJG24c4JmfBsevZv6WH3TY5JKBLCKeMbiKn3vEbi
OHdqsnlE8vGEbn/hATzt93BvNbAgoNbvv/J9y4miNyZP7BX2oIrQKxKFmBGNlXuGRkv1QQAvEcVq
jVc+3OZ7Mqhdk0McGZWpcHZn1/h3LgKpAs3xFG/J3prZ6xj6OTxoHr1aHD9XiO5IyxknWseJWfjV
t0I4QNur5T+MEroRUbSZ86J68xB2hcudmBawSJeXDjkBbPbJVl/gz4gFLNPdriTldKBWcdBCFMhP
rtmhIOZSK8ngprgRrLjlcFXnoxAgDt1pS5fnBeiucNTKbmIn2mzhKUau0daEOLmpm6BJIvriUDgb
III2mfP4OFlPAAcR4DN8nONGTJwrdzXf+WXmKTvTD105/LH18YnzfSc1GoVI+ETZbqUMph8L+Y83
R633OBeTmAxHpxDixcdIsW85jH4lrZkgUqi81g55i8u07DwgRbzhpQ5b7Jn7UlA2MxMWvW5yF9O2
zF79zXQBiKcEF5mibqBQoO/AyEM3QohSP2J6eIQ7h3ZBgM3RpIdNUTVGmmnjMlP9A5UqXip/mWDM
fEK96OSvfC+Lij57notmeXsdV6p55lv6x+aswmrymtNRkzfC19a+nLk/RmmY72M7tXkQDqzqikM5
qmYEAMa7B6vbTuMDfwIa0V7ifnXVWl3/Yp0df2ZftRY/c2VCmb7gVpLkyahxSOFUgL5S40ohx87c
aYDMnSZ/HfBr+nTDtyff/QRnOvoQx1UGsnoq32SHq0UDkZBCIZIb6L96axGYjYkdgrg06g/trT4y
WDRGk1KMmsMbYtvtvotqW3LbiVfvLdHcW7HIZ7/INq1cGbamecvt+gXrweeQbFSWTRrCnyFPuedL
i0kJw7qZGLnnCO5gfp9vKrohJw9QgEUPi+IjCUVGAdpYZE6Fi9dXY2znoPh1llSTlyDLjcWEU3vK
HTPD1aQWv8GeqC+V8a12dl2/KPdjzivSthtvfEUbmjvdA3Tcgjzrvhbf4drfiXfMnZcZWpN+n6On
uRtmziE/HRGrS1hxb5qI+/ifYPM2brZl8ognjWksvWH3xwpr1Mct7HoiJYVTQz78dej5IvhQ0ZW9
9CphLhCSWOBzTdFFkefZSXpYrPbVAS0KDXGIDB4tHV+5aHX6RPaqwJH7U0uKI5FjPLrCMJelP2NA
ylDMqzf7D6T1i1OyUfHn32OZ83bWgnS++0tbQI5tG1PhNevSRER1MDvkUU9n0/l3a/gzk3/EUBtj
wQw2mPM6LzT2gX6ZuOpSAw8FTnNCTLbnSxch2AlZqM5d8q9HSeBMOXyEFYLuSHsLSo6bczWtL83+
kZfNBed/9GraGNiYQfNAmStK9rjvG7+N2m3t/b3kb0eMzgnYzjP2v5czVFYb2o30A9M6iyPrOkgq
9Ldxh7Ap2h1n7H25Zc4defPZ8GoTqseeAGEAKeIziXB2tHwyF+xgDIKStuTjEfboleRbTk+Xadhj
XVurUyiU1CIlqc6kpuDfyUpaeJKBFOLgSM6TT/4nr1LwcZ+SOv5GOo1XDxKQqI9BurvxgUYqByXz
rZ9u8Jsism9lGxVy6bRyqer1fnvxPL3tbiLJjimCDqQ8T/tuYG7emOKZ1PfSeio+htgs+VHBpABM
WhYaSkIbHomawhj9aWnoVRcXTwMrMTq8PZw3H9jOfU6Q8arXZvFbbdalajPmO0KFxS8hElLWStxM
4ppA7MPTlZYwnUd/SZhJHFUCd8AJ8+fOo2OiC+ZrRUcsh/qFKhmcCHbAHJit+5tL8DYlmZYs2Hbv
WH+jw7WcixNwKtCq98e5qp4DdKuaeCwRHHau+e9/E8HGyLyaCx8orcgV0VNOsREfvwdbQlwq0fRr
j8d51lqT/2ECjbVtoaee1peNhMGBxehasEDWohNALjkTwkRAO/4fSD01zAYc+2xI27eUBoo8ik2F
6gA8/0OG0kODTY6oUiCN5Giwu8Q/9ygZ4CS8Iv0fGqq/k7xDgm2x58nQicEAjmZV7scg2NPCWO5/
y0YGqp4tlBS6xwOwWxPDbMKkaolt+oZ3Y557KVs8JjKIGJ+bguAJDRa3zInDDFrvgrtQdIvaEc7d
7fGIxRKrZvOkuS++HG6uLFIjjyz98vfwT+LyKRNsFWpy+DafqmfUKoGsWCVGS+AG5BEwZC+ys7Bo
gVUEVAdjJnAncnfE3cMPFkXWtZnISdO2imQXa6ciZigGZCtP8J/d2Mk623DIpE9bwEcgSpEOJhPs
ViFm2dBsQUNh5m7CdNhNirrO3DWQPeDYz/up934PuwfvPyB+q6riKmA/YvtXAUwlgnPyBwu0ZFb0
f98Y6sXOVHaI5P4JmeFnFEM87kepJzXP3kVT4qNhq41tzKN4YBGVX2RLzzko8tO+vjCFBa8ddR5P
SdbopFZMEkASyFK8QwWKJvOlpoNtNfI/WqbKSXjldOE/uFaa1k9bfxYl2BxvY4NLvzOmOsVeOL+L
Hr2Lz+GAnXzOPnPN3XGs0R3wHiArJG7c/h0Bn1UtSUh+NpiDoR0xb+XDrVmdPbjnMk272xHxYaKa
ds0os4cfN74r6h3/SoZ5yCyuvLnDeTrNpRfLl/ba36ayl3FKcfSXh0EM4j08ATcKQlULueogDYMq
ZQ1RPNiH1t/Cdc4Yx/AV9VJHFR3okKMwjht6cPBy7A6FgP4Ap3356Ldw4waUoQQbHNZmotdAZMuQ
YNTIJcFWm2krk4VbTRWLr03SDpqDLez4jyBTloa7QP96feIuIF8ameK+CtQbEkCx1XXLWbU1sXXE
jaGiYvgQfNhrAhiPcAybo1Xopxk7L87y1vh6upWR5YXHyHCVs0O4EmqVo6pR37PEYGHjr3l5KCPZ
yoRNnFTKCB0NljCyvZdJuzWPnnIiWGUqLeOvMlZo6/lwvi2dnXvjqJjLDcQboom05a8wbugeZ0PM
3JEgiBSBLRIE7u2BUPu/BpZ87Jz1Uy7q9Bs41amvIc4dDa3TJuMW2tE64BtynnkJSbsg1724qGIQ
dSnHGopVXyquq31StK5mVuZuZe9HYVQMxHh3qT0mYhAL4Ggj+CIFDtDzV1BeVF/2NRPJzmevoY/c
DyL9PwlLaX8a74orRGHhpKCfv9jQY3ALPVExiTKP9ZEGt51PMJ95AWo/6FhfWbddAXygRpZdrp0l
EPlGHdGI6QyQcd/vTgHkB+Pt/pWJoxc82oYImFkyuRO3Gcle/0KgZRu4RTifwVwkdaqfGWLjbSqu
M8qG+ecp4/f2bLlgahYITwnadSHXlEPfm/H5oYtfT6N5YpaIgGw21nS9OzqS4nX4Znh1ItzAwU4v
6j55zyU8k+d/kH658/HXfVfHyrmMygI3ZL7g1wpm3OnIycBiA6ZSZg7zGEbJlh6ZdoggcxJoTBIx
fDtbJTY/Ze14tRfycIMn/B1aeg7vnIJIAFhCoeBmIvNXeMbTnmj3IxP84qNhXX6WB+mJRZSY9thD
nwJZ2fwyquEunCO/OtZaoot/hCefLQMOLvAu3r3qnKvoKfup9XqI4E/iD6D/j6H6C4PJ1yurQTHC
6Ax4qpk1eiz/fxFnC5nRc13mM8S3PGXsK5VdT22kETNbXq8Ldk9xPsrugDR0OMij4+n0WjmnMPu1
uLz28yLqFNtR6qUBLN2Oug0/sB65EL2jIAobhDE6/N5XgvrAmpw63+mWuSPKjV7dGvGq8MjUw+qu
VFbTDQmDDwlGPmBmrnA++X2xexSMSovGvTateXwinuFmO+m7lWrIRPV6l2buGN26MAKDfIuGr4Fa
pQ45BkCRMpc4t8Q1nGWdh0sgfYZ3YHuNtuNHneaGWhIKIgFTFJQVSyPmNO7wse7DYEd7VpB3YPEH
Qz22/33NxiLaU4smn1KAKchHO+HKbJktiRGsH2T7dfaWGXDh/rpuMcbLXj7S6ajSHbB1DfFUVFHc
E2fXQxYDhEXlLFMDRzKZ9jaCcKvgFIYrzQI3fdu5QVKow1jAoLHmn+3lsRKla/JXP07zRJ0WBzU2
jmSIi+QFG/qZd6E4j+G/SkAQvjlqKZrrPXQUgEDUDZGqzJrldcdQl2kLIYtmwqmDa0R6MzBT3ECP
aIwYp4rZRCHn50TpoR4YEz0yy2QjzrnJwARAcRyMNrKFvy9K1RsahHvNC0Lwx5UjWPNJq6lopVBm
3Yd5feMkYkZaLDMOHjhrMI48RewHie3ULpP5ANzd0c3fqRLS7oBKF3pOxPk7QgyQaarjDp2VF74o
RCggGsbKFYoYwh7Izh2J6Eq4aJ8pb0Y7yw2CfNtnOp/uGWFdGBDEFBF5TbYffmoVduqWify6D4il
upEVUKfVLzRVJFSz3dXHJhm3iKmK2KhvNtM8p6esknEtelXHKOacjSDh+Gk8J1PS4I73V4/BmAP7
ck+OpzCMpiSJw5DsOOrzYw5QdpJR4MVk+MZ8NTyAvBbkVx4DVBneagYwSbPYKq+KnCrD0wRB5gvN
4EdFxyJRCCIwU7bpGobqrX+WWMi7jCakS46CRvRM80UhbFikgdCLByHSTSFgF0xQ3SBgJak/oYrP
Pu/yuVzmysITckDfefR+sLTm4ZNv7W6fLsOpzYGYbHuyrD/trqfCSEc0uWUZ34/FB2DBtIGFtIPr
hs1P+YYXg53BzlyIDhCYz53pSrtaYYL7PQl8kv7C9WOvVPtKw+bfIINrTLfGzyS+T19rcDzgYnDM
hqawqpXMsgMglfw3i65whT6wFIbmKkqylvXn4NrZacgc5GBzRnULdpYJgBrxdmGOb4sOFD+R7lME
Ll9A1PoksuXQcqILHwfV3HTodZ5E9OGDsn7NA2ufk7XsfsjAu0vOCnposDpXF20Qk+U9FSSjni3A
qvOrHnG0ASe9mXMaFmpXzwjx7sUPe4qv6fqkZxJKwH4m6yPDiAvyICjivMGBFcCqrs0EVxqc3oPV
E2xt4rbmawAbd2+2ZiUQeMFrnbBGxNr7KL/xFNeXPLwzHumBBqJFvJKXx/jUcyUNV1SmuDeHFkdX
XeFHRn9Jef1WLGu5SckpnRhG3Ni+M7i+woFI8fO72s7VkXYO++vjyeR+Vr1WFglNnCWRZUGYbpoZ
QF263wahyUoxUJWjtauF12hXoXHnolA8uGNcORJ58Df9/v9DCLnZLRO8eKbVkoId/9zOaP+7b/Uo
cdkih1NhyBOh8W2tElZRcbli9ecY0YM0h1uOQDy5O/xnDcRyK3KJzqhrZWineaFC3kv/Aw8Ja0R5
eSHgb88AdEoqrPh1WR58qrIse/9s5zZdKRUB4fkQWBJxhtPAiH2NhaAjG8ZMO0pw8+mKJNHVgKG5
FFCUS0WocLFYXhOtx7/IBvN17Bn12+QoOVyx7BFPXtuA5Ei3bnMNw6SkI4Ml4kfK+YYV0Cdsngdl
TwwwMQ7yMASdBnBWOfpkcLsAl/I4ChJM943tw0bCTon5qy+BafAg5Kf1CG3LQrqptvsSkXhUz1fx
LAT+C0blll2C0fce5Xyqy7efEIi8gM8JohVMiUN6Y+qThqzvXYL2K+/br3NOkC7Ysqq3N4k1MQdN
G5qUepe9ZfHGsHb64Q8TRWq9bvhlphjKWDO44+dJJS9uSinv09pqQDOdSnzzP9J3RV6Mv8zwkoIY
Eo7FIuiCPhnBGmlk/iaAkHZPOC7csBVRNUe9jT07ySREd2MTPikSrCfEYamxdTA8TN7nJpcWG1wt
+1Pc4dplfLtdy7KoR4970O5Jm9xyJD+UzfkpHiSqBVfbF+HhqlPjhsoTIZGLQjW/8yFx2PiYASeJ
VSp06RgjUxiAPJgxS90WwvhCCc8Z3Wb839wGcRYumgyvonnbGDgpX4a62Lc14I1pzKAYaaST09gv
mdNducrv9NciTUbRrEhscx8vV6rUS19C5zasqDTCEozvRMOxDWOD6Y8H8mLXx53wq2rLYlqA/iSU
OBcPg7LBOh+W+t9dl994FM2PS/YjHjDhKH6H2RF1271BkNh2L+zC9Qbc6uuYoY6MEdiEqmZbXYnB
ixqYdBU7J/eM2Btiif6M7OCBhldHJKXBYS2H2fChkANZpsGZ3TonWXwR6udZz2i8mPXom0DslrAk
ppxEseVS1OKILFBm4iR/Z+yvw4R6PX9yTwuqLJBrDEX89XtqTVWZ8UehK8/AH8Vt1TTvdCX1Zi1W
UCivnRJcmmoZYj/83rhmgSQMiqz4QoXuHYdb/UaPsaYlB4q26msZU0tpWYV6XdqYfsVwFDzXH74d
+7SFaeS4AUiraybBoiUsVyJHZsLcqjBmP15XGVNay4JR/t0dXBPpB38h0yS7jB8IrsCuPQ/lp6ac
6unBo8uFG6gJo4ljEmCV5AUMcdEnHfI+P70y4sjV+7+nLQMy0KogIaX6rdzT8g2TQKtrLC/sQv1s
EWRMTZF26f2EL5WF8K6haqIHADw7V34MJhfpmN4NbDZod9Tj+ShszXra/Pc3iiWNOzfI1xi5gskk
aZE5nZlXR1ohDWPCY5AXagWD0oFkx/6M61x32w2Y4mH5Pf9Og/4jxJn9L997ldHsE6yMMZ2/B8BC
femK/V2S3ijk5Df4ISnVrK4lOonpuFSehgFnQLPmg2wKoFRxR2wwRYiNasRf9SdsEg7lIg5uppPM
S2ovgZu0yJHxLhkeqLOh3kYrq3CZ7IvCODhLmFG1Y0K9Rcw2FYriiT3ml5c6erba2I8zH/8BS+lN
8dBFJYK6rnHtustG8GNuu+cIKmHXxVGfLofmLlvhwNfQLKX+B5xJoeLdW7Jrt0jl0B6Fq/zNUIgc
KsUAmRfmDyp5dqaB/jFIwjMnPX02xoB0KzyzFjh9VHw9uZEVqRC7mXW2RAV2CBNJNOIvzT9KLn2F
pGrqlpGwrvdHNLc0SU/bQAilMb6xcZBpJM/LwjVCTfcrrZC6VndCOIUQfMhme3EBryIWAOtVwRoI
yJjEV8zAnToUDOqppkfCQAj06jtdbHFONegteF085F6H1effqAdtvUEcsv9rj1Zy0xQeePjYhZqP
sm1Ro1/y1Z5dVCli1PesRwkgRn/b6KbQmRRfefrG6HFODbWu30klFlIrEo+r0wQsI1j7ZMjixEKT
2Gcgsvg6K0u1XSaET/RZEEk1a86upbjo1CL2kgF9SGmbmYlmBT+IS910v6x31UC6FigGrjS3hUG7
EgsKjGoeKHJbYpqD0iWtbj0EpYy/k4vLU+ilDNhW10NUxt+dX+DD0TZMCqJkxHaPGda5ofZpFbN4
mAxaj1mGwM/q1MzSq9sGWum805/2rDnAzcUPaR9a83r5RFa6AKkpRKB2wxCz4BWb47Rvp/BWxIrF
Num6JU1R6MGqpdQKmrISB+oJ2Vm3yo0bGxNrVKTnIxLZmfdXcrNOdPm+0xGRMHfWzc3CqUCquTkQ
HAoVMTUSQOZMqQO6re31mt9kNTfB41rYPHIaqap+qUm6d+/Os2QI3/mqJaYzgJHG1rVGk6wt6iuW
UUpqSISNKWObuWyCICO5RcYxbMQe2XXgK5BBIew1NuBxfnvFxRozYW/ykqV6tnYRGOuLkQc9p1qP
3VmOHq2XcXLEt7IwUCi8teFrl62jfYZbiEIiK39bgOcksO1WkDGO0I1LLCLAPc8n/fs31YgF+Nbn
J9ZmCWli4IKX0a2K10Ufd73xraJT8TeEjT1RMe3wBqf7wqdgzGCQDnVGsGhaY7LAW0Jtga+ep74+
0sHiKQ7UFlPIqhSQWbd1pmCh7du3EUOG2tBMrWfdqC6uI+4y2BUrWMpS3Vr0Hkw5DPQdfFRXHA5i
me8Q5zK/vOdwfXEGUMiCdFTn2fCnbJiPJM+QOdkXmPxyJKHaGcnzvRhLNOl0gEGnD4GJiwyCyTA2
lRSPDaVjCp6o4De7o01rTOMCPMewMk/jaNdHiX3NzQrTkyb9SUQwMKamnpglK1C3lLnxmt1KlpxJ
UuLQG13lsMaW/4flOu4F6UMDDWK82iLLAJGGRMotrR4xL2XuLej/4MsCkZi31PlGBLdXUv7izXBo
w+cgOgHI9Dl8ULv2VDtbYzff4ce4jPoOZh7CWZrsFzTb1Qz+B7P6qcPTCGSYY5L0GvXtm2cSVY3h
FnUFrunmxPBYyiegXhXPsbpL3KFYlMdKUg22KBPuK0cEFh+OLSo4utvoclCXZNuSavB34HlZKg3+
/tOlTJidFU1BhOx8RReyL5Uz8xZ9HO4vWSyp2po3JQNGHB88frCHzgxYqFZqGA1ZQEqXJI7t7Kwd
9hT/r1FhHD6yn+yqI9eWIUXsQl42lgVq5XdU3ZDACX8Lhb0tQU9Cq+R9np68bEuVxHu/++9Z3Psu
4bkTuQPfPA+dUN47usztiL1ta/M900c5otWp92zAIegE2MC9KFO0nazj1Y3IBtJS0qmtIvrd/xyq
nlKBOeUKBTw/uHrkpWOX8RnvTUnBxtu0U7o5LziJaYQiIkN//N4BmawUHnCHu1bANCs3BDSmgJqQ
54qVnaGXhrC2ctvh0caYTWbVbgBu6tvn2rwTu+BLJRxbEi6XhgP8k5clQsCOocsOHhQp9HNDtPTD
LVVCsVpHX2TyYrNNsrWe5ITa8UZmmWY3YY25/QKnINaBO9V3Hdbnv1apufllrIjl9/ixJuOMnqEo
moFCu/RjesAI4rNgeKvLowTubP1XAB3PzuZymY0DVyHdXq8yKictS2TbiaTsJ8+NOz78cKUGTspS
AZH87XeluZYeHVLxqN+SCt5KeYZ5ip9e40945k6ywOvbc4BjBqBDJcfs2oqWN5jmLcDhEOiYLnxA
QXq/8IOkyFeiNFrBx8IHFFwpYtpQDfAX8pp9OithiKgkFM3LOiprm912gEFf8lvPH6ZT4WhJDRyR
Cp8rOd5sQT7jghv3TVQDSDlXf6uqeDsOVLju4GgK3aWpECOKiSKXSvz8Q+tpSFYAGV0TO/aMfSZc
k7Eh3nYAYjxDfzGEETjKmc3gFeRbY6ytnokrNuZdPuml5a3EoxB9EjVT+wFnJmByx6iOlXl+bjeT
9+U5AHpabz45NvMQ/5nxccfStQACPovqWae3EehowsCHfz3pIzMJ4b2zd4yRy85vJvSHMH18ilMO
6CJXF5kuDu6g49B4FMWka6TQyetH8JTwVb03ECmhLvnRuwG3OIAC1+E6wSygRogVfO8NEL5kh4+K
UpLv71T2N5tnG1yJuVOGdCOYeKDJE/IIKO+H6l8bGU/LIaf6kJmkh3pU0Frp8aYE38cb7LTKjRJa
R+oQK1izb67KvWQ9RwbGSNi+9/U4c3j6kx8CbqVxrUTEjEAySq/lSXomoc2pO7sxLs/o1k+LSNTu
ty5VOFNc1WDAXuyykfBeppqutKC4dd7jjDl3QCpRLg+krQiPtD3umgr/Tq/RnMq7al+N5+2C2fFA
BuBTCuZ28IBKdsap9gmMrlSS2g8Y3CIzEYVFVYTIlIbK7NXroRuTwz07gCJ8uQY9jjgXnFH3+CVR
JVrWiE81mn+8xq8Qdjbis1SW78X+iljgfuhMVguAVIdUuTNing5QY2XMLeoxLta4y7rSfBVONVrd
KGxu5f9XvpSIeConpNpyle4MXcHfCsJ9L16+Qro8KTiGj5RdkjbZg+RKAIE6OvEEUOYwRakVDsoQ
+49bSB/uaQFHzTeZ15K9XoWJssAUm5rFKMPFf7wYQffDIcBJEUJcscWBfs0XBEVDCoW2m1O77fTd
72czLOAGPFo4eddby3fKhsXA7SedY/sgS6qFP/EW2QFyge7X8Twz1+7xyksA22S2IkwL9sOg7ez3
k4fYu0MnIam8K5N0wb2qy7fWZFH15Exxy06Xlo1bgj3yTdJw4qsl9IHb1KUFLE7EvqYTh3Dsiimu
1GMdL21+4MnwSKrdJGynBADLMxIc90VZTVmgZvU8Z3ViHvqAE/Klz3ddr+o/yw+GC6v6mGwVzE5t
S4NqzGT4Bd3ShFS/PBKyc4h4tTykDx8mdHGNPMffG2oMPyLcdxXSVlDmiSpTGLcKHNCYIdPGS9aZ
AgzwNJWLYZlJnu8M+pSCpEx4OUmOswkUivVETx1FH2YhBx6s8v0+4fBbVl2KvloTPP8BxVtnuIix
cFf40zQiCVfrXeyCjTlVwWw/BfF8KFYK4strYG18Pu928XqElwDI5pc9ftT/XtpgBkC9xdOBsvdW
s6VagW543EhYDH61kyYcgkMF9k6Qo0/SfaLw2uqtQjokfrx7qVl3BNeXWe/jvFCeIZq4JilRA0qg
mH49NhqUWcAu7jyDzVOm+Q2j3uJCTmDZlFCBkRwoRbQODV5au1bWgrKnPfnNBAiD75DkhTOedTjy
oxnjL63mnfcp+bQrWlik9BZnu9Ijm8m7wSkOTxPoyFtxMhPkz1C/h9yrwzk2J2pmxpnaCXT/FZkK
qwg7ZXqxPx4pGT7G0cNfpMsDwNXOebBzeHhhIFKySLqrSqwQnv7dT68HvNLRr83wta51kF5luKfR
rrcDMMAr4cy38QVDXwDIB/K6B/nP5L6QMZGzF2wHLnj6ahVmKrdpErvM2Q0bbkb+DUHx0hcjwLQx
Z3NhXX0StAd4EQo2vsLOdoSvuMxPZiQU0qkHxt8jVydCrGHZq0UgYhGrRdsOgwLy6bsmMTn8CfRn
fyxBWpUaPWEyvFnFavg7tGLhGm0cT9L4A2xxCiXx8zN31lbgWE+l8eXXoE34O3v1V9rHLFAe+oyT
PaicmTHP9QYsmnc2uRfL6G5h24L6Gz0gv5KudSN2b0Fq39gu72QILRq+WhvBXAbg7vlVO1eWksie
9FzXZxQer9ao6GN4WBmaP1dckr8BuOMaWO3cpIbzyX7kbqpT6MT9xYQdbcjDLkI4I8LA7cqH/RUK
5o/TMNhyaxVbHuHD8+7u27LWERAmnWz46rknuRcjfghrFi0RD75jWhQJQY0SIcwTlzoRgVk1vceG
zYt786Bu70TRIu9dMnHYBhlSpaaOHvRh2Rpz6694BGWnxoANGgGCoutk9feLz+MBV2tjpqmsA4nD
YPTpZ2OXmQ+gJqbVeCeEWWi7IK0b9q8KqD+RG+mUPI4wqb7UAOEni/DOtGH3iWqJb7ud1KxTNEnB
sK1indKD6DluK3LH9OFWh4Huinlc9EEb++LIZVCIn2bSDDGw/oTveJs3OS+YHO4IJi1i9pStDo0r
vMbhl/PDC/j+pHsGEFF/wMo4LPv2pwSgiIlNzhf5Vea71VRb4tU4P1mp39hFlaUJXFZV7IK3LlFb
o6Cw+XaN4vGYubREkJ49AztbEVp+kuzXQHP2Sg1PMMV4EL1vvh57mabgyB3lUhd4yDr4phdD54Rk
exxmxM3NT4yRPMPE5qPfjuWKaMuConoXE4u1lm1O2/R3W2U6YcXxQFa9j8dpUIkFFK6kwQoe7Qhq
SQsEtXw77YvRGWbTmoVCo6PvMuZwKUa0DRle3cE7IvoMF4zO0zADOxOcUBv6dR4ZQGcIymjJlBzS
H+nrzc7NH1c6YzZHVGMEwXlWOxEyJJDlqrJfTxcBQGMJwxbh+hKT2e9gYjLryxcXKmLGe/bhp3Jl
eRbuZVQDiMe0HydEWAJeROrdlClUGbybBNoBxQJSEDAUPw/v9jlRa8gaITfStB6z76ChqQre8lJs
+xQ/5jujIqjGdxdnLsLE6A+Ynu74/cfiLI7rzCmk/0duS1kpIzszZu5KBDXn9GYFvwvTpdN7UPOw
L4RknlVPg2pXsZ+4FKxpoFfJGxAVM/053xZbCfLJrINQ/Wx2yB30yereuov/K/de6+wyYvCoMHUd
Zrq9xzEPROZOfhQ1YnVjpbIsZw/8L62JV/nqMBRyx9GnOq6mVKtal6gyMdINvmOcdSem40uSVnk7
TwuZ0DSvmWNPFBVWX2QqGFHFA/VLQdTer0JLkZaw/Iacmbx0sqsNFY6TImLfzddiM6rf7CxOWp5k
nXLL5W2WtoiBQaozBTwHs9ZLCIfEemvDEhZdiIM/dji7C5lnVZya78xad7DWbQVgApNsRNSS/W/s
YqMpfPVRaqAGdMUXrTeBW2dczaLIDl2Fv2vRVhX7CXn7RGW07RNzBKGrjyFE5RzcGL60+D6PNX+M
wl9aCJJeRN5S4Zqy8m30lCy9MbXTZRATYEA9XM0q0jcFcBbi4m84GWe9Fw0Oc8N6TXKK2k7y6w3t
sjd80qr1EeChlaThY4i82qDjEIQqjdQM30eDS0Hus82s/xY4DJf3/3O5+vUMah/d0kBC+SDHPf/s
XpcqaT+r/Q8qfQJFUti2nh2RXQoVZ2iyWSBN/R9sFrk7x0EISdwclsfy7eUeWX/C2iaJtUqLHOWy
JZo3kOi5WtH2AqCySzQDgu2RVxYqXc8K0mzWMlzklr1/U9YSnvBnkPYuGXh0n0i7V2SmDeky4OfP
Nm0FlA1zp6s5P9YJ9uWAP2GmiIIItJWg5dXkRA+zZWEI/LbwrgvBkyVQrHFUFwLQSFGs+89BFnxm
KOI3515ZZMdQCze4Lrw9Gl29FTpZzFfHYsLStP+JuVvefEuobFnmBpscS1NMkqC6cT1X3nu7aHhN
pBro96b4iJ5/eHwXKj3cxWpXO4Hom/f5xXfJjWn+fblkMS5csz3CpNnfvLwv7yGJ8ec53TOLYq3d
hiTYRPTXFpNPRsLhA6PsaVMlRzkj9DDjlM+8kD1FRK3C5we24uQdkuyAv7nWDTw0xJoR4QXokkfi
Ts+0UPbc0I0c7IN7uQaH6PPkW7r4XLJNqf7XQsZfelpHirZArQPWCAx9aEK9Eo3DD5MiYsfruIVz
J4HmxSU643FpsmFbhhOoHfxJnnjNhUGY5LTKCRPlGpmnEdfRV4MS3Pw9nBUWWcsXKeJfBal+Ncp/
hx7dePn6fwCBmcbR/bfxRlJBSv1QLdXgQtveCrnVlgIbupdl6kVjykGUGasu8vF3kFsSlJsVmRXE
UCSkyCrg6IKPUqNWx+We0JMBrSxzcDVxcqZXNJcamkHeTU3qhY2rxTloO1QYzK/wNw/QdPYLNg64
nymAirBB7p4bSlz3N/rHD/CaMXvceg7VBaDSSi09LgzfaeGWFCVAIDY6QTzF0QpXi0MbxjCLUzrB
A8sUNi5V29BHZ4/IOxfc2JoZwojQj5jEgCxwg1tRP5YEoUnmVRyvbqS132W1svThwFIRHMSQ7Q6B
vOq7O/ONg3sB0FNiXBmThxYhXiVV6Is/s91LGH/r7ZT6LB45vb4EbX97aAy3kLQMbTbelHYCKc6M
n0fp8x1AgcRZqHLlR/fMsKL2KnKgVVuzfa5C140D9wwkWESY+oeEP4qcX1/pwJbne9uU77pvoxKL
r8ywrXTlrrfycgO+vmgRMGqya/1QDTPq7thBW+OOWprIxN0Gs/ZudwjcLgH99dLRmdqpKZbfNIxR
dEHDugqSXujKQMyKHUBA6FSQYXI9RwUUdKT4e6p+bPHFqQSvw7H4l9v41xDriNeVNRualEyFl1Ag
Ks3K9O9Hz+LBpAqTA4O9sWXrJSxEx+Z+2A5KoxGG6HV8zUZeUtvJnevmo01m1tKLEF2PoSn7Orl7
hxnvnfC3rrb+bU4ZUgpDtqkTkWqHNj+A4951OHjJWJQfy+wfnwb+ricVPWsjbIfifYOzfZGiYt1r
r+4DveV5G3ss/J7elVttaGhML7rDhpUnCET68RCp6RNmkLjojl8vqn+DpzIgsb8SIRUqCQJz8L1H
KB1/Inp2gvPrlpH0oG1CUkGGEzShMN294n6/1W7kVGDQcqrBt//UTAunye5OKC5b7RfBxpbEr/+w
1bf5MXc8ybVMWDJoCQmrNp2MnnLjIZlGQLeyjjDuOlp2B++b4z5I1ERnTHbfHqap/s9XCbYx9xHv
NsaQtXyeThIDpf0istmhh/bUuoZkh8mwe+ar+TLzfvkfgjcNfbvRWyhlzl1/NphF0QTCDIcRbf5F
xtsUF8CgMxxJhnidhU5QJIyzSTv8wzTuKrAex/KtzuKw1Wx1ZmlVpjZ8oFwRv8s6dvKTmgjzJGms
5MFEoXDq0R1xr7J6Zl/CTas5HgeQjJVGfjsmeZz6G6BKBAv+PTFHeOuIB8sZL0js/NfZ2+UacN4a
Ug4Syxx+whNO33EROWFt39w0AD/wEaI7a+bKmZIs/KlBLfBGSu8bWAbdh1atd5D2d8VhYDuLYR4y
xx/J8FXUDXWJxq/mjDGB3mp2Ba8QXhhZIuIlyB6EV+XMRb6LOzBmzlAN59YOB8ePS8x4ITkqhogo
xa0GSr19Wkvfe2cz7pFtOsTSE/JPIFOyADizNEP6+ICt3loel8l2hOBIifWITiSBA7okN8zIz6S+
wLWsBGj9T5JTLsD88MZ+raElgNxD4REwpHWF0Sg09tjwzVkhkUNuWRQgym1jKt2aNB/kylpS46pa
0xKeKDwh8GEEH7Ghx3NsxpG0PXiRgACsMUl5wcLpi0N1rCEUwu5VAgxdT9C87Sa//XyyexV2dj0/
36HF+bQkqBmk3ZIJOY5c4RyKhUGeEI2QFdEakg7ntUlqqL8/0TVfTW4cyc/V8h0B1ExNdU6kMAO+
8M/ioZoFMLbOWOWnbnRiJ4S79INFVzOhYDFGA3rENs2T+/e4QudLLHgU+UtV++kpGXy/b+MBR3Bk
vFhs/mTvY28POOVvsGpAF6zd6wunvcISQ0JBeyh8QCAkw4jp3W7SZ3Jl6z0mhgm8rX5gqDZROJAh
MDwuD19JXIMhaySFZTZtH/yH0Rb15UAXmzEB7reXkeC9T9vU5HGvAtBmmgdmWAXFOnP8jBQaDKIn
g4EPrdYi5W7vcRyi3txUtsJozRNjh48EIxn6VnqW0/BLzydIqMS53dKUsCK+X5tTgUll2FUcI+PL
nULNEgkNi6jFIAgHa2K0FWFe/G2ExsSAqbN74hRcXNpgq73EyK5bXyL7toZOKZCqJ5A5GysQFTMN
B6JFBqc3usJES8bNfdMD3axnzNuEyPfy681IPA5x8Dj0IF5oRy66lgsorwPNdv1x/qPk1FIc5M1m
H3wTjY7AuA8HLo6E/eL/j0/vGylmPVmBika/dVTwmcqa1GeX/+3AuHVcxZ2ifae2QiYT/D6YjpBk
E+VdYlwzINzc13btVnfVwtMNsDfi7XCM0m2z96y0LpCddzsnjfaFM0gOCBWIR6bK1b9QoOB5MweY
KKm0AHzKDOqNY1L6M5mlaHasOv3A3HPPeylwzNUZKh5GgMaFJZDayda4xv+Plk5F/LMzYJSc8vQq
tjurWTttZyGipoGz/b9yYtOrzmyY0sfplFphS4cHvXZtEpJ8lg9w5vvn2r1aUZFxmjin49YN/9KF
q0cIQTjpaafH/QdHRkW6UV3tUGnC+QDCJfN4+Aiqz0RNyLOCbevgqpzfboq4QwVXz4JiUTMlI7Ka
qWTNf+X/rbrk2v9esWIbl7D+Xdt4XQTJeUeGWxmfi9WWoVjB0aK5Imek1+XUfm8ppK+szoI2sLK3
ekKU4L5XeYnO6Yg2hMig7U2iCICMIWPlP/npLQrC3lalAbBWEQ2Jd4TeWGnNGtUYowAr4FprpjcV
bGHKMCRitDspKHEHZKNtEnnTBS4P0JQU3zP/DVfBJdVmg5Ur84QK/vYku3vzg/QkAtumxQsMfsuL
tfv2D48tRo3cRNiJMW6/ZCZUNB0BklKQuXV6Mk2iXOz+bd+jOUHmqonc73elqfvVxUpEPH6j6Cu6
pOap7pzaIjNQDXxuOrooEKKT1eTWqfugvOMX4mrPPzFfTGIGEx5qlPWRjE3wzX01oaKJXHjsVGtd
YH2NQFvO7lFs4TGMixMGcSrdcHPwyFeOfgSmC8iIg2IbV6VDEwjRZymcXq/nbKAD4NsHxtStq52I
qUsc7K5ISPrGP/9XUZHb95beqMtvtqZT2FPkbS3q0NldaFNLei1YmjXEiNkobn6Y6Bt6hzbFsff7
ejp7YIk5tgzbxJ2TZbFef1KakozW2mWF0Ye+eApW/l+5e4zjub2LXocLj/xTcA87vrGs9o9sy/jg
240xlRMe8rfVi46d1TSThhab/z8zi4jqAWJQNpeoz1l2d+59mbN4iTwwDgD83qa739HIfR9z3hcd
gIeyMw7DG/5BBaho5mAAuJHaFju113ThTSMC/nbX+VqK9135h+pRWBqCLbCaUdmvkxIP+A5DOF+s
g95vlQYd0rgnUgTCm5wlB9LK4BijRSvKCIbW6mM9NjmvTQimF3fBpvQBLyLtLiGqYwoF3rqGLW5Q
lnVZOX4EM1gumHyBrya9XXwo/Bhp6g01+Uu4QEtdcM3JBHtE6NT5VuqDWo8zhP0OGyYOa2qj/35t
q9XWL34XkdIIjXSAkYUCk8SRtOYGVZqsC91YurtbdM3brc4D3riiBqPQQ5WtP9CHFcTIJDXLfeVx
1iB5gxR6u0h1c+EvXk2mjTaMT0YcX1/I/mE9X0OlPCbdSyLaD8I3H3kUaRfgTjS8UFk2NqZ420/1
p0f/gT4U+jLcdCqqdwWfrh3Aqz5iRitMG3Gz2e0z53byls1MDS2GUDaqjLTDDwEV9wuB9J7Khonc
7kKGhkQcMNaT/KlVIyq2y9gkUyCCUPB6AmpaS+bepm+yLy2mjBg2wn4Hi+p8iMX+WTZCyAjdE+4/
D7alVVYH+Z7yvnM/htmPIsKftEDE1DWSNt9H3FtZmya/lY7/w5hYW1Eky+h5aYDzV2uB+zdQLzrY
bRLum5ycsj6DiqoOhs88JvC0rgPrdRMGWZbHrgkNE7e14Uyn+5Aq5I50F1jKOCDUeE03C6Su7SNA
MLKML1SFdDorfWtVoMK6PuWGK08tLdRxQJZrKAUjiZ7bojrPKmyVwuNSk4vywOmTPlLyEAU22Hqf
FFVvcTTKrm3L8FZut8CkbGpOj1NLmfEGTwohHzvC+TIE0lNk/BTTD2EuimTzEymXbNCadF/lR+sd
35Vlw8Lz/Qivew9bZmlXM+eJ0ngVMm+WYnv0p/Jeh1Qh2MP1DXuwTfxX3tbrPFZpYlKy/ENAQMTU
zwErIeeLNotjkTdRk7bGe0biz/V8HOuc7wvSoIFYaI2KLMhZp31SnlCpNgu/78ttYrFc+Fps43GZ
gMO2r1pZDjzXPXN8HFlVPVBUQHupzZCQrDwv/fmoCWngeI7gYf0SrpyqFhTJXCH+J1UPSdDsewby
89yDWrlcmIWli8utiCB6r9d2qsMhbxa+/XeBUVh2qSRdMGtVloXWpsVheSEp+X0qL6YEOE7d1BtH
vEpO2ds94YcvoYr8Kg0vwjm6GisnYsXIDDhRDn5W+Fv4sy7jcJk1DtU/DGRWoV7GHYi26Zx/0ltB
L+RG7XbAiijBOzCJKTjvx92k26rEcrjc7hCiXopLkN6HKa/HBrbOC6vbIcxzj0/bRwDep7/CmeRz
YdqBF4oxmj25DJhaqv1asD2kbCAoiiTeKFc1vk6em8Jus8G5z+EvZkgb1s0FksvCOsdG6PDreGkV
wVGcNXJsF24K9SLIYZlGSyUbXjaywzloiehSlDgDam1uff/ewNN8W/3wTfjO1mZMDDR17uPIUA+/
/yDXw92Ot5APzWVbqbKss/2wleczecELOdMswu0LSKKuLKbA6SnvM894qh2gqh3MK8304UAgajQv
X3DVsingCNnOtBUm/JKCeZGXiNfHqHbOPjEqcECLSAyjn4/5d5EeQYag+e8HjRVzSwZisQ49ri3y
dGcI/EV9/KB3RCGLQgvpcpXjWdCV/3E87exIDpEt4XGH4/T/lNLaOXUp+wLl1oBSgs2s63JrLOl5
8fbUaFvPrS9R3nR3gT7BlC+zxSWWEdw5Kbc5Y5MoCGtPNd/uhqP9/2up0H3QqsleGc74V/V+yxKQ
5t1T45IPddr4ppnbfW/tY9N64jey3WkOlf9uCwAGoJcIvITNYmIDaXERt0b0kQwH1Y95TM0Gbek1
53fct//sdL1MA7qz3vkU20c7AFuwJhZe4X1va/eeK5qF+t4m36RtGumfq/TDL6bN7vMmly9qr7JC
3SJ49Yotua6uIvUDmnp8em24fx2Qg2cgFo3zV4ceZqMfKrT7OpO3bY3E2r88CjX+jKcNALRlGLRo
ZcK/Oe7/VzPeAPBh/nGqR0n59dV82x7ejpzrIAJqgAZ+UrggP50HQYlC1GCWt2U04V3gA4lPq4Zl
moI1S2tKSaLDYRQU3yS+bGz+iUZFZu0jclvhI9fn447MNm/cUENsK2LbLqhSLIYSlKthNa1AcRGk
YcMetlx5TM2KouOqs/0HqJRiVZcqaddzhg16PmuFKNSwqgOE7g0l7Z2DapcQ98Q194mC8IAQ8q4e
xBfUnvq4NRTDyiOXeUPdhY7WrtZhM4XKJPqURqlEUWstBu5QkYhKoqZlvaC62mMUzzA9UCXWE1FJ
j53TY1VV0mFmOE2Q3Q4R2Cz+3tXbVu1+YeFlJiwCvJxqOgPX8t3LOuAeeVk6e1bMIdoTcC1p4myJ
JJVFrkyvd0SLyhzlqD1hUaHE72w3Z1f1nZYlMEn8dw3E98P8TuaNhYTvbROCw6XC8HZ/t1HTza4s
mMDjS/YCbOrmh2iCGvja0aZ5AyBc6uhHeAn3hHmjVyBFYEsu8sLhdQfGax9cNNtZLgzt5VAY4M/t
zwMvT3dblb1/43ZIZT0LD5I4fkbDTCY6lgYjgkdYuExU/f+S9b8pAIty1sqbRA8I0R5jsYOEWqrh
aSm9B1LNQxPIV7c1EhZsNDrnnhucszupqaS6/lOX6nbSz+Qd4whFtfTOa+mBCojdMGoo8FJhXUlB
rOXuTpojCJZu4wKXgo7N2qINWWLRhBDBCPAZ7SV5xTfuvgOdnKYhrsQ0K9xJlKbR8qkAICqNIdX8
5VE/FX83wEdPAlrEAE+q1zYKq4iOzffFgYHmsiK33aZztCGjLH4M8PcguPntD4KunbhCeFrBTfBZ
2o4D5ozv3W8SjM6ZAxx6GUXDStiBDx35Z+yJGbd2Ajr7IuYQQmimLgvRkSPw52nk9QklkzleBkfL
0UEcC8S/ylq+asrZdxY2jETOM85w5B3iqbQTNtl6wjFycdTkpENu+dWieNfLALMxZiInc6k81tLN
jroK7bEOiAt+6kn385YHizSKEypEFj71/f3n7Lo64LZUHfha9RBsTa/P6Gq9ecQjugtJtytvIjpE
JnhMQnyCq9DWWyT96BWbxGfbtmos+qRILP3Ijp/LxVKYsdajIverCh6PD+i7cEfgw7KXeNjomAkO
j7w/FcncsgyeDWTbnKH7kDxWXqcDez1Pmk1rcJ9Di2IwZ0Fw80UZipaEs/Yv3Jwy6CUwn86cQHzs
T1tvDcraYt/0lXh1dUTXE11gueIdZvAomO8ZIz8JBeqvUxP1ytTiGX+JCDB/yAGQb3PsS3XWzW3g
wHvrGSID+X7JYcYFSU5TJ7mzqjfrcoWFgnNesmVUIWlYGe+P7cDeeXrAOY8DcVJCTeY1S4Brxtsx
9SCUDjovxItFdaTN5fUaj4xli20lMutBlRchczIBjeA6p0NOos4Gg0vTuRc2WpQiOX7oy2Zq/n49
P5uT0q5h8Dzse5DPZdctoeI0XClwG4pEz47rh7OSE8cFdD2EsxdZJuh8SGTxd9qIKR1oL4bSEChZ
sknz/HpgudjiTgmddKPeH+5RuLAC9LwSFuRI+RlZOFpGHJ8xTHyOrNBnbKsw59UB+uH3dUkgYI8i
ExECkQLm7sN01reCKMjTWPa5MmS+jfZ+eM5zvXN75V8hWYu8is5mXkINaVuCxxKoVb7c9Ei7uIUR
y7nL7eKzW6k6XfOqW6MgRQzN93vtLobHxUwmHsD+Q1ebPDu2ILTkvDTuj1cYNaGLZ3c9LLC9Lop0
o6mWEHM4VcG4kafUL7VVvRuNZQiW2lTqUF24+acJB3H8ebZpsmSDa5NXhOxUPHwo+JdLQtD//o8W
5XRc8LDSukRCStDHj/XcnY8GQ9uBPjLdvFEbLpBBIMXKyrIgkFHU6FWm7gYDHdBrTzeZHNlvR6My
Oszrlp4AqfCZoE4zvNvpak5LhmxkPq1tBfeO16O8xKDFfJSEQtA/gipwMlsMRh+hjhof71ykZmjl
6Riuaf1RhES3XNyPbn/7gu2HFOP+m3lU6/PKqtz1Zkt6UIqUKUNg7iea3RZD7AEArVoLswgSxt9i
mgUuj53j9CEI5KUJLhQlRZ8UXBmaTxIawh7EdvT+ESg8luaL65KQFZQu8M4tSm8rIlgYMGcC8Ty+
7S89xBntrFFMTWR54itgryI6FjA8UzTvDBmJv6Zv/uWKS7EmHzOvcKC4/SjqFse5YE2Qa8ZUWahk
Ix6WYrtLPXqvwJPOI34FMeX4nCfgRZcHaN68ThXmJrEpPhcLX90o6YbkWy21lCrRKvWUpZtdShEt
/s3JnMExfPEx69IAihFKWHHE6WiT16PJoqfhx6ntssZIqttxnQLdmgPbyat2jHujfBP6Y060t8Pv
XlCTJ1KBO1061qXj/rAdYT+cppUDaY+u9weKYGR+ORyN3BXpRl2NTBc7QQtqTsb/5PcSS1NpaWyW
pEaRtOpmltkDaL9NbhSrHMO6pbJuiS5Zxa7nvZi1c/BEDHl39X/KlDR3Rr2Jzwo5aTSEXZU6BFgZ
X3LeJldXY2JT7p4qNDHugB4XvOIFLUxSoObIPQnBYwyPv0/nwyoO7zkHL4sZSyYz/FyXYEgs1bnZ
/VwzmPynE+7dQAy994Q31zK4YXrlKtmS8JuofmUe5hxweIEuGdLLDgxvtUFRKO0vHe66SuUq/MBx
06X+CoyKgePoHiZxs7mbUhaIbt5rwqHNbU//9B65WLdRlBCaPLfFUAtEZjbLhIjXEhtbknQJXmaj
qwYnMdAOyLp2r/0B801HQtgQ0La/LSaJ/wohkjR/We+JG6q7jdlEUmhM2AmoPWZ/1OyXw2eC9mgl
AekukCvAybnq+pp8X8y7od5xPHs06cgUg8K7fbAg/yURQVh/q/OXp5rIEJIzYa5vLuXKnYEklu0r
hnDQCX2ktJ+EcSWaDFCuGQsbQjKQAPPOs1za509fJ9O+SwIftNDrO0+b9ySlFA/qbdvA3h5gx3lW
qDqrKJvQrhL8kruh0L3OxGG/XRFAMcLrRWmng2B1I+IJqNZSpS9e9YbhCh/Wm8zDvICJSZ8sjPib
t+kfrVLZkLe0TwluljZ4JfKp+YHwADO55spMtW4HdZkJ4mA8PEEFC5gFrzwScixiM0P5oCA/lEjR
V/lV1eeVCb1OZEhI0+mEuiS/IIQRCtP2NooWxUvka6XrLgLBomZ9trEILpGht8vNmD8dKLDR1gTn
KAeVCO46DZ4p4bxAwXP1ceOjV4Wg/j9n320cuW+zIs3XPI5A1r+hs78pov1xhY5jm9lODWblSzQP
F4XXJUTCYxrY9fbpb45+WLpH1Ta9uZU6xf7pfR5vNiHqWq+yf8Q+VtRfkWAJccLx3/1anN8aGMQD
1FuhIKZaLed9KhZiUvTVPrAuBF+zNaOkyb21pScVgaHdUX+3H/k/amBY/VMEfYClJTMgnvArzsSQ
+XxtAETtEvpQDtdOKU8RD79WL4tPbma8bfnOui7dmABgSpuSVEf3udsSiG0f0nLHFFajEbK2ForR
eTipM9WRTHXCG8mXsSWgvolB9rz6oXp+mWrXPO583Oh+vzRLFqRVWNeRPdR34DlWhfK79JJl1kb6
y3I93gihL73/eAa9FPrMNV+x83aMyDMfLYXi+7z+X3oKVu4TeOcLgKS7lwsOv12V1cSX/tT2Igpx
lPwJEcq0+i6lNaMmqTTRIu/yEOXXiv/AMdWVNSKwGZZnvt6jsxovHW8lFgneKHcR8kn/FWqF6IYO
rfBxHFWYUdFollxiS3ugnFfOtwBezlRTh/uqwGibqb7ba9fGi5NgTRWm8drBositv8OHMGI6Wu7i
6qqzdQZqOmMuQr2pnC0MAWHYTbdPQXAUIehS4baAaCiIwSXSdBk/cVx1EkJXFEMkWwZAFvIVg0JX
gpn/ytXh5aoKdN/wI1YlP62fPVCDBvwT73l/ihJ//nqfJc4tqNi/LN8mHlT1ROkgOKvGxVoMfm4d
aW30esBts9D1HAvpdA8y1SObb3tRYkhq8xk+Q1zNuRZO8lp0U7+sp6yKzatCrojR/6KMIOEfTk0A
5ZHTQRs7f+YV8UURXTLb65L0a0xeTQV4LU9PXI/KSgLCyyZpXugeoUrVH4b35T67Kk4uvnYBh404
uN8Mmdlta9J3BjqW2Q5wg65pn61i3NJZBJJ10XF6wGuWduuXcenNnFoxq9RyGAtR+Dl10CvRA2mi
Ezd98Pwm9ufiLOIHfTEIyJ9wI6w9efj0Xdmegit/uJUR4BNJQbzjsYFRr8L7Fi5gMiInov96SuGc
Y0Vr1Tao8+HkaZksSmR0TX2ALekIuiGKacqCmNjdax4eQ1tZTCEYq8h1Ra2zu8ZmxT/RUACCJD1V
YrFTR2vNBbn03aJNaifjR4dsUGvCQvZ9j1dz0wZ0WIIJhOQU6J9QqAR9czmQ5B8vKVdWLkdW9aNp
3i36TZ7/93akVTlInQwZDSnUsDSvoMDIfm9E5Nb1W3iCKj4rGMqXYrp4Q12RxW8bURjxc+0clA2N
wz2aaNm6abpqe4h46WHC2bazaD4TFz79r2OvhD46snV/iTYLuiwkAsw2qgQiyDPa/U3xOcNDmoNe
T51Wc4JevbuBZxG59Y4tt27mczeYULCnLnh291cO5cv7DhJlB3pUIGw+UY8Coetd+92+jbDd+BYD
p8tU3irFGtOqu19VD8N6tvpe2LSRKgd9l7lfo/wJwEu8xM8LkGyQmoVN7+yyrhW4RpKf7rmpnAIa
tpbTzsQozMWWS5O32jrqBu/AQJtWUoFt0GwiaOY4uYoA441kDQVMykLdt1B/iTJtPnnW31dLYp9a
s1UlIZxpgecbrC0c2V8tHXUKjg/UfpZXetSOuPIvEU5MIMGvuZY64r1JTwK3sWZVTQa0ttlS1pgU
ypF7Taf1vSUQIZa0eAtQqyhu/ru40VaPq0ws3vKt7HJkZaNdWonDMShk7pUIT7IQ+r/Pwue9N3/n
xxDlRFmazQWrj3F+0kV2Z4rJaW+5ud/lSbwoy8m6ty+y524mlyhfRVc/gxXpMgyV1f2cLqrwQEPz
X2KnPKQ6wJuxZ4G7U/tpHr6nEkgYEyVHRi3L2IWSx8MZNe2mAt6sd0FVA+AKZ+T9D41lOVNDSatF
/5jYxbyDItKN9MJkCBywKO6wYJT3DhnMS6acPq0w8pl/axaYvpsvDqLdud8lzlq00gPn6gFQoZ/t
84thXlGzYxOC5UG9arzwywxEAs4wWIdy5cTRvq8NegtI0hM7ClTHZnqmwou1LTVSWVUgvkTVIbam
5zPuKq4JfgwW03ogk5T+lwbpzOMUcvKREwfcv5iAjMTwJK/KWNsHWluYYf6T5EGN5tWtRXQF9H6Y
IVkuvU+luu/d125zbTyDGI3e5JukhNgUX1G+aJaeoc0BVa8+6sxADxBhQOCfenJN8GtNWGXTmlrt
F41PVB+hUMq6YwGTkU5gff5Y4jaB4YfnGgkK71wgiFrrMiRTIycz1Mg9yGfj9sIxDb+2MJFX/XTV
zHUTGQHWfpx/vw9jto9btXHfQKO2uh/MMBEJKYNL6TiJoxYMw9NbmWAsWp9J8mHwBFnUg93YBR1u
f6/OLUZLznDZ98nheEXRsttZhihNBYmceFQ4jE6voGWxHGe0nh1t5qodSPhH4xGjWJG/mk0gbaL5
SMVwps5M/cCHiyNjt0JLHImRq/FK7pMrrBsOTXpFQCXs91FCiOCNtKiNGCrmIoLrXuDzwoZmM/Dg
OVa1dFLsbLb74TVNq+ljKRdz3ahcYvNXUNEhwHEGx+8Ec8712/ggJFXs8GTzD0M4HhfwKhs/Ogwl
zriDHSOYPxZCr+MiD2bIvZ2VONzPyKPfyICKC+xGjZNShyMqUTPyAozS6/U2YY5dIE6ujqiJzNrg
Xeo6aO8gjklQTc4Ny4ZqaQf3Uj4KjaYMdAVkI1+SsCKH7A1JSB2TBrFFn7nsdtAuazvu7+veUj2k
vlDE9Cdh+NptbNBma7ixvhWXUvQhEVP824MxBYWbQn2QqGzlX5XwQfkDUvc6HiQw5QzVYJpd7L3E
mkK7djVRCLr8GZKMUBeWEMre6+GO3vC3utTomnwpYLNrv5yDwB/abLP9lrMbFFSxS4tICwO+aWoN
DjfC9kpjCSXaBHovQboBw3KMe8SgBGQDrt1zokEZ/EjB0qD3quhv7dWUit0hHPDoksbzYCIYKvur
NsXPglgoNxn+M978xwX5CrwYnoAHqUf6uMijovkuFHsq3axWpSn+XAgqnwmLsT+H2rp4JWexlB+4
9KiVnKmSGZXG84oqVoSiwq0zYbmwioGmfNY0ZAyzajc6KYLfkxyZUJfX2mGrxc5WcdO2wDWtpaqP
i7RrTD8jOufjM1OgRiKaPD8dSfvEhg9OMigii/Zg7BrutbOKEtsWVFpINh3jvdMOX5HOILjaExOg
xNGVD6RBMrbzBRVQVjxbszcMnJ3fT1BQkdOkOEzzUi2M/r9ARDve3bnd2JgriASb5nay94k5lzRm
un2rVT0ywbfv7cVOd+6C/u/W8FZWDGUrjp609xh75p5X/Vi/6Huv1IDH7QhI2rizwiz7kPXaEEEZ
6Q/GwWo8oWJXpsqiZWqkKNvgMmOUfwvh/T0z3mLV5gPTvaqK7OC6l9AvD4aNlqlAWtp/5xRK5Ref
GYZBFVyPQFbUy3BL+jAhDA5pCfyV3gky/cMXDhoxYFNj9FXvlCNDVKZvt/E/FlVf8At/neZpGEN+
F6VPcDH0Gf+AL2PNkGuPc927txs8naPLQJMW8p9s8LQYPJ/6r4b13VPfgQf2QnAyQfgIrRYs7Mah
5H1G2FaJE/H47fokw8Wy1LhmgMWn+B1tzKRZGG2IMy9r33hD43Txi9FH/X4Z9oIRAmjODxpJ2xFU
A46MGAg87Ty3/O4ws/qccUPhP6pNU4SUsMo2tF/WhDf6EX1TilhB4Fk20uf7U4mEIjmUCmBPY769
iN4DTtx7AfpXu3ZP/Z0Lsy92E15xXNG0jWkJldgJej2iHH6bpstckIhJQsARC6DUCT8IeXWk+MTs
utHUTNJKC6xvDq2ItS37j2yQeVcvYJEye9KQcHCWffYRhQbmEjHngkGY/re04dsiAzDDdOqa4//k
O55Vob7AmOeUuPgNa/1xWBuwBy45dKPeY6J1PzxodMxcu7miBzw6tRpEnYF5S0EzYAKKEMBRB3qc
+I0EP3YwE3ZzbLltxrdZboz0hI5WlXm6Ch1A1KwEFeK3QvJSgdoLikDfHh0aGC7Cun0tWsSBQpLk
KQpp+lP9L2mwnXMsHcu7uyvYwYybYMhtS+ZRxYPsvO8OoCzncUSxBTIt2v9WG+l8v4ZMQLSWPN/l
uQh5yeXaTeiszsx6DKTKnG34bOV8yGGMDD8VScdt3YQ1yhjKXeym2fXI+l5vBopffLCGd0QkaotD
pE9suGm5ej/iNSxGLBJezcCHJhBR+rteVixnATq7CuZ3TqnBxOIafDoC749/Oces93UPoa0vK03/
nsi/uEek54WAVMyeKHN0fLD9J3NIvFdcL+Z2fBbChTO96eSkIbRu803VwDFdHQqGhnAiYnW1TuiY
4uJKpKSdaxzE+1mDaUsOLCmq6pWe0k2dFf+4srT3lvF+iQfLziHySuj9O9B3ElJgQBFRo95J/Vfm
Hke0A2IUI2WOdZFcijSlfI2599Yzj4+Jzj71a7+9was5TJJ0qeaF0YG9xBHUBCJwyu4VI0iJQjko
XEqNgFQgnCD8JC6zDxernW1iCfJKT4bmcfJMJBrXWZaD6/wY9pDuQZVygmXNAtyfr83dYihE2zGg
P85kVwV0C+Xty4g+HPqfJSmXdtgl7Qv9cxXi1NjiAmtpsx0l23OPUO+EUrcRjYNEHnrVZYC1IlaV
nOCd3hCUrVbv4ibapvvcusLSG56KFPwfWyUE5VKae0NmWVWXLf//RofCrkLeumJGGArk9lPmiC6S
DE/3sSbSMk77Td+LTQEXvGm8bOw/YHrVRB02xFdMkH5SDZmVCtFrXSWwo5kcp+kt0KFNXrg8NpMt
t+iVvNZp/rfr02Uwcr6i6uc+kPRxp2ZhvCyAjrIOhoXAjpxCatcnF7czmFAgLdlTtdHapOyMFPEp
rUozJMkIIP+FBa/eNVF1Mt/f7egEqJ/FOopLylX+JHz5JttUqSQzmUOoXvMbN9h74zEp0dEu7rPA
4CEet4L6f/lMVhxv3JD1O9+K1lpTLL3bzGYnWlhMpXspxHOIs7AenbysHoFUBM5pXUGikFp/awW4
+CYaXOimog501cKz3z+ehHlB6widZBkqDBsrbV8aNy2xhP1tGymhvs6/CJ+/Q8x/XVzMa1nJjwuh
1Vpn2nEuJhNOFDOjooMXi+pqi4Ebxp+dWOZEyQt85OPdn5konPstrn+aqXLj9QgDNbsclpjcmfG2
YJ12QT4mh1iGR8s77N2UzotOjnGyN2rCBFZblcnCNpKUf0hdiRk0luV7qR/FnoEbjbbbH1B9iUm6
jkAx/Xb71pUJ9+TNSGV1DLRjq1UahuLG6adEPj941A1uubPGlpiupfcGamsr/A3p8D54kmG7hyTq
/GfW4wEOqy3Mn2uavVvqwZ0aIO+Fhpna1cn2vP+zCjq4qAT9Tz08K1ec2R6DukLIwZIq5HQHiAV4
iR2xPV94uqAeCxFrCGCk+IaGK+9Is0FN1j4knkEmRAMXMxcJKIXdRrWMcDAX5y7FcBIShrIi02mP
DF4k6GoS9RgV0edGlrePKsXuuYQygN1b2a65Ffug6BTYnRJmpWR8pAkGRS3ruOp8/Y/LGwd1aFhZ
D1cfLHYIzTarnhXzDCMRzcyzn+FVFlg2IiUfQ8lC6Q6kUho8Ed/SCYCeI5KvJzArZXbIDhg6jucR
h20PUYP37BF1L0dpKlvJOxose6MYM2OaU5paxyp4AFqWJRFX6gLcv1bs3CWIJIFk7HQL2HWduQt5
QE9mqpY9eJbwD2N5UH2xYPvRJvmkAsVAkCwZgjf5FusQKcHlFg4n4B4oTW1IDrk0hJF4fhFCMhbt
27iM0L+hSOyW9elEJlXEL8s5teY4Khbx67IXtA0S3fwq+NbofrKjfLOBU8un8mqNWbsAyJECffVy
cecbyCyo8r1a8Om5EPDtDQYYRRljqtxijgh2eo0JWbzSneXT6wlhvg/skIYBlk0r40H2Z+WuuWaJ
ByAyuHsTPTm8O9kGCnxc3xQsk4dV15KAPSnZAKKz86jkedmRsmpmViSb4OoGOLgHRsW7FE3V66DB
AyiMQ3weybocrexP5pzgupPsnqAQWZ30sHZ9Ci/6vYCnJo9WW5ipQ6B/hNTaCxHj6xmOjt38jY8D
m6ZDdAYidzd8gh88GVT8MBY3jLN5aFMGyyDcO1U+OaL0xPaarTa5Nw/236dsF2ycGMps+nQi8hgN
HyHLrww8+8V68Nk62NNxk+fIqMSAI9qeyTaxlSW0tzTS0bq7dJMK7oA1f+ZPLlX3zEu+zwgTvV0M
8mFS5ZqdzBOOhsg5/a/yxkvyCHAJQKx7r0ePbgUbp5zec0Nto0kLY2+ViMMTiaS1Xb1qn6VvxWVq
4d0/CBfXgj4MxoH8yADU+5rGgiJC9u38uruq+MAQq/DljbEXlOB2vmvaT3WUW7rV3xOlYKV2elIw
6NgG/Z3O+9IqI+2V7y5Gdi5c//fSWw3YHc9/NtQnYGNygcE1teXxJ+zHbeLpMaxwC2zvfQxHz8PM
VZEQOdw/3WS5WWY3/AgYH5J0Ji/pifUywuCfvroX0YSDVa340d3FBy+O22WBsueDiV8JjojezAOB
I8w44eYIE42gGByo6r0EXbNY1egSN6vx2LVK5RQY3MyzwE3kGljaTLD5iCdW2EgrJNVgO+TSKaZr
/BBbC4F9jL9kesWcABfbfNIIhOG9O9SGMtN3UxIn601mhcJqYGqDGq92PjPk1B6j0oaxUMJyr6UC
tsUZ1x9HI746Lf81gWCkc67nisCYQaWkPoXdDbbRVRWQHwWW0ODErQQXttlEpR6tidBkl6C5Mk9H
8GNw2OVb/IycjLQS+ESCpzeiIW++zHYGD4dfBAz/4bqzYQPoNM2XZWzbo/Gbc2NRJUfX159mZHOg
q4fimaWeC4sRWo8XefmmdHN2+pQzUHRMeputYEC72xzsr/Dx4nRQ0toGpvE2OVAraguQEKxcTbkp
vZmdDjOb8pI6AMUUrWf6PrnXQKSS1Tj3kTK+woWhEZSpwCD5DKIOZow+n2kl3tpjz2LTtOmAEb5S
UFqJJflw2B/RiWiwEnLyqg1ryA0Lnm4gd1m8jA2I39m5sDtWx9Rfs8x7FZtidVsMIUtcRvr9aFgU
hCfhNEJ878FPeyGaAVcf0Rl9ggPp55wR3slkeJqydpriiHMlfBnpdieXY14XtJewAMNeUQrjyWzx
nuV+iwoHRRQTm9OIYoPs/1EV63BVvv5Zx+/rnww8fSgB+Xm9GaxT+14mia3ycfZE3lXrFoCPoWIn
ncBEWCAMQPT2vYt/kKrQZ/2otCxUrijmWKBw+ZuKSQdB6AvSERy7ODEBrChKCTZ8FVYRXYv2D11y
xqqOtPjmadbzjWE2ah9XbuRZn3W3hcrko5jbzAwLdTbN62Qf8DLXr8FT6sDRXwTXHiHVJoBVIXD7
X+jtZd1hfzs2Ym/brndbW44bJ+ORFrh4wt35suIVF2B6HdEUtJjX5bFygR69Oy0GqGbwSxwcpz4E
bFyawiG5C7S/AFRpnPfCD6njQaaKkZQ0sHexL9t3sz33hDzwTV7xkHnwFfZuoYGANDYpC+3GE0C9
APyF/ZhB0uPF9dwn1VdoMFO6y2XcR3z5/U4C6X0qGHuyUepgYxmgSaIEcF3q+YEcqHcie6SQJVml
T1dR2oDArVHXCY0J6BzqHJUoQW9eCPt7aGGT7rVgAFlctSNzD1aBSVxAQXRQ9zMennK5Smhgl+7z
ek87pibAugXcJyd9aem61oyNlaZxcBKxbrzqgnVwpRoxJsaeLFX1Tqx1nP+Odxe5LxMVE6ixR4UR
M3su5HwlcuN1gu8dEBtlNZ5h5+XYn0bcgf7J8UiZ3FCa46mcwu901j75mMYEXrB2zhp7ZiX3gGOk
Pq2g8NOXztwF+/5gpT9VcH7hasrN9RHoSVJMIvqynX45ksTR1emnl/HP+RugAzq6hTe2w7zuJ6V7
LENBycMImPCYIhzh25VCvZFgwmdSLu3VjIi6NO69FkXQS7kXxuJ374K62WpgVo9lb5mQzr9HQ5UN
9UTDdqp2dyqpsfQyRIqLXbEdlbscttnf+snVf3PGfk7vpIviKfec1zoreuyyRjYOeMB+qFP7ibzz
1IE2xdbnxopdOtpa8y3sUefVm8lEfhFnjlAyFUBdNqBj+s8QVVOHJ6LpVWjpSvFCzLNe3l0oLSCz
TjqZ9sTumz4r7mmYcGnwFokT0MSrqD5TwHrM0QHSSN1hgYZ+REKx2NCBDtdpWmxP4V73x/X6NBs4
ovha3L5AXLy4FfW1inBdyFrkaDeKU0mQ94PlY0kBuNhiIUwhrA1bRHF8MA976EYF6Jj+jKlWKo0y
E3CBZg4rFZq8cZjj/Jea88Un/gl4HGqA+AsE8o6pC4jSYUG2OsRU/v7QSSfDirfXD6RJuGoOXo0v
d1QRpsdpTwscYqixO4+fwoXEU+KBBopixFcoWJxO0ibKyc4XnAZJKIQ6Wn9bkojuHhvyf7qNu8ce
Omyrk/uqLKYbFbwB7kUvZ/3Wi/CwOBnu5s0FENW0Q099qEaD5TpbkuNd00lv433FYj08jmdW1HKj
LbT9y6Wedcf5WT5f9kNcnEqntPYM+DVO2NfKk3vFXcy8fJptJybiNyVNgqcZ/u6ANtOCqtttQ04M
1O2TfD4HPju5HPQ25nCncfVVfBLO0FWas1n4RdhelHGfRy1YbYfuVpvrw1mdANG9eFe64Pc9qC47
CsQBjYIRE5FfCBSJAZf59yaStVXovCNQ7KMApbA2fG/Hqt6u3pGXQCsvx50fo2Q45jQdwVz3He9l
kzfV/t+Oa4ycPXTAG1Qqlamp+q040qcpHkdWoYGEvdeppypIBpgBKW19ehpweXIy8fihq9D+yks5
3qudxBbSkiYbgXtYo3EzIcsNtr8qlyHPbrOUcWin9Rao8akAs6tJDMyJ+iFM27lWWqm3l/PveG18
9sMkpeeWJifmI/3hAq65gRVayROAzY7FMaxxr8eruMpYgLr03ns+raUhQdfRNzzGOjY/8o2yTqdQ
7FPlU2RnQDQQ8eWkE2RZUbTRtzxXQzCetSR/LnpEnvc4y8eDdbVnEwQjW4ufMLFn8H3y54ecRBiY
nyW75PIQ5eB6xxza34qH5fehwwWmLX9k4M20M3yMgJhiZEbVWG/Ifits/JXhb7Evw7FgeBeWvZ11
V4ZgtEo50zmpNNa7p2upERY6tlzQsVqc3SGiev+J9JwjdoqZy5hUtUMBdK0wlCW4ahPWv7vo+lXm
RuVSkgLiSRox4ExkNThYsAs89nQcR7kMWrvZHKFiISHxgM8e3jnSLlMzUdh6TYbBCrlGCwBtbf5K
WLaHWDUW/i1C404+RQ1hLwh5mweZBBGpDul5ZQj5zwyjzc/L/zwO+uNSw6obY4ATGvhcErH3wvWk
Jb3743sSvCz4Tj/Pl4b+0Xc86yLoun9/6xsCtILzfT8AHysixmdjkJecN1UFrOTJPjEhbkVaZOxF
xG+H6JFiwAa56pLPqAkqPSxdvSJKOICf8WcyeZTZKC/WM4Ryzb4xE6ox3LAQaTCfc8BS54YZo03Y
WNPwm5TiypCSZ8R9CFvRBZpJu7DxYCoFGT6tJcfrtTvnvS8LAxz06t5zeT7fj3AzXFwfC0mtLeb4
ZV5d1h9inDonNlQCM0Clef3KSk2iJcom8cl8ca9HVXpB2qHLWbqNrWFrDXZzK3J6p/R4BbGmE8pr
cEDU89Pf0T71T1aMAcdrTdMK//Peq7kgIjudcYMTw+v5Os7Rn2lrO+yL/a25sdSMuH4IJqzDZO6F
87P6l0Y6Yby/w3Cql6l4dxaDjd+91DWhqoHUtXWZCaltTllu/Sff2EnOZtOWMR4Fc7WKX5XxMFuc
t5jANgv98chfWL8vcPKqaQyGZBbYDbZZVguePN/hmrbpst17eAS4prU7viTjauExqrAcnWTeUklP
yC2BhYSAux4fnikWocCyLqTtYfJOs/dJaU+sQKC/4EQPzGf9A3mKDLAA6c7q51ocJ970vFEnjJJZ
e5oHbZpaP0ze431JUl+J/TQHXPswtX83/gUIULFaHnd3lZM/BvMViRDRUYaxMEAI2TeTutxpf94p
d+uJ08zdlznMR58gPvYQAOxduCpE0ywFbqrrcLfyGX/gOqjGGXLrtLrd3BYm5bkRqkI2fynUmG+J
TN8MhDBhyF40RiAfxaef8ugUjcB+wVu2DmkJZIrcE6kh1jX9M3xrhY50bNO7HIYJ4lfuCApSdDJk
13iiF7A4qzeZiMii7S8o93AnUiS0q6gdVfV33sjF+ukagcvizQiZ86suEwsXzHWro860GWcoff6u
wQe+/LUSfQezv3cDa0yPTURugwJcFuri6kZHw1eEXl9Q/7su95XarsiWW9PdztNNa+Seqr42PZTj
2FffvG+O6SAhEA76ilaY0Q3elIINHvuQnmpf8WxYilR6xxdhhmuy85Aud6u1bXP1zdTkNqMeFgEP
uo2vskAqbdCXFOz1I/24oU7eLJILk2oNY24eUuttUPvtB4ASoiNTLpeqg56zTiawVxzrNQU02wye
qgu59B0d4WuureivwIow06TH1jxsiEcE079mbfLKal80X4ROhAPZ0eXwtpwsKl8marKJvi+UHdNw
2Ie/SybPnUYAwJmoPhUrHDlJbm/nwDj/ry6ywp41MQqkj7fitNk5HPHlUaNUUx0mpNmwZybueThC
gLVB5qil2JqsXFAL1DSEDn7BXH6wgGPpCWXuNgzwB2GYSKmCAOQaLKiXBYUKQS53PDl9sYRZqzzH
+qUTO//VIe2EiePolYwYZuqZTzCFXD57ZlkJb8v5JqKZx9ymscM9JcjfFrZ1HyWgNWLBof6cTkx+
JqP2FPhRKVELn3FwZkQRSb0EIN9UTN8dUXZnCkxngYnm8UqmXFNb9nGxwl7eFlpj9xNQsOhy4+lX
ae0jNNryHCIbV53rZufuENjQgQ7DPTdvzcq5bd7pMR5+/Cv5xHKYPF8O/aVoqvWdDljymnorMix3
f67q+GqYrtIgmyTDwsae3T7e8ZZXIyz9lYC1gg1VMAFri1089tkIji3OZ0HtbN8gJTqdI6g2MSjV
x4WRY+FPL+ODhtRDjcfiEQILm+yYgkDHnQqBp1ei8g16EggZm+esjOvcodVPiB7BNmpedRd29m18
5x2XyH0mtA9TUcQaYjfVX58SAXZ7BNw5I5y3lgDFLUzduVVSlSIHmTBCDdx4vl1uQZXNEMyGqUnX
k6osmKBb0s0gtSIRh1CrRKNTWGMZM5EVeAtAbUfWO8aZfo7e1XWgD35q1eZxtsPwn0DWz46Nkbsf
iZgrHyyDJ+iqV2htz+FpUgnEGdO89pscBqau8tLRa2T2zcTrp3GV1ae9F7SZbDObRuqL6XQnzK+M
oYDKpa/wDjpFiGMviuLlXArbrZPwCLjIpEoF8VTT1pB+Deh/UI6/IvuwO6GmiFPUfMJqLH0OR26K
7am9VMr+HcWnGC32BYqBMFfA/n6rl5B6q+rpF4KTiKP6LDDwrD3vCvFQRH0V1q7Zn+4tXZFeIxEj
aelXQ1P3uF3MDz9gEbpfcz78xvRWk3Xe7H7Csd/yA7NytJqLk+MtQNO2SwZ1E0i+R1Iku4HMPzU7
PTIv5oDPp3d7CovYi0M101Xr4BBwUzKMSJVjplMuUJLyWqyciwW+GK/8VMeMhjJb9qZIttmfdC0K
Rx9JqtrUSL8P4tGhtIHuC6L3qS8pAebGHV7St2rH6+KwpCVI502v2aNgWX2Zv+AaxjqXUKoyGuFC
DF70+VzhmLrG5ISOgbfvIGwEA5hZ8xKcDhssOeybD1UGCBQPX5OSRk2soRWuPt0oCo9HDmpBlNSq
Lb6X3s1wflwUG5jUEUJTvoNoXVH2F6OykyIps02LZ28Zc7t8DOmcRqyWekqlmLOJvQQwFAIMWZwn
B5tnM9Xlje9DjDYZp3xrPkPtwtxq66h8Z6hVe+DdX7uKeQBJcsgkWJ7THVmxI8GkzzwXeOQdifsJ
mRy7ODUmGcIhFiFqhEPR20ROevBl0XADqCtMtRHlyiTAy4XiLH5XTOUwSva7AfDfiUxEQJAJs7lC
9MNjh//MgZk38Refx6oNhhXFltK6JRONYLAaCX/sg9OdZnMt2Z8E4Rg4o+g04cMndT0w1qEdkvNz
BDlVHiwLbGdU0JGlEZG5YlQvHdPub6cgMsJTTke5pQUioeGdwXSiefNjvjh+e0S/kb8VVeipqPy4
YoPPYV4KIWzMegRL0zLtHwDKXu5gSu860wPCdE/DAAtFIfF/E2rUnTwWgSb+7m+JkB8oje+Db4xt
5PgzBA6HqdY45gvqR3ulVRpA12u2wwGk+pqZWhMM8CRatIZCl5s74uLXQzYaLQiv5yaENO9fpRWk
8Sz0oiBDTkroNS2SeVUAGtnN5f3EPBjUiqSIRiJGGOjFoFnPep6Wfse35jACZFc0QGYIaWMmhzo6
TuJ5/WaJz07ZL3xm3qkGJDQQ4cLOf26t+3Xw0RcwdeDd4yzsx8jHCP2/Ujrtqb9VJ6rYR1I0RXQ1
BzchKjuaEaiGTpHY2nGxfl7oMqKltWjpsfyDKAPh6WpXDSlBx3hlGqw7Jr7F+9bbIt9PBX9CnVpR
LKJc9ZtDJQbjXaVkumAwL6VcWThqmKU74jqSHYnlbDj7R3QjGwAxvLwuY6cM0wgsnQ94oPxxbqCi
/OaKvhX7QuIxsVSDAjmloLwzVPVhgJTreUUEO9B97q+fH1F3JupznCGn/cF420+dn3QjM4vSGIMe
nwVok47w2BosC/ur3LpCXjT97FvzXSOHb0oqCE9DNwLda0Zv/u+MvXFGQG69I24TiCX2e5XgpyYc
Ux4dkxOWDCjiiWAl5DHKUOSEA2xqXj487b7BacriEj43dOEZCYm43cUNY1t2qD14iAytVQlHZAiJ
2hi5SDn8EsjGHfqFds5eZEHPnt5tunu71YEjcsOdzFifroqeu3zwaludQt3HWabSTtJ8cvM+2tyD
zLZEENPgKf651qj2VUy4ZjO/R/1DEgochKQKkP8ov3DZ6eyF0L7zMAB3H1hzGKzd2vTGXrFGs2ZE
1I+MtQI7XsNA+8Mv6ae+lgMHCQ//ilOjR76SkMiYSMutj/8SFc/GnozX21vNHMpc5l5+zTdFSzb5
nF2Cxz3mKUN5tc0a81e+pMkwGJY2QgsHbH6e/r4G4m6RoaahU2ouoOTHBzsrTxDggWPdOBI3ek//
j1/LzV1cI3+YHtxCK7cE8jR1ajnPBbdeHg+1265cWCwonQ7atOdnU0CC/Qap8gFnJ/QWEUtYqqAd
jfwqTk+AdXkMHdT+NkJpGayKiRNU4GzrSqcVHDz8vYNWeo74yU014D7lSyXBA9D4u9hexKQkcV/q
cey1CPFCDNj80JcQoT9KXSfuaoQAeF+O9bBb251Zwd0fvCxuGMw7p0GT8guZ3/rNQR9tpnonowYs
RHDnEFkp/0RLWGtK4AJ0FHDO6zpVO3m6ZYH+JlLyjjptnXgAF18NkHC5JB4OMFcrKLZmtw1N180O
eCfeWjT6iWYBLmhIAhnNrvY05obA6wVAn7kXg3t1nGU0LQ0bKKXxe75qajr7pqkjRFe9CNmy0Zw4
wgchnaFz1c+ZfDU3niD3Vpp9HgGTab/b6oN7/InG89aDDjHd1D6eoBbN/9uV70YgmvY80r2PpTTf
lqnJQJXLhYKyCJVpHRUynt96rdR1+4JCYvLJ06bDGXKDjNjV819AKepKe8BsAu7yRG6PtosZUkcl
LnRdXF+crW58wXdzv6FRShYMnAjekdAA8Ga7FueO3P8OkRdKQP10JaXkI2M1FWnp12PUGtMoBOem
GRFVdODmaWf5pxo1IUoAWj51fx4UEjBJp+01+xU9VcUiy+1FpKCEQitEv/E2tlIYkmgFf9yUqKqt
1rBXsZqjkNaMjSHBjgFAyC3BzVNFNwDDDIL6DdiGUMsdJDM92U0uXqpkgu/3mXsEqiHHVNZQMGwR
z9NfnDx4COuFGyar+S1VFIhPTS5U1kNT6qTkvnlXMglcJBb1H74WJBrreN0MkRTVjQokztPDVC0G
xcLZdTNWhTJ+U3nLBbhB5XzZFQ1ZoHlm2QAiXwIcO9TNMczivwTUZ692xLN0zTbw8L8lhfvP3GmX
sgxl83fLsFojcIFQQ8UTLozN3MmMKh8LNkmxaPt118ZOQjxUAS7eLvjSTsD9hYCYOiXc4EbtJQbA
LAGaYaUfrKqkYaptN2+BLWYhcvmFf14upOBnJGUGEiyE4f9d2768dRqTAmVlILUqWhp5l72h1j/i
TneeNLhYlWrGESk9N+8EnZpc/E5ljyo8deQPeUkFRXOKhdz16obS3kcIfjyZogoZc4W5rWeNQutm
6O5eGQPLq/B2JitNgMYgM8xirfxEyGBCU8z3VGqR/mD3e+VI+ij4ShF2qXJxyEvc9awZD363vge5
aGGUIXOW/6yn1yAO3uFjw8lD9iScM1l++Sdcc2aUQ+Yeir2NIdZbc8tbMb1AsgmUso5/qP8IYoXl
pRKCoe/0Uvvm1YkgHJ2EIHG9jeEtNYgL1WpmOaSmzKqwasZll3F7IGSqdp7/4eKmd/M+jP45t6op
pfjBzAkObWer26dJP8gXp2MxV59kWsm9mJ/DbvNPVHDVi6tN8N+836fMZ44yOFmeJtEcgJ+eZPZn
LHUY+ZZQJ54CoHDD2i4OaVyU1LahPGfEpSyLqHz2mfNvdtjvRlSYA87D+WF3lKvKETUTJcBzgaAt
tcT3uvIqC1zASfmt6W/amYcHjSXDw2iJE2Ma47aTjzD69gN4XVYkoERBtXzTp/AYLiS8sKhqrIzO
2dMLtt2qjCyPFq4VTdxBFN2cMiIPbopOBnK51q1UVSzrn6/6I+RlsqrL+LcPExSzjSdoTfYaW7V6
K/tlcH+W5ZrpLf27VpxyQc2zuEhU8DsCh96/nHdZgU9NT0+Y9O0TKfFcFGdgjtQ+J+e+4FAqnDQB
XxF8sDi0krBS2df2/08oxmGFgdzm8II6dTKdUAxZeFUxYelVxiFtwjxtGModdp4TWPdlWHH8cwPN
TPnLZZfMzUmTdAyhK4j/ImGxeQjA/8EcoP1jtEfGFhBVAeAKnOVOaa0vw2aEBoH7HlO5Rkv9tjKE
xCNJKETiPXMoJ5UDJEftnsrCPHG7NXhVvt1lUOhGas3QvbE8B5paIZVqS18gJ0Ej/HLEJ9PgNzHN
7pjBf8kiRIS2gUEavW7YQuIqkH61RKUjFOVPSvlBf9MCtpBvjELWS2dsj+2gtJPNpxSXF5s4R/lR
I6snMiG3xpCd2Urd0vwUbrozUf9obHlvk09+ZNDpDOebOwnC7iwaQB8lTvKcDB+dqouvJIDUBXih
+3AvR1jdNkpFm4ioGVCnkkEZeK23+WKhphaSBYUlZ1uekogY83HkyurLzQYhpH8G4kZ8Z7yVeCub
S+GZD9fvgRGEop9ZMlfQhWxZ3+oCRrN2AuV28GfkrWUzxXlBsW0YAU8+cjNJzAurEynj5IgjvRU0
BTW9YtG20QdH1IPEXSjNJGYRek8fKdREEQ67nVE/zQKKbYS2/n8Co0mOAoxjqu7kkZhibhifwKWg
FWWru2MoaxzR44kyV0AxNS1gZELHTkrV0MNjC+rWF58XTtw2HukSNH5BLmGa2D31kvSrO5csX2P9
0I/n3x0RMuUEKlvoyO3+N/fa1adRRB5UL3n4sNeI5pd2/2ZA29zZtxsMYqAYf3GSTvd7rFAHL7UO
0VQUXFBnpcTHavTTS+zODuyMrdtD+Qdk02BV8F8RdWQDTiKxE1wjBObPhnix4tWEf5x6V2AJrNTl
jFT+nR2LHb+EEgNr82WqWpn4PN3WrWEmULRGxbfqzws2lu8+hDUWZ49bef0T/6nBkcik27hXHTZo
ZLj+8DvCSWeuf3N909CNBA1vEO4FLdz+pNnfsPeVb0EKACKyH9DXNxLgzH2TFvI/BVGOOQdVJ6bk
0sxkHQmcIrUfgWPU8/TupUtea5rpFQquAc/xqOCjOhvaiE40v0/wwW3kkrdS2LlDs67uxZMXJfb9
odYke8yPVHbV9RAlgrrfOAQloEXO0pZMKhpfq4urOLhlJ1PXafqQxCyAMi8IbGRDsEnMhHz50zzi
WiCm17XEkxoFpPWKeLjadfDPFb5sjGVV+79rtXwLis1xFRqChw2D8HHBzqAlyOLFglKE48tgmuEr
hW85kCYkH8UN1nUt3q5CqwDzcA5ZBLnVBIz+9WYo38GII2VRu7N+j5GPHyQvQnPFg5J4zFb2kNSX
n4nhED1XyipZKvVobJkgUPzICzxl2vaUhwBTrCu0Fm0T0LaXmP2BCR3/92jezMALzqHbrQtPG8Uo
MSx7oIz2t1yfqIP2/UU7ff3CwkUdCsKDJpp5oGMIXzSHJdCkNXeDQD8k0LJqguM/7qXCNTlQQhRy
6PBG8dKB0cc2CKZ4ef6/oKjCeeb8cxIom19UcWz0IMXDsZifVUe+u/B+2eaNyN4WLS7MpXRDDVuD
24e1Q3lFD3S53lQIUCb+H2WJpisgToBOIqfVrstpnC66b6NyJTLi1m5cCv8Xh9HZSRb0tFSm8zdG
dJc2e1Ik1eX/wXgIrcV7hkDr2B6KorgRf67EsqP8R69H4rwUF5aVKeoOgFjIRF0y/UBFSUmMJDCg
sZbAyMj2ccHicgdFPkvdHgJYCI3ksnmpNEvLWIsrgT3Tkd69mq3LsdOmfzyutpLjXkrAA+didqRR
TnCE9a4SbMHdA6gP7pfKVQSpptBCk6fIns7x6KNeFjUQOsCAiXMGoIwv8O2Q4S7iryk1tqyhNYDt
fp17sk0zwANjvyCnmQ6x9L51ou8+uVe/s+p8Li2YpVkw2u500oOv+96fylYGBx3LutuBbTy5KQyd
va508GlyqFo4jxqOCw0PYLHWcAF2i1FkGCwStTtIIH376QuSqnDNe5lfyU8NQkizos83RYlvDhD9
7ZH3ftLD2wsJBYmy+9d5U4qkUZLkPgo1QI873Pjp/WKe0Wk4QrHwJLtelNfPHnjby2nLUvVdgPvk
Yl9hHV+4BrGLXLwHyBZYttGNTQGzj6C5kzCKYbRESndb8LfHm9l6b1jQMHl5JFuwSf1FsoI6j0Ou
xQ6oNVItuqkPJv3sV+vzAWnrST7Cq+sH9pSMF+gT+TIPqIEFV/xZfRgBIZdZ8n81qWiN7noJ7G75
n9Jv8Qe8KvncMV0PP1zBq0PnkPQmwpAej0Co0oKDRFAvOsHQfL+wKXYUcpGi2fdiqxZqzxnDneup
TAkpSmw2GkFH6dU5dN11woh26DnQPc2vg+Ri4gixPfe0TCVdu7+vS7AAFq6cMTBGXQk3uROFSN/n
TavNom758KqWZkjnigr2KfDvyjcuscDoRHgs6jnRXeKWGacdqlD1sQtWphN2Wz4SNS6U1XFKL7Dn
awKcWD0fLIbb2Z0Ddl4+Vv4vbHDI95iP+DCd9uxRk575EBjM4zH71AZfa/jvNJZLaR2/KtM1eq0I
a9B4raOBoYS/foRTpKQqiP1rCupCiWrsbxR2P3KP08aohKTCYxaQYQipEa5xkgT6PhkZ1tbS3aib
9W8c8JVeOHaBSZNTUG+z114Io7Ya/BOK4ds2Yhp1eP76WM8ZAR0LRNrGWmiPc7znAM9fBcFSS9qi
O4ToLFzRQ2mnEV9714BSIedI3YjlcdvcbnkT9UT3d9XARvhKQYklrvNibvpW1xTVj4YsPtyOOIuC
Lo/nwwRveVxRL4dDS0RwSabFN3NjPw7o+Wc3j4d56YN2bqLakF+zL35AXRRKgBm6YAs4HlffvG2h
ezP1MJhMeTqi6/4Kaad+mYf8oAHq8jFNuJSBPq2YKxbI5AojtfDGgLyK6d0lU4JqsFVEaroAHIz6
5gsMUq82HDQS6aYI46D3uXj5y22PeT+02fYPTqZWXUAo4N7zoyyOuIwcFMCMRSBusLFV0Z0RPrk9
0Mc0/awLsGkfY10joiYwJMB+jwk/5tT+pM6qx5Bv5wJB/0hQwGKNOLE0wPVR7Qu95tAMiVL5pnMv
Cm6uHEyBdHbvEjdu5Y65OMoF19moYw/WaxMbBCzJEG3l+sR76fo6f4Ov/wtjEQ1IUvoHH42IZLic
za+Vg5ydfyNCl3EQk9g8tNCyGEG+zO3Czq5FyVxVyTQec19EXnbeWouEZeRauQW0Kw2Qxw+g844E
wQW50HLVnuTiyFikeCtnc4G29xRYxdKQNPs3LNAlHAI+CH1lrQ8/fxEy26jVDmBtR9jSr2BzSRwz
+COiyh1sIp2o9q0YAxEBh+uDg2yolGpQlzzcOK6J6D9dNN8AUcCwe3P1bY5JauE0/MuQtikZiAN9
QdwR0ECDeKL6NjFfi8ovyCH+ZEUqo0HSD5542Vf6eF54Aq8krGi6To70ZXM5sIRGBMMtTTICKs+S
vTyF1sHz92zhhxKYUUyxD2PAo/TJ7UIddX+E4+nEoJimWj92/+rT+h2JtNYhyYijthBd+0JuIZRA
Sl4qy9ZdDH1mP4XGWUq1uFSXDSwMhSJ5DL1wOddBq7yE6g6hrmCSQ6p9WWAUGsRQHy1g7Aj+wuOX
lB0rxzUyEgvYr+b/3Z8MseAIEksqlSre/xqOdQUvQ2t+Z/PMP74j8usvjBA9mRrEMplZ/+WB81xO
8/35p7c15s3SrHaeCmrujoUeDBgAKX8xsFbfw9vi5smdyzxmoux1W4Jr0aAHXcqfDkcpbQ4w3jSB
ejhl2HLi2GdVwf7hroUs3Yce5EIEMs4k2UAoU92OxvwWRuoTTn3Rcm5OS8OmGX7lK5IH+N8EejsX
k57woPVfsi4uad1rCYZudEecvlGGSFYGieleoCRvefuihxzlzaojjEic4Rp/hYgtiDku2iKlwKTk
ukpiqHnIn3b4Ih/4zWQY5spC3HKItC7YuPmf2yq5l+z4HBltrO8ofq2bfOzcT5yt5WCrGIocFfVe
GDYhdkums6BK9yfKyz1e+mwlPEn44soHvnT0h0THRjWrg3lpRW9xwjKhYNH5RmlTI2KmEYEW+GFE
0RpjQGc9MsMzCeaHhLzixAROLKwO3Itav1lCFKRrj+jnZDEBn174/maBv/07vc/UlgF7/jmVFt3U
D/F0BidWWH6+iQLVxx7jUt3y+sjMBOJG9uHtffJMFiKQzC3UwFBQUHGNzDsdIDFGLRgSIFJZydls
RWxoPiUn0bfwqivTRJ/tp5gicLG0ZwgiJwoZprpozz6nF7wH2Hc7Gk9tf+cAeAYmeHXWx8W6E3s5
+JJtxxhzwLpvHhBCYKHHiXsyX+sE6PwE5hNWwhkufiPzGiT6kgFQNqand25Uxwcl/l72PBLgdI0Q
GwrcoPaTc2LKctDTeO6HbRdPJEsyObOsznwDha0Um3MAAt3+CJ5Xr/4P1E83UIRc7zio0jJ2BExV
PjWA/c7WTc+s91XS+0ioRSKnuniew5ekHU0K4lyRW2qMGzAKPBsLW7NgKUHOjD75Dga256FqJ0O+
jgYHEIGMTLerq8zjXFM5IdeaqZc0pPfX4Tzzdl0evp4hwHGasFClvGog5XgEW/1xOpKFgiv2ydsy
YzyzJrqZiTumpYRMUfvUpHka8mqt/htzjB5rZAXw2rFdUUHUSGQ/Myks71/0oJr3OzKQm3rcpjLv
m8r/eFO57Cn0PAadCnUvjr1KS+As0wxBN1WRlzm8QwiscNQrIvEsmMjM1IWe2nm6I0um4E3nYdZh
9gTjrGuweTZh5TxVXD3U+fkistkCC+LK8DYr+X9c1fCQbX9bCuhyEPP8hTnqO+6rzbKIR/fL91+p
VkazfJoG0o9k7XNyUy7qrji89k7Pf0AIp3ADorOc4ijOgbIflsV2fl0ZJYoybDqUFR1vEd1Fgg9b
YfoRc5Gz6uFcHg2O905LvSITlgIZPQx0iBQ2pAQ3hH5iPfORgqNkTXMfnbIZD5JbNtJutpY8Is3v
Dx8DFsyPWrttMDcd4TLZWlQ1mPDh3+K/ELmaSFrfOJpy7zQax8OWJXxUpch5UhaL0NI0iE/n0XQ2
Wq9pFIBa2YH2JtEyWx/OFZ5qgVi2dOw02UKIxmT0qUp60TpW62JQyerV8tCUY1KFO5s29PHEIsu6
+4kEXkrx1VCjpM3PkjTTnU+0puID1Wpz+QZep8Cjjam9cxHsTB6BH55ZaC/DPOQps6zMJlRDYT0B
POsxJ0dlVERQWEMmgNs67Rw0piTPlgJxULKjYzfGhPF545tmas7a6YdU1yPQUosjrR9aJC6D6LuT
cThNtXz3qk8DNH3URuA0l+QVbFRdYPnYCEfUco+8mWYGLQfyR9hihqYxLi6skf4kQp+PRzGYWOxT
Wfui1qASta3B7WQmqJbDAxev1jD+iQeHnqs+x22Lr5HfCfGYHoa50ShTlt9ihZUTmmnqkBMGl7P5
PtuBcy8/irnmDwerrNPx/iyH4ZHmejuH8Afo+1kBzAd5WeQKfCSRgy8RNtl8qbQJJmSz2VqiuV4O
6jBXNfX4M6gccy1Lzy5a5ag3apsvz8HJKeG6OhbwdSTF424ZEQaa56XBLd1ihg6ZNpR1VPunT+Na
4D6a7rFrjmQ7PtzCFiUId77NsqISuRGsIHh2UNgzPNlrysl0wEUcxEL9DVuUxU1KCpcZzRpsBHI6
+bal31Dqz2T0cGaBCIUL4mrzHho5x0Wc3DkATTyNT1r/7umWuuLAI4EJTSMqL9RP+/OXGjT1rx2Z
QuD9EgwNDefy2WQjSqmm/TEuBBvbY9T+RKNvwKv5M30O7oUIJP3gbx0be2JzGUuqRpxqWr/nKy7R
EPumHXv4DY+mLELesQVzj05JOnbiYCVJtAlEt/Ci2w26z5oxwdmOmXeDDBeT+1UOYJDCdUNidOYa
zGoSR1ERVx7obg1it+j5RSSBQfUU8WLAnPO1Lu0AswXbBwzWMlileyBpMu/pebhtdNOqw8sEpcZ2
RH08VWuDlk4RzZHWC4+Rxn/HbjY+f6diFMf/tE+ky8slYx7J+eVgbH8FQExSMq8OinGcE4s3qGVf
iDzlAMyd9vg0lao4P+F+5EqxLa8YaC/cRBZqS7txFuVze9BjCMdq71TvA1XX+BYfKtTQv/bnPjsf
+AKN5GtbdXqyGhu+Wl+PlMXZEqjfxB9QE2EGIP4KTemoYnUiHQzD21aCZLRE9aBWT6hpTnGICyQZ
u/gR3byM1dW6lMEPsSkD+b23/ZIfEPtEmkRTpzpAL1Rf8156QLlsneS9zS+3ONeVgig3OJx/xDxj
+7jNEmMiyj11Lf+eVt99W4oA2LGOn+D7xGgmV5xETc9L2AN45DmXQmhIwsy/aeAVtM6jWqY5qEpM
bF4PvhVaupihdzsYW/r7ekkVtVVPTjgB8SPzJkA5ZefMJgUuJ2o1cDr0hrqrOTDPa1QrT+yLflFV
flPrlAUG/qrcGnhLzbX/aG86B5Xd0eFXQ8GcTxOaMgF8BKJeaH9cYn86AWXBLOg4fCDGUbBZmv9x
maiAmbibiVKSMc0llK2joVICl2CQiiFMt4pVvsEzRYJt0f1HCgwNWTAMzL9poLHj9IU8N1oW/3iH
XthqKT9VM9xWOlHNZVdtCyTI6Fpg5VvXDRkgnhIpw3LuDsU4TpyOiJ8cAxXPvyZOAW5VDUpHIuFX
oy5ZKdP4sE14MVAv6BD1hQwmeDBc402o6b+vYJmLAiZl7a8rhDaOe8FBWadcLjWoTCbUWt0KgtXN
2My5pXguuTYzbSFpeO4gbnCH2m1z5MpOAbchz1HnzfAdikFpaD8g+O3zBdF7Ep/Alj/7p5PKKygQ
qXuCanN1GRTQ2fzMEBWO2f6hbmsQ7aqOw38KxIw/i/I4l2TBfdY9QtH8CKp0WGbIO+Qq4sIGFZ6w
I+KRt3gKv6gIWZo3VVZMuHmuZ3yvYKL585E+FcYKYJLnPnzYCZ0KomovvpXa0M/jTsjXBHsNfLzc
4KYyal2Ympvmt9f8CaihCq41qnAAbw/wa2rGdIu/EZEdOrIv05unDugIXvT2VAXvY0TXuKOyWAfR
Du7CHjAszO/TUCOX2UzUMwMIXVjRJnl0WNZU71ubWfN0TT/ijGjiTkNK04QqephgKESiKOH8un1k
++Uk4lW2LUJv6NbOuGMLrzTgsAV8WCAYsnhcryDO4zh3EFj5CLkxBI/qL+hZ2bNDOto6CRvwkw2K
/EFNe1siAWxdXOBFyj2f3LiJ/zpeaz5oIIhhj+BSU6FeMJ5MJCTiVD/cJIxq7t9r+QZrfSKM5Fsc
QMrsGPMi86zMdSvZha/M359HBbFUkhfCAs5wgNEjCz32CJgsQftA6pvForAbFxs3YV+x0tAqU0iZ
Kj/m+8QqzoMO+tPU8BEd7UNaCZBEDmVq3TkFFb5DPhhFo+KSE1UrYHyFTm5p4OBxXnzT5X6N+09f
qADPAauhA5MGNraRmmIiu3f5OuYtOVpxSXLpjXLv9JVfmzdgbnyB3DkrN6fajsTkrB0KkSJyemEz
RD+n2yGTwJb1h3vO6Qjlz5VYBF2Zv7ZF9RUnSAtrcO+NiUaMy1npjxHqKJeii+Gs+LS7Cozt17js
Rwa0dFLuCIYoNIPQEKmNfNERU78oALV+wz97oHW6jAigFXt50n0D3QH5rPj/85EfUxBHuARgU7ae
2ywBaJ28g8MQ/V3zuy7gVbQzG0FtbcauW4Ob4BUHmjUvg023ykW8HcNmzosCsLEU7LZ2gnVOYcXD
cW2wyR0Sia9C0T4Fc8O9unwGcY6/eH5XK29i2zVawyzvIMgbXgm9TWABBA8w1dR3kMJS8sQyNZ4D
nlY1QtQAaud0wzNKdISxj2hFJcLMqbgZpaCgNueydZ9agGHRcR/Dmsdx6FV0epjGg+fXtHYnRk0E
h8XZRErBPk1djyKTm0W3SZQ5kmoOnLdMoFvd5kqO00OUa8WmBWShRXAMlb6c1G3VxdcAslqev7cS
mhYb9UXOH6MA17X5APDrRYSFsVQU+YmIGOS2Yy13APgZ8+51/O9vaOuHXuDg0cfFUYO48hYJedKk
2UP+JavjMRCI2qxfxWIjtIGKSYZ0z0je2DubRpgxNT/yFtBweYLm3j2UElZufik1MjhjFoc8qucs
lhg7XWp3WgVAzJSSdRhHda19lZjEH6fPv+GGWECrWQIH+VFVR4RCNlFi8HNqUOvYK+w0InTUu4QU
3kPPlv/MnVHWxHPTqfdpx9qjXfrY905d5OjdE0+rETxwa8RAw0nKFprBdwnLNN2ahdhq6Rq/5oOT
AyJBxeabHVFp0Sx16fKEQslAKDyo7JktIQFJgR8RIfQGwbmkMBwVu5wLqkcrhokmnF1A0oVwkliv
w7haJ6VAr/gILcQYdXTn7IrPGjRYif4iNpVwaAdD+2aU2JFGJ6z5myOkdGUCuOpNgj7J4h6QPSM3
pH4ZoX76uliJaZaVF9J5tmtIuDtKp2qiZGUA+AM/6ku0Yx43h+/llyh8tIr96+DC/eoIXJv1yxt9
fE1EkDXm2bDfQsLMEHi5A3xq5hW8CJ/D9dHQCjn1yqp2U2v3vYymzvR6RrNGIb/R3y0EZZJ6maJL
6YozJbT7BtCYtlVLNZQ0aijnAJen2pvfws5mKBNX+Swv6W5/sLYewiyiEr7ssx8YsBD0eeumTRl6
6yCK1VivTsy4p0Qw/SmCLEqpbZSq1B2RcbVs0QHc1tqiUnZTvUO77Mrz+BycGUT/j+NjAO4lD6LY
Tx86YENeT170ij3MqrFf+kv/xzSplWuhm35/UhQLxGCPsoXc63M0uzo88PQfrODndvJJbBpX8eC0
0xr2D1nmRW70FfkNkQqwF+CkTJ+OMFeAny19n+auLEKeL2Smg6TD9q6lNSNPo8qyJ3U4ZS5G7IUP
cYJQDDa8fz9aD4ywiRNExmsdTSGy70PlEf0kxUbZOKnDKsOWBz71U/8viLsoITybd1TuoKj/4E6G
PWS01SQX48oSnykgcizZ02R9YCznhw6/v+fYyyXRgZWUxMb6ZZ8CuLUz6MNrbl/diKBFz54kFZxD
AO8qOT2B/GVlPruq6q3S+ignEUGd1Wp/TBSSGKWKamsF4PicHn0mz7CctiBiq5t2DJZBnOtKUy3J
vxM0tbJ43d5YLkCS3oFaab/47Z0oSG+cLMX+egE+hDRAuFqu/Nk9xWzHxb7sfyiTzriaXep1U3Fd
hFV9Muoz4PjbzARaIytbTIjaQFy68SxMW1CPt6VGXQcz3RJvUFi0rHU/VeuemCEALHOARcBaMTlA
oOXhzDvUXQJwTIFbzVR8EflLlLKaJilTOs0TsbnQRT4zFzj8pPYZAZOVPiaTc/V7Jy6IbsgZLMfj
5E4noLPu/8jCyAFhWLjfumcmAW/fe0zPl3MSkLfkPLuVqAdP+e1NUhH0hd7TAK+ioYdlYoRTzrnR
jhfKYgSxbxj1Tf7Lfeq9ut71EcFq3g7kOKUOhrhpP2vpSblRGZd/gR+QKVNrgYcmybUTvPBt60GZ
r1s0BrlLYQbHnf5Jd7nxHT/cnxvXL1jqaKDfw5cChtVbDu9CiGMLBILnYdaUdwFeuqSQ0XShYW2E
Km6VXjZcEfX/Mzh/7c/8OImRj9dDU2gtGPevFjKDmWC/KbjpPTO8/QWuYPXv7IEyL7igqtvLDnu/
6Dbvkvtk01mo+k6nGrx71epr/A647IOcG6ndJ5THKSy4QSuk9HDZNYusMMQP6nAeDEhw0fUjekt+
b6nnkUHA8syvA5Bd0MGoaHCLBUdl2y0Qr918KqqSPC3qBKUe2uBpoF++FkCB9Qq+sMGzsTrVuSnK
2Juf/PuLRe15avQH1lBfhJT1bi5xeCbhre8DTebTG3m2rpuG5MFs8SMrsEo0clNkjyy3uyBCN3YG
KZff6hpM1VN7MkTyorcPAP//fwuyftOks4K2rX3Od7/5myUOLowDsF1k6t2TOW0OxUnkrXL/mxyK
EMmKZnEKI8lya1mrUE/UzyWXVZ8I6fjselnHMzQogueuMW+mO6i+SlWVmOePPCAbrkAWCbIhsGCM
86+atc/VCL7L8gcJEDG3m468TjrPPPBEbkJq8sU5y9KGkXFDDRUfxdYgO738SlGYAqksBiZt57c+
8jEYmXSdekJ7bYtAWko4mQFNchzZXuYEONGlKLNztnGAIwfWXhIrIKgH57gXteD6pZ8SFURSEAvv
URWVS/MLlCxT6QTJqLOU75b9BOMSbLrP9fd6Kjv1XOprmwivlWBBKNoFcSIp1D6NZiMWyP2YUt17
127y5Uzpza4ozYbgAHmfMjJ6zv3QhQ1hHu9vPxP09Nbsx7NzkjQ+lcHwU2nd/tUbGZBdBgzkbZ+7
xGrEqKGnCoGI737rX6vMQ7hklygr6aZMto70+vpWVvSm+wxemBji2zWyfrm2mPV6Gj+SsacM3m8Z
Oz/sNTmG4foicVa6uc16GINWo4Nb1sMYDvHxJQ0fXczRqjIdxWG9TFJ6W/zRqVVwHSotkD1n+BVe
B56PR6Lpw+KVa4YhjIORk25fAEeyW7i6O7Mjqwl3FsYE1HB3DnKA0eKrim/r31Wak+ezSVkBg/Y7
n1sgFFds332xUDF3rJcDgJfbNg9HXJpqka6phcQgIlNvkUOipxjg046yJ0X3u0Yk8DN8uvyR+UYD
e1UhcvE+N+fTbesG735jKKQyayKaYZmTOOuZILW0nP/EZux2VucL4qRwQEdJOpdHyW+o8fZVondu
ulNfLdmLwDPyqLWVhkDmArhgJN4qoHXkBOmKDQj/fILgBbwqqtkmeF+hLzq389L8zskviLqWTnOs
38lwoXViCbwvx414DxupG2P4hLgi9wXt8IMAXVxb6nWmPD/FiZXhQfYyTTLCltYIC1+IWkg0kkNW
ze38wjp5BKwLaYutCcKmMvZ/JzjcO0nlQ/ROOjeK/RHz1bERNOMYsTyrymlicxx9DX8HoKF8lySr
ASc4gc1+UCXq2YxGJ94ZYw4CXuDS6fgJegJd3P2ICjPLuRfEk0LRJvPD68AEaTtukBP2QWg8tDoU
RNA7OdbRZR5B4AF5jXi6aM0H+cyWB2D4Ljh+WktiIJJIUcz4pY5cKNP7ynjtSv58sOJW/0eIOtPi
3dOsA/Vrux7DYz642suuYim+IscVp4cvwhYJoZIc99db/zMp3wsWmf1TBA+Pf2/tow+VhfjWdGkd
IFSDHS135UCDKrlCBjaN9O1aQDHEgcfYXE9dRUFPAokEuZc0sJfxErOpe02Y4ow+X39AGYN0Ut9s
uNzIP/J9ykgu+CSrOBaEvv8zMkzz3/YzEt5D7TQVDF0wZ/LGwb7gMKNdaJ4lJ6AKaAkBTjFj9LJd
ujiIauE0ogS0HF49gNhoyMzwCK8uNWMLVlhZ4WLYIrvcgNcBwUxthHXWS7MdmqnVwgCKrI+d8j3a
7I9Zl1FU2QKDACY5ItYWmTzY2SkaVoPjQ4IY2cfk66aqSZtW64m37N0ZZzAtFgAW82iV3UVkysyN
dUGLrLLpfmM0lSfDLj+IjZZbR+9+VKIaCNlUv276N9+byoMFHFmNl89pKTSdk+v1mnUBm5YcbocF
FaBkQvzEg3+Bm4oclcRhmtWKWiHbNWD6THhVTE+zGaYSL3AEdjF0UlIt3EJ8xcnn4YwEvjtowG9h
pKLbM95Hw8dPO3MOMN6aLjUU9p7m3fOA43n+Xo17rbzfeQm9tACSR8E571c1l/ZRL3exHTxrIi1I
U39QAeo2DXezzu/vqiduiKqULQZ2F2zuo7dc5o91ZIJ4UrhYLl/EbIwArOpFDyH0rL8SrB7I8K1J
QnZobc4mSMpX6gLCz8oIPXGF9og+voOpWZmYveGm5T8uaVIjCBoA5qa8Uu8RJnzDY62uQhGo3EsS
UrMLJcAWweaGQ8vSymTXDeaP0oIA0aaiFyka4aIwEinXCtacfmRH+b43eGsbPxQVEmXiZbN73qRj
qFFi+judgzn24dJZHNkg3XvUoNhRhD/FlsjH9qGyTUJdjJ1soZZb3wseYGmUwDOUv36xYF5zOsnY
0R6cRmjH+sXqv+Ch9G+PzBu6HDDFD5v9xDJngUFSK3tYfNq8ayFEep2Y+9QPH25Ag8Bx46q8lGTC
Xv/GwJONNidT3vddJQ6WIgubnwegVxRJe29mfN7LnJi8OUOSOUwGFhq2Jhry+DMkeytPO7vgS9MO
weRe3grLwd/2Pck3ENSozvwGPS3tQRcmqR9wpyOAUA8cN/2gDq8i5c7I1LjewNEkaf2v90SdOGcu
smBA/j+RnwB98AcR5DEjhem0B3k+ZmwaItmYcrIX6Nbg7Py4XZwUJjG5bM2fNS8vDB7GEIwFuo+B
x6LnpJsydMbarSs2yyW3NyYuFL/Y1ytrcBJDFbpOv7zl3fxF2UpNZkd6RDOxO71Ujzk7dYrS/Mvp
LS7f5mYvJNCwZor1ocfwI1oEqVVtMzj62Zle7CmIVGLn9z9frPy5nim7PJGgoROATVbY8xkDkv7D
YUdMNR7IftEX381RH6uRnpOgoK+0A0PJTAyUMtH6TSeZ5xgpQbUmEOo8yCGxTfT1BeInNMz3R2ij
/rPt7BAO+kRF3bq6X1umqVnUb7iv+9/NXcJNZN4UQfZYpz+rsQ/sGkBX+3oVQBU2JWxUXNCif3MH
bX+ygt9Sd6O+xAI8cm3js89j75lTit7HbfgFD1OqvnWGUpz8s5hY8L8znl/F5IoMUBoWgCrwrGn9
jJfhcetaXpCURKO5YE8v/aShn1CjV32BLxuYtJGtIE35wbv+WpdJy3C/48T806Q/R3lJBICgwhN2
5mjFEJhN8uqLvsiPjjRn5mGkrvCNufABQ0ThGonTZMuKNRavPt/4lEzeodrIn+3Kyn/NsTVWoSE5
rs/9ErmsKJA8s6mnV3AHVg/3sqmQv/0ghpTt2j4mNlyOgz9OhI2k1V6mNK8JtEvKyaelbTKr5X9c
f68fQMdBc6yq2aHjhHOMWTffWV5omF+VtoebO6YDuqMKs3r8qNBbnPoLFMz4JfGCWqe3KIqUJljB
MzmJbT/aXhtkjg5tOtwaEGg8qAbH9UcKF3GTv0oIeyEz1H12vpsrTgXs8+F1eSkexXm50q6NLyib
AYImmACLXcGvgOXnLA9r6qKAqsLudqGS1d3HFEDmYLkdDKdPKC8W1Kyk1eJyqBcPkHga5vxNv8lP
3cQAbWLlpBSlgK9SFOdMzyoQqjSdhQXEbAdKccyDE0Vd/mTZZkE37q79Rs00bn3ACAMn+/7cLnA/
P969l469TQBvqN4lN5ox6uKyp4WBL8L9RZwpK3PzkynP4rquzoSiA57CeiEIoV2OpO2v3ixJXyGz
tc5xkTslwuJDRyYKvL/czGf6rKA4+uvrPgF6oEBd6n21dWB0TF61GvIi88YHT3tgL629wxpMEtIn
clANsVZoZfmYksPc5MiNnRegrcFND7hj/jwUtnT9OgUP0ZQZ8GD9VRihgpUMn7hESh70O3fxG5v0
ooBdpu7kFOysvEtYWTj2bLS1WkelZZVIRtVfTn2m/h8UDgZpFAz5nAKS+bGnfjx7VXbIEdDzjFDu
VjhfAkBYijpIVPxemjb6kuVILEtKLdSKck5uWKhEA7niY3MDcJq6DbuUO4xl1fNHpq/vm3WDxnMB
yxg0GkBpHwj8XLc6mx0OZRZ+dBRizkct/nfz13/2DDkjWcYf38EH/rlnybXXlyoUwwMR1U4o3gL8
vgK+acpdNlAylo7u4pSuJB06Dn9y0fHHKlFVUArSDFFDSsJIGxX8g++qyOu1/wLiYrkXivX2ZpQT
gP2+GgEgf/yZ1xhUGKKXVbk8Pm2117e2bNnzYq8PfQN9Q5kMqLcoEJMhevCyhgCEug5t6MIPoNwV
5Dnui9TQuzLUwnd9Q94uK+CLvKFstVvpYaCIJl23bC+i6K6LnU+CMwv0SnBJOoKdp58q0iUKRZXv
8O9YqXiBhpyybtXeNgh+xTRqDc/W2rGkNnyFtv9gShbOiH8d92Xo5h8YBMq37c/zasqtchQmRmKK
yLcKwdzOyINZ7sLOZcJCitzAYYZ7P5lDAE5ADVQFKgEKpK9Oek2ERocVEvodkP6hQCZIo8ng4zFF
o75/XBAmEcurjF5i6HVMwxr3g7Ij9AF1Mv0KsaWYE+xoj9kSdgBzSpp7wTETaAoU1y2IcQfr40bh
vK8eDSPS8n6KcC0LrBg3TYDbd/P8ZhW30n6vNdoAObA2+Mjp26ffmw96AmRV40qv/aZelXUYH5vk
/heFoSwJiwldT2+/ZEPXn0D40r3nJVx3hpksQLUkrtoyar6mWrD9QkIIZv+TTpdXGOsU1vJOAqny
m2EoZ0tUZtScCt1IrHBx1VM80DIY7V0spuTkW66fIXYQ+EWI1G2RUSm0I3Vkdo1aujxeeFRXkl8Z
eM0iSl6FcqmZroUpzEToJTx1WAxJkU1RHN+X1RiQGITQtayY0nfdasfs/FklO8U3Og8thdwXrgxX
Bda5vJ8XH3vdcIHjeK8BYUu95iXB37pga8iDj8yoyUwL8Ou4VtSrC6LMV3zfkKHKLmXcyhm2L5OO
JI06V+e3r9NnBqF0FxAKBAHarU+ZRv+6nq2hpWz+koXAwwIlblu/GJ18lf7RBYc7YuAF24W6PSsM
7slm/Vp2uBc5zjXnVtDKk+7Y6vjOYu1/2NLxEufIbyN4mY60NX4XGv2+0NF7zqjBFKpIOPrnyyfp
lCN9ZT1sRNOV5Eu9w8kxI70SA9qDoU7IBQeSBRxeV7K5ysNj9jgkXesHFXHcBRLJpE5j6y9GdpYS
21cjAVqtw4+kvUmLAY3wv+v4Era9GTe5ltR0paBlny83Sjm4YlAiavo79TKtKFi8RRHroCAnNqU1
4jHSukQkITbfWUPTm+tVHyAv0Mwa6cRpxnDc5JlUzQ4AwK3nnyZNX3IJC9zZxR/CMFnKOfFYa6SG
HKlBglZV6jSnKAsJNQtibcJvhR1PzrQS3BALxVujYGbOnLHfbEkFQobRwd3Mt9AQaSDFzBEJK7nc
IfWklVzsxmeXP7EdtTLCqQefgYbwRNs560g2zQtq4/bBTTqP6LvcCuMA4I7/qt344BBxfghtU5KM
whycqEQcyr8CR86qg785RYC5c7ksBBtSfYYWPZ1r/c0IE5Ds3avU6frrml7zFRXmyI0H1s3xu1mo
alVCe7uqmBSCn1SBX1i6F+FtB91ktCoP92ApUT/q8TRmeyEdwd1YFSfXPXwkzmY9xev81DnEkkWy
XKC3gSo8GW7D9OoFlKeMxhrM7JD8243ZBWXaaAPW94sM5s9DjlpZjihE2ETUS8l1TMlPbqF0AWCC
FYGxtKVHY4nyTEfu3oMKYmzGzNNocPtxNoXU1pycF5pcS9SpgAEiHTc+zLO43e9JjfEQadDcb8u7
82tLRrdpggc0CuQAbZWyphmZNqoIpzcsTGAhNyNz0xHVJpfg/OINdgEh023wyqQ6wPtP4eRV6TYm
RoS633eidFBKvVZFYS+up9D+DOQkJqRXdo7F0XystoMeJIE7Vj5lOWJY8Hae11cMjrIr8sTqTfrQ
KpOGB2/9XI36T32E/oK6qTDPEYJOwgQQgTWMyGldJhYh57iFwdNn2Lvo8fAK4kocjoDD7SDUyoue
L7cMs2ypSZvj2Q5vQJvKUHUMdBWvW8LDNk2Oh/TX3VCF78s1/GgYia7+uzUM17AUFaksiJ4EirhG
Ia7uFcS+YDGx4hGM4e4cVJedSiV2163VKcJQKIISM3gxWbcqNy7G2EP2cUII6b+5W8+oW3Renz8M
rbbxuPawUxn33ltZsKcgFZFRQsSCZWYOZYdtf9SV2NqtujnZYX5sec65R95qdbjNAQbVpyYs+qcP
myUiAJPhipqiNJr+mJfV4TYSy2OwQmHgGTjm15V0ryEBKfqvv0G9mADAaYi4ISrwxSKq7TyqJn1T
7p6w1zhpGLZMN6ZNe1UAUo6jMIedmcltdChFLcEPDreGc1H3Q7SyPLoMjSHtnNfXF7UajymP1cIY
L8v5kAaFMF6YrzdL9f9QUbACBH8oZTSvFzrtrQhkbdeoHjEldveXJR7G0BhqqVTjO4PHVHNUoeni
A1D639w4hEcAxLdGnOLBQ0gcsHQGeYhrzrCi61jNiaY2DWzxyszIW6KSOi3YPv3gBp3dQyPCVbke
GYzUEXZ3QEaOgspng5phr+m/bKL8uk511lMiWAo1d6rtgYOQnJarVnGH5ih9cnvSr3NuKlvt/Ou1
ffZGvfwlBLNHZFvxP4FqKR+wkw51ZKQjqB2i7+yl7ky7oCAdWC2IsMe+FF93Vf051GTGxkkaYMy2
mMDq04jWXWjweOGuGKDYCYRL3N469ph/WmMzRL9CEh/zrnt5LXdTMsBXC8aSx4EEmGepazyx802U
WB9cl2tXLwj5PnhmW5M11w197laKKwN0/kS1oS/Vst6ey2qC8uIeDD/MYTVxdtIMRhIUYbEeSm/y
BhcJjdWWcYcFdW1wuvTPL9/bpRtLdi2dQ3JfUBzCFrFwJa3y6CUM4Q9AldISWzA7uHu7oTQIl1iA
JGlDljmfs7NuW+00AOjquIPGyJo+AOV5wwOXYKTA1mmfxrm7UEkXs+vhJ6GcG+//Df0Vfl/UKzXC
yhKAFSK7Kf43H4GNs86LOAx11Sq4RepEVk/RFWPYUQQklK4mbGdaevKRacPc6HKwP1dGPmR7Pb3x
PYAEj+lfwbvvl1VW1f3BBd+gQSo8QKUEAzzzdVagCq5cbwVvOX9G7T6WZDFSAK6I5n79Q38zvybV
LPXIKNVFvSGah8rpm9jK/BDIKbCcKMz01J4CIyQHxWuzXzfzEo/7ohlmUgWO//8WcaIZum0zN19n
ZUG5lL/+U1zO6Sru/WqUCt9nlWPcOyhjUUI5tj0xvcQVcGR83EekZcczdn2O0jwhurK3fltBNTqe
xh61cxpzZ5qbz8urboRlAOu9Qwcz86Zla7gl4SVRxcylYiaSBWzhdOTNMZB+//OqxxKRVRkCkWg4
Y8LMeCDp4+Z5Hy3O4DDHq0jBBTJ+YtMZ6mcSRMVBLJZck5irK2WHjJuAQKMeeDSB7UZxg/XQGWj8
7yqqUJ7SfEuQn/hkvF2Ep8ul4fywLhmjDDuEVk1Kvm34Oyt+NnUcGpbxyqpoeU4yC5UU6eTnNQWb
kauifRgsPaR+SfLxwGUa+jx7jPTEbF2aEMS0WSM+GKm7eycDq/hPakCmxg1LuZRer+v6nQB+CBIo
FUyMzd9dW9PK6js5kAjLR1V8953GZZNmCBv1Rjf5OCWOwE0OAZfpY+eYjx2sP2qqXDonvFwKjjS/
7pDG+mQRsz0kQVhvsNxzMYMUul8ItKeKi31Avow0dN/B8XSzLAocAPAEoFh0pN3hyYka11iLzB+m
/RsRLhiHOjvA/9nxSJkQrV//yyD3T+ti9cF06jzqzxsjlVq+E4YwppR0p4MoGwCiSV+JOxT3InBJ
WY+ZPEGaYyg6pMKS/9VTsuidzmzPHnd7hJEK2Mq4tBUlpXd2054/jKM4JEAuypfUHuhpVrG44ISm
9LIJDJPNCMWkihMNv7TpCynB1otq1nwh/yflL9oZL1Md/+gNfNdK9YmqgdIcdTVfM4TL/uSAec3t
3y0I8gtfATRp+RYTHjutQT0Aa9nLNN/KSkPHqe0K2dVPzElAj+Iz0bbB9JQWmla28wgBI8TmZqs1
pLgfZCsW+ULfcrvVjndFVjbhZvflZIhReAvG+yIvqpwXmrg5Qk6syMzTdCXa4OVyG+Vy93dWJ4iJ
qTmCRTV7WD2R4vk0+9zOk5i6Q5rNm0zbuUSto3DhwkbO00jdcSmKm/Ko2nQmVnJMyW7WVGj22HeW
4+ELiEFR05CK8gM20Pbr0gkkQiEtUvg/kDDyucNAhNpiFVQsXixHIBGCDwZOkRPl4+dOmI2zJEBE
zjuqGODXM0buqnvhvQwrK3eqWpAeYpniMMMwuHgfT6tWvyogg5LjQrmqNFvzMlAAML1RIjlImOPB
LFKDirhL+cV5Nryccv2crG6tHTVeDqqVh9Ccc1AoZWsfKHHUQcBvFtYJj/3XAjGGORKRGp7nijXR
vEyz43kf6zTtjygjoVE8y6fr39qBCtW8E0DhyUdCoD3mLU97s5tH8zJpn5jP6ncxJoRhYQMVm66f
bATJxHW7y60903VqZhF1tcvFOjWRx+KmIpa8aUCSC/8TAmRM+pm5E6SWoxTJ0NVML6Sf7qPxGjGF
1VXlolc+ke+3Ew8o5TYwn5njetX4wS9IxHoyB1BMmfxnlOroc0RjnHFBtQygcWgm5yxUImJ9WPyW
N686aieZUYN2mkjHF0+8izmGCUiARrrWouYxAgmQyVAAOBRMXYFY39EIQ15H4jr+EdDVNc3kM6To
CK6quf672cCG3henpY5ndcuwxEBO8+856zL94JrR1oc4o6Ekso6jpWiL1sAMblWQxE94jBmE4K6m
Af05GpsLER6TbzN+0MwUbZI1GvdqGPw79ADYkMSWLyOQ3uxRmeBDw38+quRwUYafshmgevlXPjW3
387B4Pfqxq9sbqB3oCyPlTbKz0F2WW8jzaRbtd4CUZWACRfjtEuwH3Q1aRTf4urAR03ONSUm+4C3
c636QrmCsBa4l+Rd8ew+GxFpd97SN30rcCuSOde6QCXXbkTNCnNBDjSj+erIoyT/+OQPy0hSUD8A
P/AxI+ENufjOkGDHO/wG7yzwd9/yTZNkMTWpY4kcYX4n9qm8T5m/gfFYHxOeuvZYraOHTHjc2Qnq
UZ0wqbUMN8jrDB/lGihg7hjpH73maNBdfrtUI8NzkYB0qcjNgE/pVCK3gorEcDmYXIUZTqFcULuR
dCNfjS2iEUCtxychhIBWAZcftC66RnCjXcIf7os6vKcDHXWglt4Mmy1dD2gprHfWgr4XN4IRq2gG
7aPOh1oJop9hWJK96/ifR63REEG+E4ZO5HHhfa/rooYJkAxkQ9XgwP3mH7DWeK0dsngop2nEGaBS
k+775Gmoez9jmeJmvzXylmkn+jf5CfSNOcYijcDBMOTF/nEU0WSEBXgZ7J9pKgyCYtRLlSpMAsvo
gY1kOQURhf/jRihBYUPt7keEasfuroGWgXjXrsQfQjD3MdcqbzKbxo6bzmME6DPUXFtLLOYGMBrp
qz24LLdEcWd7IKuR81KWMvnPOF1csTuieAj8KQHaLWcmQx2m9hy1izeq/gohBSfCBzKxgQ7LQ9XR
w9kg0K76MojO0B9iumCrwBT7X15VZravWSmN76T1mG4M9VbYrMOJGpkH55FISl3LV84sGkrxb+oI
PNOXqCRYftmqnhCMcPDZw2XXTFY9Xwh/YlIbDAKUuj9ugviLLZ1HEd9uBMNIDNcC0I69ozCuYZr/
568ysuB8lUnVy46KpZ6Jbz7ynMVoZQF+JmPonEG6/HmdMf7VHfHOb0yGym4IAT70bys2ci+em2GF
TkmPZRjSlIDciM9+TMrRNPiFvNZ0KMugAbdnySxifSw/jNSAPIQweFh3vnSskOaMiJXab/zyyriQ
+u2clKqOWToXy0aYo94f65rdCFptBzzzVaDBKjg0AveTfkp5mpzn0Tb9yyEpnL1abu2vY7Map7Ak
UhUrEZOk/gYS40sYQBsroPRiMWw9WKT2FArrLMII4PWzmlTQ47xsnqsR2V5MIdriPSo1YlUbAKPb
VvisZmYXptPupjDvdUB75UEsn9X47JMAaMrKToeGp/7s7m324EiZwIFBBPG5fPAezrnzia1aF9Y5
S9iQ86eZiV9MR+I7OiSioImqDqDXoJNItBAWds2KKDXgbosHweZJXLbWjQvi8WTymPM0GmiQxGcy
7jnjp0WUCLcNqHlNXySk3NQaeYZZMmoRPheV6i+7smM37frxM/L+xICjXqqSK32JFSNYSELstI5g
ZqSHbYLrGT1rqPQs/g97oTv70halQclbjtby9JNiTXqWJXU2fkWkWz1chcw2nZQaswohOFtCevIU
Ctj1uRrR0AC2+PqznYCteuMJtVG9kh6t4FjGh7GmcDq9Zkb2PwuNuj73XGWqiB4uHrKsRpcE3Aez
kYqf+axnOyEP9tHdJ/BvNCoKAdb5eUtCrwm6NeCuQUbkPebvHwimCN8uUxrjglmD4rbq6+IetlZU
1zSUOb1E52lxuuq72A1fTfXaNBJ0pYA8WbfO+WUL5xyrjVLPK2Cmeq1RtkiaJJJ4xLHUMYzTVXNk
9krOrGlACvQUIrf/UErva7r3NXCkrNIJfYcu3svchl1MN+XZItJNL11fnnSaI4tqFTNFekq4gT0V
9uy66r5QnrwOzHShAy7e+/b6qMWknUjMNSaPMHnLrMiUKc8fIXufNRV6KbC65TVVqx3CZRzbHT56
yoMOfGdxOvu7SWiGVzn5V+UAQuUK5OTNQWpAszdBXfWHKSChZeQSAR0KeT1Un7GvxqNvqamFGq4A
Cdaquwzp02Qsoa/2da7+YbxllT1/KVc4Exb3U2ywYfR8+Ct+8DQPPGnHyd2WWj47Nyw2BMF6/D1L
L3rLETX+kEueUDlOOhuh1j6wyh9wFuBcXuHWlcp5xkAH3GO1tYlxURe7GOd80yeakjLaOPkOSvgD
IcKbXDF56zY719ATXzWxZ7j/OanrUNu1f3BbRLOlZbEfuq3zqzIq0YJq+uHX2UaAJJoYN2wrBAKf
X8a9BZ8lEbveV79v13rVkIwdKGrQI1vVkaBdGH6XoD7K4jNkxdMfihpit5nsBl43U7Br+hS+hA+s
whzAn1W7tEOc2EYiuQb/mFGvnK00M70nWhoBsUWJkueTvHxzj+Y1lLcXR1vIn6oJ9/LABPVPrJ9K
ylRbcxuvtkQHdFGt2TxvukJQYwAM7/IBwZEse1zz6dTWhjktwAV/UJqKMBYj96eLTzOZ+xflLQ3y
58D46Q6f4k4WlDfA07c4EJB557O9thDYVrJhoDHOUvrMZQ5u7edp7eCHBTTLlrkGiWEAgIGeyrDe
pHnz3L9UumD0OUPa8Dt3AE0ja6mfr8PJ5wJ9U9CFBUyDP2mGnzEWHirEffp2d0+7ZqJ+LyOvE9Lc
edKGpqVwXl3BuDJ2hwJpyilsILhvYwhd7p/BxNyQwy4FkbpgQ9D+pieQ+Uuyb3qN9eLPe0HZ/Ogy
krpMFoXOPKprSWl5KuFaGK2ZOaMHkeFnb7QfeLdWlewVd0Idm/QAO+hRmCAcrKDoyXg5bbq39kHR
+m9PToh04GeAiRR/PSPK+pxA/6GMQ9TzQiEIszV108dvZJAUVEFPIKZCRzvrLsjAUA/cBRvf2m7I
XUsAuRJb/YcGRiq/3QdcwVKkMfPbi5GrHvUbqgEnug/f6XgQPmntqn/DGu/4pQi9wLIu5frvHvYq
ZZoz0c3ia19xJS65swYXmMuWw1GHCvdHl8iDvbADwpfddocsNij79TFDTOmJpY5A3mXyXLoY1+YN
ggummny93C0EITrhVjjPAsZy7K22dchf2G4Z66INmCJP7rCDncHsKA8oWxNeeWjMGgeFU+GX40hL
m4CiRMkNzrLq3dWEJHQ1DbVNC1V+pgJFRTFIc3wSSVR+xQytkOjU7Fz2w2g3Eh+a1xqr2MwGtBxB
ZmJ6tmWt7bVC2I9gLNMdFv/G+niYo4w2qw9EBmrLdTRHsbsa8yzFAcrafCwHPVmZesb1l5tnTwir
UUlfS5y8h7H11Yu9jCPDaBKXdoEQnJD5N3mWDjkcXmq2WFJP8a2SESj61tsrqXZkuvboXBwXvr1b
s0RigwHnK1/RS6f2ljMZVCtEF+9Ah06IlXkdZ+ioDOPxkcFfwHaiRD9IUAQlinbqxgR5KCqc9x3Y
45eejks7czBp5mX9rNwH2LWi5L7mWNPL+WGwHHXOlA1OAqGP7hKSWHO8LpF9um+B8og1eompm4bO
0vUnWWPo0VXqNNH7zcvDGQFllNjku+YZSiKLtrnOpB4npN+v1biDlNFte4gju0TEIPrs4LQLEX9j
1Rq58064GLrIrq8HvnWNbEiRRPCDgy5XI86UuoJrssRcR9aKIkkNqJVH74dulZsMKWbtS5yO+g05
BYXDKU3ZJgDl2do5H3BGHb7RMapwe4GimyCcszzgVDGF8iAv/jGJddF6BzI2m6ViMGX/jPdguoWa
mSgqYQI9rb1TF+ZQJUN5QKPm5SaqPJpTUymLZInsEbF8yR31PFIJkN9ziw95uCkA0Xd++QIKSSYk
1qsZhzIem5K9hrgMMIYp/LlPTIwwLCF8ZLmo1HK1TZ0CUlnpi8ZJDskpzEgfu+vtvA/5JjWHkl1E
X9DNx2nCWzGgKRHlAALK2oI2NJoBmPUpMZEyTsiXo532rDxSvxyPK+hZD9Aq1Xt+pRv7FYKSKCLe
IxYMqe0wO2E54fETsEHJqS5u6LMLM/7UaAx6pIvaY7BdH13O2XgkOEiOTWUZnPQ5EEwW9D14qwdU
H388TCg1Ym0pKsGHXHfemBAb3tSSt/mDeAcDDmEE3NBBlB1VN+WStodTRtlVqB2luRVyF3srGwnA
gWy9Emks9vQi/lF7XGy36+QMHgUNdx+FuTIDByeYlPIPl76X/NZvpSUbcOgUizVn6Mnexl50++NP
ALwGbUQ0fmoOOCiCdEIxesL1txEac88qgbXVR86A+49JVLVqnYfhY/iGI8m+MIJLR72bKn34K0qk
IrLJ6B5z1CfxoBnMLuSpHVtf9K4Z8JMLFeI4AN1ufSl1bozi/OR+RLfF+7cxSpVVbfxdYMphV2jO
T0juM3O5VB/RNulROgH/jh3ifyYqyRCbKngmh5rte+kcmfUQ0QLEnS4wThRFIbIRLo367918JYGK
FKLyW7qwq4RauSGkh817nzJodtklEWHnhk2UHoQEt1+B17soRDWZQpaRZFMYujb4Umq5y0eivPUr
UJYlTXfysyjPT7GRNsKQTs/SRUy3tGfvbP3AOOwcSzHjnz4v17hYdy2Zs7F6X5yj40PbkN6gz9Dj
ujeftN0gVz8yfcBlN19ZK9t9DGomGJFXh5VqyzWzfj31yDb9nLFqQwZ24Xy1MLDiqM9b0psNkdOX
wQl98ZSHhgHq2us5iVqyb/ZFcg4RefWvNSazc5RQkRYBaIo2LG4huoBwk5cEmfQVrNmJ8Hqhnf7f
I8L7Y08nCLFOMfR6bDwQAcGs6RJVKSE713saJuVtDJaONi8BpWMWwLB0y3gYmsJhkbogvGYli54O
OkDk4/jK6YmEg2oThcPmVPVQqRisNLbvsfIh6u5vbfkigqkP/yf/rx/bnjSwYWBYXLr4dCUlEloD
5mJ6GDWF1wkJyeZBYnQH6mHWGOFb19Xe6NSTHhA5FHDGTmIu3V1mL1qTTNDe6M7N1j8APsMaeI+t
kRPnlXHWriKCpVq74ICZr6VDTXJcIa3doczLbEkA60s9xNgNwVSxr/32NuvHUvZvfZKOrVTU19H+
h/8GYLFR7Xq301fH4LkwkU2WYrv7X3NGiFTWV7iuFB3MWKxds9Gjj+4Ri8l+3XaX4miwBc2TKa7d
sLZxfBx35oShYmByjWBAWXTa2TFUSL2s8ojViPiO1LsR6WAGbUYe//oQ7xeGI6lLyAORgZ5l7jat
INON0OkE92m/0UAW/YTSdjZEFfryrN3AwmkQifRKw/LxXS/vG4beiy/kwk2JPDKcdkt+jlo38a+k
esa6DVpL42rX3P0xTlv+rtun42hj3BowEdGRnF69vd1J1683XDKG3K4pVvq3HJOvlXgwU1Sim1Mj
pG/TE1E4eq551vCjzUGiOIPE7OvDAJRggge3aYwyIthN2zdr5hWiL/kgUqLFWov2TWIfaB9czps8
mFkUQABwrq5eskWpbODmRTiMeVjJIKCn/NDJx3vXMYM4hPn5DAZcuY2Ufi+pBaSYi9Ol4H8F1itD
uW53y/ig9RnQzHpVSuwJ8DubZKwQQrY3mYynkxQFBDTiiERYmT0uzne6h7XDUna2vU6AZ7Itl5O1
HfMi2cj02/pEDNvEblt+Mr4F71xU5+BUwL0sMhGSUra2eyENsI5O5RaiY+mq6qmAe8DxC0LHrcyJ
jLofqgBcPCCinh6dqQDvYU5wGrmkF2bbI0ySPfmZ+K/ATt6tNS52u3U+Jvhlmk6nnleiJ5QDH/0e
sMM4alau+v3KzbDl05qO1ITOu2BYsMuL2Sdg68Inz5Rn+dDaPmseUn41JDG1rcKA/YKoFPk+APBr
ryLbrrnWehgECKZUdciOiXtUJ8U9Dyr9SVgTmQfNL6rJqargVFnR4OPX9yUxd++NRKOY/bKQNVsu
sw3owDEFJ820ZxSYUnj/5aBvpkn0rzVtbN8J/kVq3S6nc02wegONJJDDfcdxT01u8PL8gk2+rqft
XBrrscPmY1UKNnaVlttCc0L5dP4mHAhcLWqqegK8IkcP/ricShfPZni/cNAzSR2QuIvpOyf3xivL
VuvAxEKeGCXrjrt9Q0FSj4eWoh/S3sCL3ZhVaRGqDdA2WbJzwuB53M/kEXh2Bjw6aLRJAmxprE/N
JYY0HhZWgp/3dbJuT3sLlhdrEsN+HmEHEsIKgPYcuUrP76OlkZGKyECWk7upZpK30GGtG8I/zVfw
/Cla2ckMFPk6o0tKZJvsSemphpzhMIr5DMojy40rBXnkHoPkSPxISb+9VHdW+bydVipd1ALpLFsi
c/bv0pHX3MdNosYFsmO79NwBsF20Ix011cKROyW+d9rX/HTC3Ot2RdaVQxuIm3eFDJgGmu34rp8j
wJpmTeWsjMMIUs2JsMUn50MLCwmq0E5s6wKWmkU4usyf+mZYTbGl1bX++RJ4qs/hRocPE4tiiAhx
wCNTLRhu/i1wnfPbELj5lNRYXhMqB4GKKyqTzqhmSBGQQHIpyb/D10B4nCCer3vPbqkf8xLfpgEg
95827EKzIxFYf82fakbT+vQ8dDaXpaPz9KrPdAeSj+fWCYA1Qm+OCAkyhoRGn8EXjvPZqiEObgxb
QJdWmoQiZkSHSBugJU8PjrVPs0PCteKk+2YRmViW1slGdTy8LSuOMJX91yQ0rk7ExZSBSntxB5DV
K8WsA7QwbipIthsaaBsd9PU/8gXFAuqzYadhhdol0SNvx3h+Ec7zYrJHhOLy0OCk1lD23KDxF+Iz
behTv7q9HHltTLmpLvVRQozosdtDuFAMHBJa/n8dbkIwskY/v0fXjV4FSYXbK/Uz/5KWfYQ+Niiw
JOZlpendy6NUukr4uEKk8rhuFk3GVlLxN+ipdCI4RAyyY8IKSldcn3e0wHVsYKDpStt/0rJuiHbJ
JptBXpK5+jpdzSbM2qCM2ymEK5OcKxFYcBeIxtDydvMO2XmLDQqZ/4ZTVMdXpp3uV2LmEq5diHPJ
9QJKAbJ5AmQ0bkkJa1M1jKyiEa+o2thIAQ5kAKV4BTNkKiVN9mv/75ijSBqqpZqZNRl6gj5+zkCT
wvaCfQFQA0ZdJl3AkkLDVs5gUm46Bfu3QRwT3ViqhYrFdMyJ4IXkwK0RnlRQwaEDuXFOKfH4/gTu
08MvXs2zZ83IJX4FdegV+8TsNofJDJ6yLJQaaiUxKEVOkeCmUl3n4MgQihWzu+n1UsY7h9hMH+F8
+T6vdtEkhNHPMHKL7PODR1IwosbzfiK64i2WwTJwF/5IFIUiyKFFAyYFQ7cS9oU7UZF4g5qmVeZ8
ROYyDh5TzVPH3UB+dJJppqJkm+8w2GE8ZB4qDoaIVS1KJTM/fXwwAqSEzX49v7o3L+nXd79yEvWU
vDPYw8upu/dNYe6eagnDA6VTlI3nXYfItgaPl0aLw/f7tMkOwUae2f1ThMsp9ZUBfGpsLF3Rn5cj
xklOhwEQlyOP4yL12oz9FlVzM+ouYSXoD7inPFag0aUqqlk5c3YmV0DG52HbxdI1F7Nq4YL/xyH1
fw92gA8Ku38A4DAPyRwqBdbrOGcTdRDH8SNSJsFvOU6I86zRJM1NFDDNBuTRmVGnKFGO0MeKTzcH
J0td/jUPaX4O0qwdUmXukZbUYGE3DjhZpl9GSLiLYqiGXe1yfSz6QTe8Zk247MVA4F+A1oSdMi/5
8KEd/En7KifhNKKGmsep8rxHC/M2YFaFq1arrJT+zPYDrar38Ndgl3t2uFZuhzPhS9WGW91WAPyV
Pyk1dgjxP/Yat/azhSlAz8Id6/Z6Oy3NWmnDOPynDp6Col7iO6aPS7WFVOKlTEm3ZfZtrGwwM/6q
ptL4IE/lSEa/s2Q1qHgFsfj7A1XhccdNHNIKIPk3marJHYPLIjKJKJAErfmWsgc5zq8qFYZ+RE8N
O/ST3Nd61Ndw0JTFvoBWsEnPHK3BsNsDwl5dWpqsaNn9WH+RV4Y/+kgQ0JUrfiNugGgJjmzmi2TQ
WwmJmBAsv3E93Oc5f1v3bDYRCj0WAXPut2bSHvYvY0XdAgiRrqyPALFri0kbz0xFXNsjjEJSLN/h
UCEr+vvPl4x9BiZnLW7668OZbgwaI+XG+pYOWXmyxAdFR1trkHOif33RtFlQQg3FoIlAetqGLYXo
YlxhQKQacRa4/HVazw8E6jpbutNDULI2VNxt1gZkXQ0IniLALRlsA008cSHYrkWg5iIlTpNVD7WJ
M7Ilg/3nbZWaSS7KtTX7ugQSjcr3GhUGv8yIxzsP5c6Ya9ltNUsd2nhIT0BpnRj4d6EKgrL7mqQz
cokJIWYqhW+/8aCM1fNerQWiIDcGUWLcVkE/uTeWA3H3YcoK4BbuZhiPR5nsjsxNgzvB/ZpiVi+Q
A0FKVIvwb/3+YI50k+wQjN26UWys272ps2+2QI7B8EsC/2sFtyN00BCvKCbuH4BQ4ovqSKl2YZ4Z
1lCMg+jdtU8DXIsUTCsnI2gA5Y4pyt35NZU0LuhuHYAsohkAajbRcwHRqed0BmZ5OXWoMwLjsnB9
j1arhtQFt5vnPAITgAQFgdW5i98Lm/54hPLTg7B4sXKo8M1PDISmCR0BvtXXOah13RCY8uyCvdMP
yjTYCRDguS7dzxVbLUUwGxM1UE3i4S4qnlBfULHSxpwqtw1DCwEvDqT7Z7Y19Q7Ch0OLRPVc1VRk
YeB1u4oKCajxwpARzCyPmqvWTDYgyX17wVS7IUeljQVUsU0Hra0hpg+ggcaPRSev0/QLjYc4k6s+
9BJ0sdDOdeBtnCSrLW9MIJRRBUeAOonePW+nNbGlWumcjrZ1FBopIa1QxH/VRkt3rP8LyA6DUK1P
9MRmoA+5csAjFnZAAOHhpJFayQAwCumBcgo0EfSW8qPUDrtbD1X7YAm/pSRKdKT2WUuCQCAMlADS
yuTECoZwcrsGSyR1NVqLySVFXKGa0zMfY5XKVDHY8bxBs4MV5OlS2peLxyvqlWJP6qyJWhfnTUes
qZ+RpLIgUrF5QWE7NY/Dk8zTq+ALpooHul4wdaM2tQm4fp7yF0Dr2Rio7piQ47e1SKL5URkNTDdW
Zb2FIe9umkHgggNS+uvbmSZR5u/gDyVcSxU0ByoSgEdjovFKgjl3NYOfyFJygYLmcGLsEhPxwdZK
V9zaPOm+GEUrSBmbBMPkQ3crAwnVisi693c6DS4WtddzDkBjDLvQHXOwSlmsdXpYelFtD4rjFG+A
aBqcE+UYdL84psvqBznJbgn/CkE4A4zULIGEbSlFQHc5G/u6FP2xdK9P2s1IUgXXKNEjb3oiG7db
g1eGtosMmviUWBPppxaiMYSY3dEfO5lVMTtus6vd3wBfMDB/lEHSyA0N3wMigvv2t5xmnuiHdv/G
yz5Ruh3NymmRKY149Xv/F/5O7NQtwEb4drMXu5ILhiCulPj9FbylTGRCbVAW8zVKaJW5zHWkHrEc
luPLoH0ctLUErqZX703u3fmTdp6c6PQ81rQ4JbNBSdzDqYVBhefG9aG3UOWs2iD9Q+hSnKKf1qzF
LexZdP2wysyvKVgw89y2yRhIu7OJF3ss099zT/Rk0yaKGXjnAK9cY5J6q7vy8AJQPX/yvugN5Zdr
VvFoUkdR1jmDkRlg8JECH+ItxHBXh3ZrKN8FhHMkn7YzHirj99+5zkgQR6xrkN1zjq+5zbku6FlQ
IeGKZMnkSutlhi8QoVasNUS15ypTt7CqM2HsY4XrCBJXAfeqwPDwEYW2GB05uDhTW/lQ4jwvhuRv
fgJY2/xUDEaa/8O+vIkKUfw6816siKRP4uv1PMSrO8pwXT9PF18eSovy44T5e4IlYBYqyvkgR/3m
C4kn3+Y4nBqMzrajPeRROX/FSwCXaxztiJF3N0l+jXB+M7Mch8sC72CKSogUOGK/sOJ3nuvFx7J9
xEKQaGdjg1up/VS3Few+g/0nxswTY/WKX6VDF6yQt97H6F4O847kBpindAqt/NbECyfT64qwtRCC
6HfjZrYcB278mhoXmdCCuqOLQCN5l/pAp81MZMipf6T3gDosCuI9gmm2T9a86iK1WRET6YLW1URY
X7twXV8vj30rbVHTC6X6QYE5gn8HfnKIq0Fg7x3a7KySVb9M9umoRUOi6wHWDk542Ljq9I4CaEuV
vLe7toGhApZgtDaWQfJofGpOaVlq5PFdcyUuv6uDQraCZaLB2RxlgRst7huiE3Hf5Q4VBz6LVsVy
MDYPPzMXbsBYMPEDs3pMLN4JsJCB1TOVSNlHz8aoZji1sFJ0X6zLK1AV6SGa6s3fzyeU/zUJXO8n
/EUIIMwZaicRj0ktPJuJnyFgsYvWTScDOOv339uYpwelku2WlnstXm61nYwRYEX3UkmRpafeGhBu
ExsA+EjqyxXBwoFIrc5TUz9D6Lbti34g2smVV2t6RVK6LGo7mYdAlFQ48KL7z4ttHPxW/mTLe/Ew
6QnwfwTeXXXGMzl7BwZ3rNGauW0m9MDavKMAao+XTTF4Pu05w8uaykO/dRLAOF5yc4fgjJQjMr4f
TwPV6O3+P3xg6lmMqblrnhLjX0LfbEv2Ho3VGlrBws0M8CYsSJjYo5aapBkpxDiNy7wc8ayrEfTp
A1k2cC8u9YrWeY0Yg4B3jzqeW8mdfxjA4BYas/own+XUZYuSrzX8d0gu8uyVzMvDr5Cj+irU3tZs
fDfqsX5JqREY+TOU8f1Mm1wzL5/Jv/euRRWg3a4Ebgmr82Hk6Y09sSkC8NdX0CwctkTC0E7CWIy1
D7ovXZh15ar/cHe1fXIo9e9cjc7mLaDN+hMpsVxKwDfKmdmXD3VDVBNVkR/0Cb5aqNTiFeBj8t0P
EZ8gEaYkwcZ2gaRPqMS5XrjAaxm5E2JdaDpI0EDWN/VdZfHSNLkSa52FgiZ6H5IdTQvLFH7Rl82t
7L1mkc0Edabq+aTyKSzaB/HIeXtZjWwjxU6BdfmUhvYBsMSPffxs6BRcRc+apjiYreUuS69/bVs4
Hwuxcl9PXvn2KvRzcsKaOGrNuymSVupyvOOvrng8mohER8C1VG/KQByPDzDuXnY6+EslJDMucaO3
3pnl0aeZBxTd55JXQrnauYU6ftIrlTvfLtJf5sOkfI9OI+KwR5vNLZLX5sec2cm/bO5qEhEWhdmS
rLvICJttEeO9CUosoA06WOWX8s9pMWFIJHMbKF1nMNAZnhVI1w/7lrjjhc2VKAhe06fInfvYc+6L
YB+Il8MwYUTDBMGu8bRXCnovpm+UrzoTt3d+9kxsIca6AGjTExPCJ4j7I5RTanJwC6RxhIwrc/DF
9GKtkbI+On63ctj6/PSB8zK5RkHILFMSsvvfr3fQJ43WYsewx08EcMNRh7Pm7KI/XxyqnKxdAqa2
wBS/4y4F4qUz6s5G6tqnDn/cD99rKRG6D1iaJZn2SzaN9A4pi4qbB31WPZry6ov3VFcZFLgT/8tI
owVKVJMygdwyO9VH1GM3vC8ibotTo7oYZx454bJFy27E0391MgiOBljzsGTUWci12QdleQTQXeYq
Z0MdWLuuzGcH7XT6gJDSuQ0uGR2KaBpRhK7JeMvySFhNckfc7wTja/XeLcwBkkKzXAi9WGPaM5lS
CB0uJ+5ZfhtdSHJlYTKMrsvULLHkJS2JqCMP+sfQqXtnWBq0AZHVw/8FaJ5gWqTZ1PQ9hYI8LzEd
ZJalOT6YpjIik+edI7jxLWzjuTktpU+flHltlNe+YT9o5CnD2OXkIQsusyzV5pbdwKm4b34jIord
ywbyQSweZY0yvTwRK05JkdG+LRc8++kCbxtm3x/fTC6PQOibxc9q5BrSnObgvcQj95xCxtbIZUg4
TtvuLHv3FnDQjHQdLn0EQ6WywK4XvqRti8C6LSZXype/UWNB9m7gAnrdx3EnarmsGsW4lYMTFCKA
ZV0PD1wYwXdu1k8pjpbwFMyYXKxO6ktBtVkzcNnR/KScyuIuARK62/VoGklmi02DgOup3B8qhxm6
os2rb0zIfzcFP7Z4vEJU/tn3z8ipLZt1Wi/sTl8TnsMgDVw56gSRa+fsRURUZDfD/NcuzmrD2lI+
tW0fHmsOvEtC5NxfmD55yH5mOTBvoYGBqUO7ZNOHCWg4AFk/NnYSImCBT/jYv2L0ZTNPcu1pZ3Jp
8VBerUPij0Lp/9oq8qGB7xM6RpX/NYHcNMhz7bBsrnqFc3qKthvLmUF3LY3+QZ8r2zc85BLDBIiG
9DpGHdZ5Err/gtIL8udcOktWz7gbl61j7p5kByIzyqRq1Jv+3FL4T6fDKq46KyoIN1j4lic7q9kG
82TXOivaOk1MjihCllwTcZ++EleHxtlXumIleDe0NqQm630consEAuxyHitj1A4k1lhiQX66kRoF
0/yczx9g+myFHOni2AkAhSZ9L7CxmxcBiJ4Hqs+lYb/Ro6fOe/9uHt1C5t7l19Wp0HQjBhOju5e2
fQOTua9pLGhkxaUYF025FT4Bm6X0P44vTh0vlq+RbmIoUxAK03S7RO6eT1pF8I3R+uu5+tO6VgO8
OuLWeOjaMga4c67t76GXfDqjWMIakr683nhGyBpXFEmKGu0F+wV86+G1oG2FH0qg4A7d0JgSq6uO
UFFmj+1RXNlggRWpoKHfFaBMZQEtqW4o4KXiNp/IN3UIweflG5d2Iiaoks62ZUZCc1C1+p0t1dG8
pvtSd/RzzdKwkpy8DbsYZj8bk2AExp2ZfqnCnna7pkYT7qDyZo6uvEnGsi1hOWTqrrCltuvFU5dE
C0bFyDvoHnJde9E4P2mB1j29xofLJVily92TfBTzBoXjMiuUxZXWo8Hpy2Uf0kz5ioZGdM5K6XKO
hFlWMlfa8EhKSv+Lti58GU4IGtuJMegMD3NCVGtgyIhG24u8kz0pkdmoG9fouZ2NbSHPFYxlf5of
H7ZIeSp1uaDalUDI0ON/+SgCuWLhGDF8TRS7LkC+Su76ze/YxbVWvjt+c6ze/Nh+sMw/pw+zinMa
T4XlooisbOdyxv9UyUTxx2qpGCksanjIuprSCRfgW6ZwqsGdZgiRISDzeZl5T1rQWWi6fitS7Yt0
tdLCeSLIIudqHPuYvb7CeABDlDQ+voHzd1C2w1o+8I1JUlRK8z1RB5GeFgt2l4VwuMff+mz7sj13
qS18yNDWlrPRW3Gi8h4vlXtvMne0qtRSXjaYrgFsXsqLyF/+n7/etDA+ARR6ekc7eRvUYoXFkJun
uExmLKj0JDZsGtg7HA5go3fyU97i1ylwOQFo5LJHEFfucbUzhJjqT5IxMJFjQnIKyExWkdNngiHj
aiYOmOquopCADPrQ+ujw5JMfZMsolFuuAMNayFACdXQqF8WbUvS8YlHMrmaXew1BEWrkBf9dtnrz
wLRsTSs5+Y3nIQN3IeGZBp940S5RDbcNGj6A3fLZFQwFI4rsvhS1jdqHJ9BpDk2AwTKsDiCOReVM
NcfxsejHXT1zC2BiXb0IaSow3HRYaYQr1dx3/wXU0rE4gsWOgAVlfzJwjiuqLhdPT3dpb19RKTDa
q1wMy71OaQLIm8K1kFjqsySzqSnWjyBd2XdOBLNuRG1t97B3vyqIRBNAQ1ASvkKAZ+N9j2CfwHs7
1Slnn0ZY+N2tDAE44VW1Ib9q1+/Lqj2LZ+7NeKdwV5K43HbAOoW2o77xeKVSqDvegcIKcjvk4Oe0
dFS6XBNWaWyWIHVGXqS4dl8ryK8xGqWV80SWOB8CS3tdHg9gBtQK86ilcQusryovSZz0H+TfoKeC
ZhP4x53KRf2n5d6XIQvaAxvbVqipQWL7c/VUr51/w93ND+acPTPCqYdQbAPt/+hqCAND9JoqKduh
TbMIiNm/MJE5YTwfmGeUHVindah8macIG8XzcoRLB+HEm9SM4dK8r0Tkb7fSWLbwka9c0eL5JicQ
xtG/r1QETGSrzUUqplcp0yLsWBsN0GYoXkPx6uVdYbU7FvImYGrJnafzPvMFhJ0SldJL+7xJH3hG
MhVawYwlbDSLrfpWeCDYR9UCF8rCB456Fret6xJ/NhKEmq0Nn39Feb2aXnfNEz6OwLzbKS0Do9+d
Jmx2nDB9SULUbAEmBQWrDi55GafA2UFCvRdiZ49oWfIe2vFVD10sa/kd8VmnPdONIv7AARn9svct
UnveozFXDgAPkgUw+USycrYg5HpeoKAm5fsahtKDindSnXF5xaEGCvFKQ94u9n7ECxkQJbYlDvwz
9iKFPABjYC4cJ+/2U4jhfzFvqH/WmiOHVkDIDfqsJYf4KpSAf/iCdVzDd8yWiPJJQ64l32fH6MHL
WkCNOgmbUhdazbRzR0Bo+EiOTcyGS82QteO1yYSOg454z7cABGWUn1rO1FDsQ+IsiQP5+Ga3VMY8
bnJnYBpwvR0UrN0XvwSKmcU0HrIg7qE9ck9PgPydZBeQdkVi9NNGPVqRcCBSiaEPgDMGg9hXQEVs
ZsMl9LCNk1x9CBiCmK/ZXMG101Rk1SIu+uQaVpWAdaJIc+eG84NoocNBebjLG6kHe1P6sg16sbaK
L+c0AKaMigePLE9MWWJAPGbneLJ5MN5nnTt154n/AH/aIewT4JfHf6BS61JaBOS9RSTfujkpiJJg
0I9czPHyT6WOUm6XXAtO/0udcHi+ZUfrls/+NlI+aN1w8I6kZd6fWhJzZLrc8OZiasPiktvIlViI
YZPwxTF1byRBHXNwalmZHpXZGx40r92KLuYS7IPfdRzc4ySg4+SbM74DPVuBx2UjLHsC8x0dsFEN
Pc+2HkqaKoE+DqGVNtS+91UWXOLIWpQlSxepgY9UR/CXwzK3hB+1GaQPAIQk9I/6CCnw8UjFy+kD
UdxJcW1q0WW3yQvvnbvweeq28O+Rjd8KWBQtL+zuj/Fd3mrGKhFyK0YQ/C1hAZV5e2Z0ZzXuYoE+
9Tw5OTup/pLsJdYr/EwwlAAjyTQIkTLlpw1gKGIQy9Vf44t0h83mkxPum6PawvfBOVVAVYX4EcKX
qIez/BFLmZEpR1dOFi8GCoqdQgWzwE8h3NUZsDL1cd2adPka1wLP3so279fCTxf9tZzrl4idptSl
ngbq2GUea4Kpg2Hvjhy+W2tpbx5eIUyDamu6EbN604Y0ZcZdLnTZ5WKOA8QYl7Uk7/CLYGcCdeew
zClNS3uGejbyUI5Kz87O/5qf/cTC7Su8tEjFHkcI77tJXs5t+Y8JCN1xzVVv148IsZHUAs6RRlRF
q1BUjUoWJ+3VMuHm6S6lXCzskWK8l1HnDJ4AC6NwlBdoL1rkHKBciZPi+TOJaAmYxnc5RttwRsnX
ORaFQtP0QZ6teNPEDbVMAYLqgaxl6Eqe4pdY9vyTWEgDTkVbr/BKy+SUt9kabllu80RPWVSTEc7S
UnCOh0AYynjp10HRH7WRi+SeV7df/ZgAAnO0ZgRhILSVeEU04XvnPkwOpPbOP7vfT4CJjYqRkwLn
LDrltltvXhuJ42rYnM0J3nqaMkCgNN/PIrzO83w6ELJPq7/Dr+oO8Y4WQtawLpA+Uo+i3aVRSBmc
Pr8RDJIcLB1OjPuUUFezLez0uDqctVSWbiwyfs/60wUGyo/KRc7f1ZiFZmkS++B16YwN1UxITQ+P
GUkv/PCEz9kO+JkOOfXSEAgN3m9K14Krt3uYOv8Xxbi/v3Rzj5rspH7OFg3UoK2c2ebBkI1WQK0N
tq0pLmq6FV/HZ4BC3xTYoqy+fGAwnQzmuTOxuDE+KBM5RWTjEqkcFdBr17c71zqEeJ37/Xuh4DDQ
3IAYP68uqf+ppHLLfAUCVJ4/wHhOEjMDKAIpa0CNX9M9pbidLESukwLZ2pnFLVl4ICE9WhgvUvbI
hEgpP5bdUJVhwJHedKaXytj+9tce5xvWIhjQmbI91B4isM7Mu2lsHWkHHV814tYsNK7SOKCG4oWk
iFB1VOYBEALaOgZbYr6IYRbP+NHv1S7wp9HrRIUhaMO4slu/1dHSwzMgzLZHMbsxk0kB8VWoMU+w
3oHbTxcUsjijxuvJhR/15qQivQoOOohvAU5DSpBQ5OKBzID7YAy8YIPu1cf2WaXqTJX+ai9OOQQb
qpi3WcQBA6gkj047xoMHZx3K8zKHIDPlIQ/ri1oOl4p5pDCgCfUYWVeE8DLqbhX/8fWkU92ugGKe
HwR5YAqrUnqUYMXHxKzR91B5mNrVoLx+t0YorTsOh1C583E1/EhQKyoijj6YA0zxbCDt59bpxv+v
UNsN1yxXRJa1LrIb6D14Vzo65GE95N3pflRXRo3JxsIIXAunSlMdx/T5om3PJNDa4AXOgZNyP+nn
5oA9E6KIer4gOOOfLKpEzAoDmG9D3Mgznx+wHpXbZ0MnX2wNBDLCsAfa7422+7qDFbGj5Ly+Tw3w
JybVvvlMkJWABj/doMwjMJ1uKioy1Syo/AJjgn/7nSxVYfVPuqiBxARPANNyKqWSk9qVyYIxLmt/
q1Kov8ppRBkTvogdGTl6WYASfiAYT/r3pO3tjlQ1HtOooRwR8bBxoMp2wUgKMpIfRL7z3GiKlAsR
Ev/kpxGTqX11JxVH+gPzeqj9EJRk+K1jYThgN9EjVZh82PjALEmWN8quH+ERy0VZYX/4KHPHXeCe
k4N/BANJct5hoZ7swtW3vfXq5e7ja5euRlLrfH/fAOXrAAZYTW/j9BCyBEfK/kLE7Y8BgmsQGqdN
Ltm9gEq75xNjcTIMIMMbuq9+h9/wyqzoCcqVTHhifgwO+oxrw4hwYJ+R5Feio6McmlM8xP9kF8gX
P+r8QSSAcOle5qTclL2q8dy8D1ceazwrQLkWTtsWD2M97PQXIpBLQb1zz53LPtENvilb4a8X2vic
hoszQUSGfCydgQWXK9bNVwNgsYX8GFKxvaFNoLXwBBwkwB6kM0QyR2NEAO5N7TXexq8HZSx7sNR+
lzWJuGyE1nkC34wJYG+Q5PS6yRrABeDIvMm6yloQfAfEOF0IyPsgAylAt5fgHdGFQHo0XfeqUtCS
R2tIMU+wxUhtOw7if9oQEHspsaTxm4pmEx3cjrhJsvRqpVlBvTquw2CTX5FwS7kTRhi0DYDEKKyN
7+tAopXEqBuNohuvnxmtQ/H9+zGkQfTMIY70/meDAui4leaSppfzjBAHLDIoN4tZIgBYRBalutnc
saj47+HQgM/2v4dSiJtuS13+GsTIzJ9GUdgJBCnndHXevya191OOlltITLUsKhyZ78E04FhzPdie
FqT/1ZaRi875DX1hoSKixJj1kkqWbg71IdGBtlQuLuEE5lMv5gOFItQVfqpDRpFoj4oN6WDtmrP/
TEx+Drw+0+EjGUJm0BHszavb5WZ3aQ0jaMOyhCtDQMIHg3xueWswNM9JR05tAH8FK2FUsIv4tJUd
VX7pn8FKI+m8V8v3CwoDWEicE6jIDkB1rmIGgFa6fsybSJM/hs4sl5YwR2lGGQnnnqiryXJJbDb6
R88SlUWic4M+XvT2J0TwOAX8+sV4vdvrvNMGEOJ1jAGZM3+I9yCsByKUnryH6/t4SB/Qtf7XonoU
p6EXzxbZkohGvqJzwnKZm1VXTC5chcgWogu6Gq+K3ehHGXEDAZw6SWrHz4Pt2qgUzy/swUEL9Tba
pjLnucvuNeVPZ8vX7jA2XsOT+W3Dlws+GbXiXgRNF/5tmJSQuvrKYyHY85CkpDzNefzfFzcSNyLe
ydu/NuMVkg7+sKcRxLh4e2lmglZp96dgPqNJrQYpYyrAedOAATW/mdk7xOMD6caPAUMTk0pWZgxG
qmJaM/Fo8BS2ZU/4ueZlkWMx1rIsuE03BMC3EziF4GQV4yrDy2HYG6tlWog5bGfJH0pFsw+snpRr
p9ZlyFaGINtUh9gM3DhQVtx82Z5OimhoLjcyJe6A5+IidBqSfCzvy2vPHwtm50wJP4I38/LDx+cD
Ud/nyCLm6N579B0y6iWqHr/AwcbdsJiLB6eD5dpHKRktq2Jgq8LTtuBrsMESmt4HJXYfFLyB9ZuB
j3tWpQ+YjfJ3dwY3ELqv8u1/04qzgmoE3kzAcM0rkNfXIiSoEnS5UNkASiL1Q1ZtamZJUd1fMct1
pn07jvWwxmMuIwDqMeMP7C2SeCqebxgTHyFyfn16wbNVcFjHo5mFDRsSGtuBiBNjaDKSM1fm5t+7
w2n1luzp+oDskfDyJ4kZn0DE7knSRHp0TmwOOeaauPc4gBF2jvanV01s4WFqX+lEUx9qKaLgrwNF
9RSHByQ4IvTrl2ojAhmshRoeyylT7eSr8kuQGh0tM93Igk5gGjXaqanMyPhssZFa7iVOF/wEDY9q
x0oGliZmJw4awjrJZvC4824u6bukJq0jB9yq1d+IGDK/30ajosDxI2gk+/dgrK4e9fQKu18SKSOq
s8CgfSNBnZT9mCEOyXZ4m80rng/YAVaBXcZXBE35ZlAPJoVceKb2WBLH1cFWIyLfF0RtGIU39DDt
vyyxjYTZ30HlV7YurrnhgtxVCgAxcZGWhLEDpIkRrU3Qm3rCX79FD0DRRKWic3nhTy6HTf6YwcyC
46x4F9lNjB4M+SVYU//5dFJdHX2dq2TTj9l+95nSsOnMWPMZMvQN6Oirn9U1dnPrrJ/h+utaN5NI
Hui7x0gOS9jL48g4ljh5FsTFVHf0uCr/2/PxQWEVeb8p8qVi4dMSmiWWm7n4aeXHsOZtOxXeWRwE
nRmkWNUe4QAN9TId0BDIRW7qkEBl5sJw0BlMN6zO8sLUlHnYJoZOzk745DXrHRlALUGViqko57xg
/89Al8ABnjmI8GRr1V/9N6jJpoGmd+LNXPyUI7ENJqrkiU7/i1A3m2yfiiyTVM7Dm2MdVaEkb34C
fl/GCqSCuIVajy+pJm1WttnudNg8FvUb4QOqd4eWA3QQhwn8VOCtl2VSRlVy5nckb0dvQTp/ZAs4
6kOOD8BcQmecdcazCiaCaALSTJHI7YmlSBpESA+NZkWrftRJEq71k2kXq+ExXU88QRMP7LXRgN5H
7tHZ1vk7cBQiYdQmIRokqxEbI74zVryltFAD2Pe673GflUP5MLNPWXnReOrB34GxnQQXgJ2GMdX/
xmMJT/FHGf69VYsurDyXOct1lZD+7B7Fd5WDM1OBp39sStIY3XAB3FDuuaKB+5SKGVJl/O8UQNAy
hN9EhYr+OKoC/Rd9y/EkGy2rTRacAvyUALvniSXcH/Uzm9D8I3SUYbKrLTtRhCg9JDmh33vIAa7i
PWYrmhHu7WfZuE9N7tUMCiLh6DAPuXsOThrHypAvqc8BodzNWA+fVts5ak8OoBkyL4FX7irSOLNz
b73OTF5XovegNfZ3Du7WW/bb0qhOgYAeVLnPrbOiYzAD3tIC94fcXn8IafcpuY3aFzaZcu2u+vp4
BfSWpwGWRmMdKtpBHHkcrPHrElHOrylRrKLy9WcP4wm2ZkWTR2un2PKZ8J6N+Ayy1p6OMHbDAZVg
DbjghGDgbOQMy1/MtsZ2qiSkWo5GT3qJOAqNRuw6rQQXgHRwsRxSiIAjLZ80qS2CX8QD5E4ZjeoX
bO0CcVEczWqt34vAFM+U2Y3blSupkEXCmseI4THO5NW6PEM12er6JmKgf2xCPVG43R36O7MYm7Vn
8LHoVXUYABNDXKUkB0xHUcH9F6wkzWbqDCfDGB3I9AvdQFdaZT5lAxSoEz65rVr0wW70axpxO6Xt
Df945G6/w6EtreiPzV7eRjGhMDEaXGlQYFpYfJ6JKFmZefwDr7+HYrQWGfr+iWQOvdLvoMbRLsly
chq1cwFaTRpEVZyaQll7ppbNVb+f5oovXiwbXDd+5pNMKZo6KjZbSojppERZGmgJjVDnAVZ/MCPz
3GL2raCtFTMvslrKde9+aw3sWhZB0ZBipsPTWEUrsfugM7CD/Gdlgi2J3brmkdzEXZ2xd2Q+YgZd
7K/rOGknvEBO4iFqwb9Qb9Ku3milpkCiHmwbaEslhrYfzarMM6cmUjUwKFNEIF62GrRu66NbPS7y
B/aCgsKiCV7NB8bkqcr9AYEGrvaAVcM1ePS7br7UBskragfCZ9qU+ShMIH2lQ7NPmYeEn49kfSTC
RIe98iSYbVOrL5xddZ7f++7UzbVJTKhIxXZ+tFTbDrkrC7HKh7SAYvp67QWTZWDTFdL/ohySiqby
odhG192r979YyqBq38t7h6qlRTscsNImUPfjKKuHan4W6RPpdvsnr5iLBMowJPOQHRTzEsqgWtsB
RN1Pox8Patt6XG8Vk4y0q3gJdCx/JhRoc6r5URWsOY65rDLElVJ5/dS3j8CF0FjkS5gzAgn1G9cf
vrZ0K/DQwNztC/VyExcEJ4KddeStiAA2lZWy9FRqS+HH3Ki7U9XNe0YiiYbIgPUpGtRiFg+a44GS
8uzqlQ7aS4XF1KU8TlnkVlz/ejTUzxPC/UwSJ9+O+y4cJQp6WACLQTZ9qj2eoOFLKH1a1vPhf5Gg
8d3AjspOJ+doCRzrWE1NY2wtIBSQz7UBAc3eZjkceWGR9jbc3hAhIhcBqJIPu4jOjeLAmekjlbtH
SHDEq3eo/WG2EnrtkgZfb2WYuZ8VFIsjg1uC30aE8XGO7AH49/6iCrZSo2VHhsfIEaR0+5nOuMMK
0LtLK+WXbZYSNlm8PxyQrASL2P8nrXFLx8b4UimsceBmta1vBmy/bUMKRrVOoxrQW6RQC9zvZlp0
Tltyd7pRPfZUAy4DxsK0ZFUz3YBDqpSFCvQKHtoKk6zuPUWgY+LS9nLcEfLNsp1KROaY3JSmtmhQ
OKIHdITC/8kuM8XiN8IToJb+9lMyjUNGhD8Gm9HXlagZ3BNlI6S1Ld0y0E0tPLiD+VhqfSKipFpk
pHFfDhlpHOyQpUFSad8wKyPhc8iSrt6mrdjeGEJFxM8fftHo7A4aEtF6mUvk3CsGtRRo9ckXYHK9
BWb7TcB6JzbCrJxUQK/TQO/gdB6uqJ3V5HQxD1Dk+9cL5AprDk6wJ7icxdNTKG/aaTfclHQU87iW
JaSqn+9aI+0maY+Vtq5GFmSkpfuTbUiowK7o2mibbBxAu8+HTNN7V9nbULWsCGoFlYWnImFPVKQ7
P7qwea1dIpTxL1qYcGZyHygBqRfoAOb9oJmo7ovSUVZMX8QWO10IRQMqF7iooSzypUaGIEfx0UVN
28qJaIii46P9PgwE1O7DPHsgZ5DVsD5KuDufYlrjv6hxH5KJijpyEVCB0s8lYO3CrOVa4qMbrHUa
MBo7DURIMSXo/yF4L40RYBqM+2c87jNOOW/a/p4m7C5uOQ4CF0ec0niry3xNbdkV9SwR3yRX4Ulk
T+JLeYuaJqOms6lxjIasev57ZWcLiUtF+TGGT4KJgxKxVP6mb8DNFUfSYDvnuan7AAPsFWP68Tcf
DhehuUCJJmq8j04OXAVCdgBREJQM9RF5uoHudB9eUcdeIgq7/jWQsFIksA0I/pQMziBc7myo1kO7
6HI5BAy8l0puadjeWGXWaBxGmPZkCbk3yRbx2YLvSJ2klu6cstBQZ3LGjK0pod/h7SO7Ynwgt995
tJNfIzMK1MFs5NSzfQpqD+IDGD1KrC5yxpB/cmXK7DLwOA2IWIGjIPKhWl3XvkhqN9OnKvgqPAda
y2pLvj9A1CHeNHzKZy833MrHgJfOI2kw7QiQsA1u8UpHoLXGFhQSaS6Khengdr8ZP80pj0/o6jQs
z6JYZkJ8sfS6HFS9/g1IE+H+DsdZg6n+5gkp/d+aTE4FB/8aizisJ/NJWT4mgwpKhGpZgWaDIemq
nEPb1EgIbn99T2t9Fw7LrFVrMZTUF1xgxS2Zrz0h7uw0T6KLMwvtlCkQn3EFA6zEFZVbLcxFxewi
TL2/VDRy9UPwLIuWME6RXmiIVzNEo/E6KlNvC+xkQE4STi/S6oR1z5WO1IHs9W8A/A/gX0JZolww
t7MPv1TWCtmZfzchhEF83e3xfuM8coIgHIusiE3UgnEyiAv9KWpmcHIvOWpiPrPlGbStbG6GM0j0
+wmSaFA2avncFicUpK73H+oSa9CXcZPCQ6KgYg9hYieEUAlmLtlvRInudJBqP0cQvFvFosKuhLrv
TzAT5w6yMRYwDAeuAJPsv6TciDiMBxDYUfsDTS2OCyLuhKJysR/ufUUYzf73J4y3m3tpAG418y94
Pr/urlp5/6l73QWEVmMXXU2QIQ5AuJFR+VKw9hEnjASCuByZRD7tkDaWiCTq7DgNLLmBtGwx4o+u
p9Usnk9KfOfT9ii3eY+eHqCCyFif2NJB4LFD7EwhtxCLBP7U8/A2CeiK3P7UKbN/4SvMb489VREm
ieFxRsMzT97cn/cXOFO2sy7H/6oSiA4H0oChLkaYWCitdYoz6N1LyrSZEu/rzHCpMx11R423JIzi
bICNBNzJfvNkx+TKFnuVYVTsOwX36fMY42sKxeGoEfixM34RTSNTE22axmROUv5pfFAek55GpJvn
AnYNjMhlhVn04SZOz6TKC22D02KD4QIjQsHa7bebTu0xKBZQfZKjKY7mLmvBWarM2tznxxTM+9GW
oIxLyfTnYrtk+8hda9heUYM91CDfSns6t6QnZEEi22+29mOdlAJQR6b+ATszQKyMCKKxhnBv/b0y
z6hck/+J1sGWBINDlOKdG+7PxFlm3hu+7j3nF6Z4Sp9Wa1QwS7Q7cPrVnGHYbGVQbMszREllHugw
jBLFWaayzWgrxNHuxOl1ZfHhziRLfCYYuQyFH+vWmhFLxrMEQ7Kp9VRJgf+gOQmpuEixoaJ8LhO/
lmz46P2Gq94KWfK+PeFCiNjRM9zihW42OgvdRnBWG8/Y5OLosODqnyGmN49wSHK+DauSXRFp2lcL
82Y0AO9UNOj1v04IFOt7VHCtwaQzqAdKqHX7OsUoAJVBvfgOD7ftanHTJc++uIo4sOi9X5X/B3by
SAsCdoVeFyvq4vq1ukdWSprbvQIJlYNSW4ivAm78vwqka1Mwh8ad/r/MDHN+k0xf3iBcvohBDbnw
Iz9ADD6kDEEzZRGnzsGLQaRHRTqmFixcmedNYyZwJT0wXAtmv0h0NcJCamrSLSn3aOU0vGhsmswR
AIH8SeIAC9E2iIbjMvsEh64fbfzAnNCP2bfarWzNGGc1qJWYKFpBRP5aKTIINJDC7J/aBmMjyD+f
+v9G/PHfSIPPiWKRBYzEJId2HMaK4AogJl1VNXkYwJMnIBUyYNV6sODLfToTPdO82rudJZxyyxbo
uV9g2dZyLTwVOGjgRWlz1Q/QWAEgb5Io4dbwcaEZ6KeDg0Yu2XZFLvtRr6w5ewbyOztO2HtvaJsP
EeI5Jh3YEp8x9k/HKUb897+5E9j7wV0M/7hiDj2w1rvQkiXc2NT4XzxPRQSDcT4TybkjxBFmqo8L
xxlKa7zP1Y1gsjm7o4YswW+Po1wguffaaNF1SlCP40go1uLuXwBSUGJZiqSAnFbsVb7lohlOsVZH
+8+MXiH+Y+6yd2TmCwgp2eF/whry8CTlb3kH3RpzupV+aIth914M4HYm83uo6In/mUq7GHPQmytJ
5EnXB86Ou20wFUY+KWk9yKjr0Bz+VOfuliZlrb6MtXya+irIm/AtV5dvCzIhubedIxQTbyrpBGKl
1MeODbFSoVdrF4sYM4bbH+sOlzQ1ITkJRXOctV2+SMpfEvUe9bLCmShFkP+pzZEtDACwPEoQNCYW
uyAnt0Nl9TzaXQGDQwz9O0juPfy7XZWbsZg8TbKqu9SxJrUE104f3U6ufCl/+RC7ityHc5w4f1xc
Pn0E2abDpE8+QIkEukVG4BxEbJjgGeh/e7RGlFzMFn4Kvv3fyVTKeSmiMfB5tdsKbYE8yxJpuEup
HeavP6dRTxGguCAELc/tVTUPQDso7EvhXA91ZIf0qzshXttEZsiz2hEq+IbtQqRhGO7H2DxRQy9n
qlRbDNvkBDUo4n4Y5xqPeN1QunGY/U5EKmtXs9R7bt4FrMdj9k8Makw9MiY8GkcCn7hjyG00yZAs
9S1B0YqJHhQ5FzkaG/dEDg8afXAOBVdRnZACUFCGot87ozv5Oc8Ij0+BQgW0/sNAOA2N8077xwJs
rNYsgib5CK2sRJ3DH/YbV6y5DZ2ykX5TmoARSe2VldVvL0jmtDn8WszE1a8z6pQwB/ZtAx/ixWBy
Q1I2d1cZkyZWCJ5iR0TayFhx0plcK5Qrp2RKaDT8ZNa5wmkehu7dQMzane8EglhyN6GntnGK7BwP
jZJ86GM0yDocK5cz1D+hz1Me7Y35ERlyoP7EWwmhgYssRmXNJjbqgeoOj8bF+0zrkUlHwet1Uqtn
fcT17xlCF2EaAUssuru9PjeGLbjWfLnTQvnTfTb/pbc2f99bxm6Tgeh5mllyFq/PV7ln4W/N8ezp
tGFbgoIII/iZKPVad4oGCeRGwrdKbX+z7lxOSBLgB+vhsqO1keX6+FhbFxjet7Vl9+Sktl79qwWw
5KAtw3RMs3B9/FrQRN3Jv14kiyd6jWzq0+jgfDKByCbmGfUBX0TlvQ6ZUhxmb0h/FzBNe270Vlp/
7q1a96q43I4HCJNY5vlvwtH9A82NITZLQdItpdLnTFgO0R9+1PGycgV7SEHyUhmUd+8XwVvRFYtL
PSSouOK+sdRTB9P8Qs1xVRjaSpcxNvHlBBNE0/NJKiTznWx4P85DXklva7kvVzOVwVFJjfw2yzqU
eT+szUCAR9co4sVeQjGhPsCJOQJuLBULIimoIqkBKuHmEe2vnS2Kax5mSOtqM2QPYi+stg9HAzBu
BYizoDFeE277+GgWvxb+MSQshDkdAzC3Lt3spOb9I0uEgzTGCLUb5kXyzC1xsPU6Ww+dwy/Cicd9
0A73G20euoDFboVNELdtE/LQF5WAA8zbZVF7BOazomkEcwQCJqSZJOCm8g2zJUJ259kMBIzXsvj7
ilhRcbYAFQdP+A2jNEaMmwGZAcGDgEJRg/vxg4ubDUjvoQqWFwlNqMELQRwm1A+fPKfJBtKU29p6
uiGChxuch2O5T9nmqL/cwma5ChVB8j0Tjjg49cGmcic49XmKE0BjFzO6vjYnS3SYDEwyTWec1JR+
xBjdX1uKhP04MMg2w4Frpc0UjkeijFwvOQwVeim0UmEYXlu69bywBVAEkR6zy6fZJts6UZ8KOaRr
+tz82rR4UBaRU6c0nm8qh15nINS/26IcLFGmakyqtzbxhlIyvSEbry/9L3PESkraBN8JvFGyOP39
zeUJC5wHCd6+LwXUdlZfIV94qmOgJhXwCnra4KeZtRK57nmSrZSImJR8Uv/aO/q2IaG0qJwlaHUu
/Iw3d/IPX6BGed8pPhnhAzylec1ytGzRodhXuXUGxT3tkLulVnmQ1nZs5I/Yc3gqtt1y2DpzmpZm
GJrAkMADnOJBIXHbI8fi2YppgMbHcScFpCIUBa8Vb+RQY7UbIOsnXw9TRvKH0022Lf3UUr2T8bPz
16Sf2zrbK9dU94/W1so11H/Qkh/FY2UmbI59Ybw5QhENVV58/K1Ue0maXcDHVspOBaiVb5oH+P4W
LiPh3qXgGD3mLZjNkhVDCbNpu1SQWzO3C8Wbhykp2XvYC7onMVRGrne+brq6Xu9f6+fb8IFyfSta
awCDKXjJoDkrwBMuOYtx9P7u3iMYd05pigvsSFZwyR+daPqnZLQQgOMKSOgHLT/4gmZHVp5vr6/K
rNcpYXH9IU0HSkL6vmCYxTUF74UdMmOFvAhyB3tjHg6OKZsnkIqkV6ouAgPBHdR2MnQlymOp+bA7
imaIk5qzv1RBCCPKOK8znWOJ6SlrNJgz02GR5LkFiwUqyC3Szzmw6nndaaamgISBl0Ma867IkfFh
E5PcDRPP7uW1fcUmWkZa9GOHRi7tHMyVOoLtbGWwYbxXpBEtf5LwRJNw0A6URoB416tuvdWCCHMG
UOwE+6ukQwSGp0RLjEdqXG6T00WQEUEkDJkooHjXjFmXzU1M/l2neNNJc5tHweBKw1zaNh1WeX2B
rZlisSOI/iUPsdOvN7SogozT4wnmNV/evHTMxXFI3vBEYxsyqWZW+WHcQh7Ll0jDqtMVJw+AwlHR
o843BpmgbTTVrMKeXbwnER8Pq+djyYjRqeDbJNGaXhHB6j/eamGpjg4fuXAIRR9mAapbyLV0/JiR
KCkGPBFtnipb4R7uxL2iTGc+SvS++v4IuINzc8GE6WsJDWrZYwC8MhGzh+s9NgrmfmCIpOhS/4Em
L789QkzlVIV920u2Epz5RiK7cFwuOQ1hKAHPsjIc9yTDkYE+FS0h5ZjDNNEZ4mOLfTs9kFYm67I+
J2jdw6HeACsyyVjxkoaqCl0cTT5eOEp77TvOHxcADe+O107Ntj+sqQSoLtRubgm+gFBoNs2zkPZb
7BX5kYJ9RLllyUMY8GeE/mqxf4AOgblv40IxJ2Axr0SF9qszWgw4oyPIbw0FUpYc6HuihVbJG6wv
CgxdeqSNGZ4GyAtu1mTNS35S6LvNtnNq/HbOstO3GLorLhY8o4lgmBUDMU7ePn06E4U0gZlIAvi8
VmQH85MhNWrOXanSEZSX+aYLqz0CajSgKsuU+tHq/76t58j4B3iD1NKjagv1Ox+oXP5i5d1nUZX3
xVCSsqc7mYEceBMeGipH1btFBH6fbXyxdh5ZqFNu+3SvZd66Wy2NLJVh2JWtatVCvueguKfOnAqB
1juAsInYjqLUmoLf1GGETtDRV0AxloFKCivEuRQYMHpxMSCDHzJ14uzjyPOhZXrmQ5fyyQkVsbOX
Jw/Y9g/ytnzONbrI42UBkA+FcwLpQrLQbC4LQ/TCgq+AWqfYRkdWPjnpgwMdKqO5ybg53O/HA54z
MRwmqHSi1Ihm3KSVNxXg7LOsaMSvgeL8Ag5aST+ehY/PldB/uRG/0xmiwNkwFEXfl0ShyMxImfXm
X+i6l/EcS4YXGM14WkcyqVWFH4ZqRe2Jyvb6SamcSm+I+FjwDLeU5kQmYD4YN+ZqXkYCPnL1falb
6OWnMJpsEcKG9sKurDrhpZZ9ebpdpG4vgJNitKTVGQytZWIjv0roF3rlHvKna4/NE9RV2oUJblOw
mPMACOV6u3futaSLNqAxvE97+yzUO74jW88CSxLKTwM+VittvLtYgAbTQdNgcRZJc5TaSGSdudpE
p0y4n3mIaTtbedw6+PBvkJ3DnAuvF9AL39WaGo5eGt1aXdcVD1Eu8OE3WOuM/fXIo+Zs6t5q1xNP
fybDeA1JsOM1WKcwvFpw0cq3WM255PUNNqhtcAMGE605oMZ9f5wM7owshhMdWi7K1WooEn03YPpq
3KZM+xIVDq32JAhNVxTeMvmBmY1Qfa2LuIuz5oHZAfrX/Pp9yltV9Evv/ICsLECsJhhQYsuHfC5o
mIJT89RMgbKUrFrlrjz2ln+K+UEzDW8NU+fpWLGt5GHdHijdHDitvIbsTLsbRyOJGQRxdWQpyD18
aPbeHO6qrym++s935T10eOY+3aZe9+C8HwANuBjhS/eF3p+TZ2gzFhPF3pc+vlq1BHBer3/7ZbMr
C37rjt1t9R0JaysGc7olHcRhWHjd8M/bls/3DNaIXVqRGvETcMqZz+R421GfcExK4hEvuHx83E6t
mLwpnGkW9G7gmh8LcqAsZvFdIiqJFUXdoMjsoFUgZdV60r0sXhF9i4BmyzlACURdhtZZWyc+c/bR
jpoRgBgsRU8mhdmeb3E1oZYPPfIbLerczYoWxAMQZBBYiEu+pp+NkD/H8WbfY3QIULHplDlmj0W2
A69pyq1VhLPY3pLd5injCzOuIYSHoL+eTy5+VPSOfVTU7VQCl/AVbca8FIY8qh/SAs5mPn4optdy
N/KYUUnMAaHH8I9W/R+5d9RlzfKWRmK63AR0J/RR7BqAPXJwm3L3x9zUh+0JtJQkrpPV+ONR4h51
Xoc0Ek5Y08ntaXOHM5ZDM+RhJlSesejLb6I9K8OdtgSsIhgwx3A/vUGIcQUS532kyYgH+1rjr+8V
X4MaO+8Ep51iCAIfVXptL/0OhmsmxGofWCqLr2WKJL0+K8Zb5/IYt5xmj6eStXkgPmkqLRkPHdOX
ZNEtRjuNyxB4mq0xn4lavZOgj/L0zMYotoLyHlfs+LTURdTespBegVw18SZ6NEvRHDtKxj9dLfk3
PYUhQyJIKEoSASorxsxg0jC421o60l778m9MFlm+tZCpMPLq6LjMNFJpPMMob79DHfd5AJLHjIMX
3kK5vbjAHW1LJ3VCgIgXWSjPvmCM4yoXL1Tewit7/xVGxhzVsW6Ved+XJdytsi9N5D0OOf0CT7T9
L0yaerZOzcujkqp2Ejokli1yk+J9j3dR/YjAyH4loXCo3R6PSvtrAC48vVcElHv8KqbpvaM8mCd5
ypwSVI0VxgmmW7mctZXUAApGKX8zo7TYy0BOsIdRYwgFUUI177SDwsNG8Of28YOMT6MNlDvQ6jVE
DfBZC+oLBJuYYMFScsXwmOnzsaRQCvt5t9jEyIM94aZiROMeEqlXdDu2RA0/41K+cAhTOmSdyiPJ
4TI9wDHjdrRVK7Hk2tMcqYv3Ybl43zNT/JvCvIXN3qNW/ligAClL3O3w+hcPbSaKE6YQ12se2NyG
dhPratMfZnSKGmZgIkCe09RtEQt19ercHlyxFte3YLm3vPqTQJbPQjxtnVBgcbFDePVZVpdScaTz
4llOq3j/0t3OY2r5KT1Tzt+abzehzqpDFp3i1kwVHUwIQAr/oyJXoJ43do3YKKCQZfb5WLjxyme1
aNQmv/lqL0jj8vA9BDtfqavb7xMNVkI0mwxOI8cIIkeCXSbG2/MKAWsY10vIe5myUzvsjK7VCkLJ
enGLp0rdhx3W6BQECwARw2Dv7jwGQgD1n1aT21ZMhD+OTwrYlMnZ8hzTGaqxqZmKLP7kkVpwWNgx
6LfJxd3rqzkjDC7QSD82ba4Zw0/FWh+SQVBkIMTbqbv+7r/xMLZ3UJvLzSrWpEr5kP2Q21cQn27w
UTZ/MZ5xGJ92196R50ISXcdG8ckHtbCRXqFFxql5/Cka62orrn7YWoJY8zgwVDalE7LJR5nHAfLv
RoHCuEjLnIxDiViDFD0rm+cvG7gDs8uMSznP/yAqCO7W3l3Zx8k0R3ihLOzE+ZPlMujj9EoLy9jw
UTYCSI8YH2pMkhF/jWwmckkzVxkFaD9WzNonvSfmpU3rbO9poAB8JUXKe4d0NWK3IYv56DpDr3Qg
PveoGzceTGcM7pPo2OGQS7Azug1LB3Zb+xHk6GIDtLc9c3qV9BTvV4x42nrGmnwb26SByGyT0DPu
efkkjw7Cghrxx/PrcmE9j974QUQRb4OgLSeDdDsxIxUkvqxnpNVPJGSKFUFcDXXS0gVNMABb7ssN
eQBu5pIHMJXWyJzi3zFybRojBvwfXpk4b4wsrjGidnRTCJaMLxFhdyOjhtJiCC0zOX1Lnrc2GSnY
IY9sDC06RnWLjFb0PoDge8SIEJpyTWQzjOQPPeAepJQUi5nENu+qI8a5R3wbzWaaMuQK9BE0vXgT
hdEXqOCOpe4KrMi7mj7U1OT1gWGHIo1Wzl2I57zk1mENU2GZAGJEZXUcay96vUwJXmTnkFQD3pAk
91+DwM9EeijaMFet9orcW9+9i6x7plQaD0W762N/P6ARylMFH9fj/0dnwgqdvVtt3sBB+UQewuwB
HGQGGk58UMd0uqDfDNf5N3D2kpUhBwc7TSs0s5i8wUkG+BA81AshyTadAZF1gAHLrqAPcEleMFEO
A893doo8mtYSRNyNRz5wCFdHz4KpFgZnOsJrCVOpqmd65QxT4V/XvV4JxmPkXxMyAwXwm+e5BRDW
80tcRYDy9EGeBdhGbMfdGXEJTjGh5CjJCUm3wQnQEr0L3abwbU5bI9Dvvfcgb1syUKPnTaT5xU+y
US2r92vnQV4u+Ey1Cr8Pg+a1NHdgFxBWRkStEFyBueJuFp+l9OuAQWsV3uiN8XJ5vngGLGsQvcs4
+jmd36ASXY+cfpVoiWFyKHhqLeaGb3AMJKwx932d+IleXs6IxtKM2boYeB0g3+M00ea5ftDt0gEH
BoF7yOWj55W4wyT/HHMezJeHONS2sZF4CFQytc9AAceNcZSnaU/6iLA6IW6TY46i5hHcpQSSp/ya
MwD8KWEmkLfss/S22OvLTN2QDRIiwCPxwserKchzNZfifuBIupyotW8hxJQONeuD0PUUTC50ktlV
ohRH42Fz8kMG+YO1ocJO4kFJ/jD7ejLfa/nrVzRTM9Epiauht5FZYfZy0dNsWoTZVscjlBUs8+yo
1uuQy7Am7ID7sdFDmQEfp44NL+cq9KeiGe+KEharNEhni0uT7I9Rix7EL6Ne/22EXbeAlCIZSulC
6YiqX+9C6iQsgp8zu0vLrnHiivb1zmKMOASm5gANsIDQydd2FC6Ol3LjYa1oE81+2JN30Lx7NvwX
U+L/uPjWxTOE7iLPAwMX4wvLNEuTTSNzKlhcUN6n2U5pOeVIH6GcH1BV5AluEYsgeLRFAHoWftjz
NTQhtXT5RNfkuqunzYYj1QIbmK0Kku/ZU35LNbQzWraghAnj7JIuw0tbOSqI13NYEQRICI8kjbh1
tGpW0+IBAxKQUPaa/Dfcsb3J9HI4IZmX1sa6+Rv69Yj+fBgmQFTQRRmQLjdS7DTk4p15mgG15uSH
C0wA0FcS2Dr3DY4fPvm1ndZ2nUq1hdZgwK0BVV8dhHM2qYe5hOL85fSg7TFiegGHuBuXNdhMHr18
3bWdBwuH0ZC+M+4ZFCSMlnN9ZwkIPqknxhamLurUcYtOebvotKc9dxU77i6xGx30b9NHr1K+yZgx
y2fvJfjjRdwLtxSAvJioyPqDmg2epZq+Ci8WsR/bOwht6FSdfJB9Gr7mfkxTjo2PCb+zZ6qQt4ev
CJa0p+FdBcLRXmQxh0zfboak+fkKHwaAISweV4k8cfVVRKu/B8g/4bceEzoq8wapr3HJ25OrmZPN
cb2S6WdrcBWmDpRu36dMP46CYDg3WLscYZ0qNhooBb2+hjHjkEtulKWqIG2/MN8g8aZNI6lP7k9r
X9jLuFs5sQwSOqAr32ZGrxocawZx7dSvcGqDE0oYi8/V0/QcmW1PKcRo2G1C4hBzz0fvMuXHTZ1Y
QlDMNwfHu9vW2ntwtCJmPlldPiiMaxJ04uN8yBCNRdiHGBicwyvLE98dadjD7jK+uq32EP49nk9O
hB/F4NylkOzKHE5gCjIVoEudQjv6xoVyJTDi7u42IBxV5Ugh8aYW1nEuWt0ye5DWnEskwQSRV4lc
7BVWI6i69vdRZvmITQXpoTGYB1278SX92/ShIt830TO0r5IQ+kvVpvgbtB2VGt+rt0YU41mbZ8KG
czPgr5ZGBWp2/JnFqO0dfWjdgrBKNPgJK4PnxdImaWzNa9+bA2xOhmYjVKHP46q1XBUoyQkgsoBl
kHNJyJh6miR9SbULPcrvKi/ABX7xCHbxya/tkLBAHTazDC+2+Mx7rjSozKE74iWvStX2r8pVdubP
jZS9PEbmGiXL39DVoNuIOn5DP21eL5bmCnd+0WTAeOEgO8gXaQ4BtdXApIv/FAkkx8jqa6pUHUa8
mYl/8hDix677/bGHXfHcoQvlumB6CoB8TdkoHMHXAde+MQnLdutlPhJzn2mKIXgyI+2OS6IQwvaN
/+MNIeqiljteEkHxrY3XsbOn23Kx666N1sdVeV3PRSpjo+YIhdB7vQKV/iaTq+wZ39O55EOA61+w
fbcbEzC2zFH3MZEKuomGQItR5SUgyaYNKLDagiQOpd2GVoFNOvwhNhqOka2ZGg3Cm0GZGM4ULzpQ
LBHSDqQUuMR01jlmOzS+veppE3MNdn/gAti7Ra5X+R3jF2ZyapQHg3fWoPvn1uff9KzbfqbIIx4H
qEcDaxXvrtBjIsMp67wKcXSjBvWTAs2DSO3SNHN/zP2lAcrWnCkkXTAgnNiMwnX72iMqU+Uukkjm
hkoqp7HX97nh0w1yjlqpjTGNcrPHltWce1tolvKyxpcSrL+CfdrJw4b6yZXlIBxysYoani8Fvbz7
pNO5Bkq888IcxDfNsyd62EsKfM635xkBDyJ0DucNUUbWc6iC9Oa/CgPTyuvIRNN/3/Yzxx1228yu
IhtJuuERNsgwVjDRm0clFMzgd6FmPh7jjj6UjoGfwUBZ0r7zSSbY/CBIbGg5cQwBXIJK06MwlrJL
c5Deq5UqURtEVHSYUeGkD83/ugzsOTEcku4fGhIx4SdLjtNotQBeR+dN1E3OKOSoP7JCINBFKjOh
FfxXF0KNLApoTSBDSQTigGrnx6nYdkXtfqY2f4kLAFaRe7aE1YyZYQdGbhnTGlDSh7hN3tqaCk+/
WNer/mZ31wXDkLmqFK9EIv/7BszTgDPHMcQGEEZA1jH+ENEPmUgZLUjHaQFkpa8DJwg7HsgHEU7m
+cC4c8gXBkJa9DYhtj8EcCC7Yf4YTjlz3CguusjH5hBxaidWKAcZUHOJO3e1Hb7I6lTij74TnqzD
C4QE78a5nUkkNk6B0So52wGO8zJjzKESSqsDxi6JOx8dKmobLEpCl7aP6Q1GMfZbF0+8BaVuG9Ee
lwLesHaR6/JXuWXtgd4ya2e6NhIFrZf9jD4LGXKMKrW5r0f9P8B9D2AFLqEkLvljg2ft1Y55ip70
/41t7H519Yub8uYJbgE5b3PstkinSoebLHLcUYbwqRiKtQxOX+34qZel/JKDzxrQ3par/e16KTVF
6IspAyP+i0C23wsUnXhS08OLDM9k4CygQ1hKwnzfTAu+0km43KiiEpy3moHu4q0r35k1Ue+zGL6P
bJOtPqfskuY43qVWyl0tBWFuJ49pVRGXf5nWnat8IRRoFibb9eqQ/bLQc8UqwHTYVU3K5WdUCMba
AAmQkl5RgZuzXjMhDQ11hniqqTqdAo4JWewSkdJIc5Pq+QCIwCQ/zGmcL9pkgUnkbVOceNtFd85/
IVI7VK8dPA59ObuJ3VnmGmYKP8fSRH3jHctjCi4CM9a+cVWFg/WhLBZZVLZYpWLctT5LVdBeGGx9
/6EYzKt6gh1XnjDKmrzUUeW6xPEbA+uZY1YdE9tqPKIx2HH9CdLTUkWtnj+CLhbZT3cgR7+moV6D
/BJGyBtDmSFSWUP1FAL/jDtbt4GzSzTnpP72HvhJMYtvSLwdX8N1YaELbu+47Ilpfn1vAhO2R2+w
sr3YleuXGAa0k4CeGO0gPYRzfLsIQoRHv11NQcak0B5MpdoTwSkB0sWsoXVuVBZXBC8sHbVsydZ4
W3cnUJUl5cXC5E0EcIEL0e7aw2boaXTbvpOJ+yDH76NwSVTVGGgWeTOsM0RO2wWDVNxbbHN508tW
FqB6jtCOg91ivisAwNQ+HLaFYNsC0ZP50elYUzOxgloqKmH+Sr0rKyaeWFkdfj6o+SRr36hOb7Js
XWMzQSJNaHPBZRP+He5kuxIgC5h0Pe2tQBUeFs/VwvPnl4VZ4RS2HUBkVIN1o7OhLZ8p5iCt2Npi
ultstxqhzeumjYnV6BoiJ3Xfg3dfBkeH5HKe+gvOrBiqByHvwfnwl6bMZ8PrpYf2iOl9+gNwyDFl
9DmZfGLL3mpPqqMA8P6ENrxy/hTC8OclIBkUTpngGNKgdSAOOmSyqALb55x2d+c9Ix18VlR8zX3+
KZZ7/T3NOa6zMOEan5qVg9k4l7zR128bZjebx/qJ15weXH9hJz9FC7KK89mH5CvrBOpzm5SqqIIo
d+xt/hL1swUYXAnBA8C+0TvVE6zeKxaDSgxYEJi93wGACEsreczQDHMzKzM5qVnezFVatETByafp
+GJ9zamzggE1M2TeCyPjN18UGJ3V1PMr8rPm/e+lVAM1eWE1/WPH5Nq1gQCxL+PDTB4YrL+oROJK
gAwzwvdvSJ9TncavzYzcSEHllDxcq6T6PgffsuB8ZYnKPKQAxQOGouWlZfBDwKH76JM4ItJ8D/rj
SlqbRaz8AFy1gTmOmeGqRrGR9r4AjKQznF6CCIwMRDF41aLLXiNfNgyxU82IWE4n4UOjgBn9wwtX
YpKwTjmCNvjw8QojZw9W0LLR3deM044cupSnha1kRUtiGAEH6t/mglxR3+0I77h6jgGaqPwuwnFt
lN3LuuUMhjT3cQsQ8QGIUDjFOoobSLCbHBVZHH5kSwkvo4qsjtDd1kUfGOUx/4aaibi+vSu+DJU/
gZAZTE0fPm0CFL7yn4XzOqqojE1Q5TxEx3RYgjt6NbYuHYqTP4JGARqlhN3fiRVtWllu6SvD205o
wI6tXuKUtCjjcYj6uX/z9YdqNI0ZphTtHSu+2pb3h53hz0F/xIojeLXb+SRwHCvuPMP6m7Ng//Oq
jBTm/hM5nuNSLb4cmWvpdDnV1Cz+ezr/kD2j3Lth96En3k4lDtrl7jL+HkDowWfckMm8VsUodYRW
g5kVB3ntA5GmHL56miqpZrVhsT0WP/u2TcYjaOuoECuI7DNjONEmD25peIf4shPftAa4tgv4f0zw
wObjmoPHlzRMLM1Z2aJ3DHgXuXKdgtum4RBN1ncn3+K5ebLaPC6RTFCEY6W5k82bWTQcerljzdNh
/QUdJCDQMXww5dVcm20CcgUPEsMjlVnPNwvA9gCiGi74Fy8MPoCSBAdDQL1tbYKqCtZ+NrH6SBS8
0K26FiAzX6rRPUvESuTlvNt1G9TdMzsE97LN4hU3wblCxb93cC1AiYauuaou2pqJ2l3ywEVC9zoo
sUA3tMyU2RkqQLZlIEGwexbI1x6INAt3TaKZ1tzhCJdTPu+oeD964E0M5fUmOCcqKKSpi0r8rc40
m2CFsfKM5sVxe656TMkxEkGjMcR8x2qzDTa9LM74XxoPfobh4uzlCA/SS8EARsa8kEv+wl5Jl26v
AZOHQx2OubYOb1fSJmEGTDqW+F+ZmeB2Ykbzfz1S/3M85NjT/5tsUXDWG2dzUYjmo+wAK0MDzGi7
2fmTVqnmCG8kUEVRjyJSzbExjsjMUsgJjd04CUxNMUa3DUeZ3AiK36JXKpXkggC9baRXXOQao55F
8AGh5mE1Xpo3QD2fFRq0kV9FcsqVY6GHj7YrDJcWTgl9UTDfQjsm0q3LGIPfK8Dh2+Z+lP9BQqG4
OweWBXra7WpqF0LZaM4vfW4FWD8t4TGHi9My9hmcA0uKHhdB30jIXOU7zGcA/0iGd0jprX2Z+rTe
NpaFwkbRVe7BhEZAi8pu4TTbKKnPHnkaM/+iBO5vBBNXy7Cm39ko0Ed8DEHFcX/E7nU4+OxO5/d8
FMDT20w2VzSEVStp7H30YI2TEcdZ75HQ/p927CfM79aL167Ue7sr8oSoHpxTMkG9C5aXwzezG2is
Etl8O56LJLaZ3hJM4UUB86NMc3e0IaaVIWVb8gxrQRpiy8QEFcZtgE5tj9FmEDwvq7JSqk0SN3+o
NxJbH2kNKXm2Ml5EU9BKS4hxhNE0WuveCSHkoK5itAHHMxu4Jzx375MdKAQ+MjGz4eF3ZLWcr8sa
RFCUsVdIPyzagLCSccJiUy7MXmQ11/ZozrdbfeHBAAPPFuviuyJMmqoI+57ABn5JrDEzGyiux8gk
/gzQingIB5V5pSoKyr7NL6T1tWdSUfbR5Uj/jEZsWTQOUbmkEBHnq/XhCzIh1CRQiI0MSlSLWW5G
ikDjs7rzk7Ym9MxTCKoiJwBo4kmzU+if20EkkV6SVoAove+7V2XtxQ8BTDFz3s5oPjao79J231kW
oTVp10zBHGqRYnh/zp44Is4yEnlLJ64Buw1gHPvCv8T/5CU5LURWzkATnYsoxOE/V5cgwimA3tYl
85ODUp8f0EAP+YJkbGflMoXtEy3h+Igf8LKVVzjRmjp0x+7KxjlftUsGusWIX8WIrkBVH/k9TeZP
YsUWbflYNgIcgEU01abA6IB/N65qW3oviMzQU/Upc9KDF7F1P5v9EkfG4FRfsS2DOkZHtpB4SAXa
R+sd5YNi5MXdScmplbpjZtwJel7G2s9k31fav2KBewN01nIuhT+Y1gQCGrNFckTr0d9OfINnrDkO
socnoQtzDLM8G6I6bdFPtJRZdHq6/RrofmU/qIMHd6AXf0zNU/uUoa6W92WEllmoEJmoYAmqqhwu
T66iata3dCHct4CSJchUm3zw5UqPB3ROAVIihjxoxgMWtZDaOQ2awYu1BUYowDO6FIQnqZXmJotb
+RTcCbYgOWLi76hZCwOuDwlE9gEJMpxW1zVeJQP9ziS2CZXKIB+affuaYJryWrzguNHnl0u11iZc
DexlRpaa2olROSZw0OKCskGA2C6IUWszt9xXp4esFpkf1Me/cxFFDY1Sw53j3vPhGQkc8fLyx6sO
P7oTnuL7ktsluKYLnlWnBMcApydaHollnWqyBcyEncDrHU7RS3nqc5SwMJIL9mssv2gxkHtjsaSB
EWGPfIciaGYL0mEIuBXpwIcxlpPtcH8tgawmFlY7H4UJ0uOn/raslKYix8m/19vW1/HjEghO8C4l
CFeqKl0yQgzlzylZN5vDlklpepX+J8lVLq6y5y0pXlTrvq0yq2oL9G9i0a6xmcSvTuXBXqDduEuE
TIkJAtjVRRDPqg4E1w1GLAhqx+BGrc1wc9nPWxdKQ1egss7hUtZVGZhHH4Kr1E3I331NWlsN2dZV
br3Sg6m11FLx7NuMH3FZvia2KuvNSxJtt2LFHmCiv3mSY1J7QV67yzpPzJqpBdyZqoLJn7WK1ZlR
07eUz1ychCeE0Mgcwu6PitxtlUGMHtE64PUkA0uhUnPeyNr0bPJLDSTzONfNQtX3u/8MBQDXPdNf
WTmosSyo0EnCQw43o08i0QcG/008JSDFIh+x3HwIhpUwPidUQ5ECMOYfu6mQjYNn6P1jtClu49Yo
RB5ZO/NXX8byEim7AGyF2b4jw4n5b3HBSoDSeUmsMDVxtJhnflTagOgnRXP/UyPMGZqjhCt/InhI
FmOGqO9GE5oN7UdAn9md0vZSX2DoIMnTHFJRStXh8flQZ6s4DuXTtnh3zzSejnPwxiif+GCvv/ve
E8/qzOfh4XkiQqFDmWTUANKvLKHytcVdkJhTz8mJ5ejf9joIZiVgXV/er/+ZWy71B83+MU/N69gZ
Ll7kW0cDkiqXP8N5jMn5K9XGILCpJ4E6cOoPd02lUR0ZCj9krDnOB7wLQwc+BXe5HpyB1U5o5pws
CBTkB7Pk35AldMehGd8qHN6UgOAJ6WA1m7uiNt9YyeB7Qu1vCupL7VwXKQ6ZXa1NPRsxbnIO0+r5
qxj+/b2qFYSBz4a0F3CptM8gHHH9DJSvozq5n9T+pkjfrc7dxganA3J4AJOuN2lL44fcSVVz5wGV
32Xm0PWyt0dAf46dyv8E6jzhcmZ0pvX9KfwmFZFhj7BARl5rogaTAW0RKhcT/q2bWfGdbcSFnPBu
7Cy+puTKBnmXLPtJ0rfoxFTuNM9PKlL9kxk92gXvX/dmYDVBLWw7PsG5BVkgNyeVi6v/4CxxmEXw
8Wk53M8Lz0ujrK5rQQmsrCIt3y6IwR5tzEQu+N0OmjCeb/3Q7x/8vTx6rlDM2frMnzwjU93bKgS1
tEcqxOaHTuB6g8hJVPy9I0onj7BM+VLoTRLmWLLFNK+eJ9S6E42tWxNR9pag1V0VVFyaHbjx/0NS
ZHBfJJ+NR+ks5fBkQRqVZ64aMhhlrGd1pgQf9dZADsnoq2Yic03jLcPPHoWhDQjMEs6NVKlnkTa/
/A0N7gidTN0f+Ln4dUcs7L/bDT32sjWEa9hJtUL2cJhAH+rtFhFAKNK7zK1W1pBx5qH6fbVywroi
CfypkQJKaWHNFFyqm22o6wltypjHouzQlA/RCo55NOIGJqrfeFFFZh5RYLZLW0Ae6rpQGGBAC2aY
/DjDla7el5Gr9bDp+hm3IaxqMPoDw9c8FiWpYWbdM6Hy8z+JOYUEIGOCV3/MttEOV4AtJI+kBRBh
EiFnlVGFZ1J37tpH5cT8g/kVI5ww4aEFKG/8px6b1see77jj+6jeA0BsIGb0m/7dp4xNcNGwqjeb
kub/McmwofSB+qLn4wsFqHIUPud9ceBhLVj6EoVf3JMR86rU9AtcT1tbqy0O3tu9RODWWF9ocvlQ
8qwV2/V+KSp1pY+xdL+fFvJATH6vlA7nyrJHOe2IUWZL5oFvKcuCMn/R6hXJfF64X0+iGheotIg5
fBFP/OA1CJ45jekIdfWD9EfQN6BEIuRK4KcO8ERmmvzpsy2EzvHnF2FSNYTW8aFEpPXxrWmU1Wv4
C3Fh9D/F4jbNuJRj3c7c25adPHdUuqIhyomdSlZq1RUpbl3/iMSb9iXkytvAR2hg7nXo+aDfiBnN
R/r2MxG4QDiMcvenTUKUKijv6cGBKqVZtdgCXGViDeS3kx08hVx2iALv3ORVV1Nu0tTgiild1uad
4NlFxXUjrCRAj6f/5i6KKw7fYeGAD22s2QBRC3wxoVeLySQ+h/AhxrdoCYtGoZWHOa6ojxgxEQ4D
9ZT5BFSaxtxvQNQgnBVkO+BMAA/zrQ45Jw371Brdr/LiQp4iae+o9AnKPSsb2PjsmUb9IxuZNUR2
XewYeJgoN/VeVZNIvl1Lg5QKl9Pon6jRGol8kyBiJOHlypmDYLn8oCGcbk04DL98c8Dr0YXeDXUf
T+0RxwenJ2WFXnK+lKGfqmfV+ei2A559Jknu0wxozuLxnxrSDomLWq45hV0CoddRuio6GvCSt2yj
defPib56R6N28mwc/vc6zhgqwVoasPM5UArem0vVRx4UUpaWDQx6UIs5Xn/vr0XiNEOBAaDfnWCm
WrapDqAwnR12YSxRtjRl2VKyeSgjA51/n2qQ61zDIIdioHdWTR0qXQV5VdHuT8lRtD3IXOgO7B1S
lOR5sxUWHPo9IGLzvPqt/Ztli5jf/w4/0+ceBX7xrdP894CMn9p4etIYvQcSxoD92lKjy85Hg19t
/oOHfvxxMclWdhlHut56EOnbhTmGTB9fTZKrPPXW54MAEiM0UguAlLqJP351ZaWG/rtgSSQuQbBO
oAe45shujOxDgz0CUGhte1CkUZpbhGgM+fg8+wjivENjpGLS0R15XWUE9VOkGEY4jZVutLWW6e4d
gjHMY8gJyEaKbKBzmOkmRl0Bdn972uAY9fQoInnJ6AhSbSLRlC8DqsMMa7UgQE2Ns2h7moU0ycga
vjU9Dhgrj5ibqa/AKBFDQUfcLOZfuG7skDQF+dSQN5jYgSPlqTgkQv1tc8qAaXLBEtWL7unSs9qa
letk7nLywivG8xqpZ4PTL4FeW5szLgrwDGbd1Vw65S9wtB6u0VmTmMU+qKRvVdZnLX7hz8/7Z+sp
hbbWEJUKXaL/RuMrly94n0S7U13wt8gsorK/Fw6pus3+cPbqSgnoHxe813RExzlAMBWnkSvqppqS
ZtmV3TlWOnQWbHPxsgLm8Az25Wsk3eai/c2IUJlGIBKHzPQkf9EDHojvCiJiCqGzrFizMAHwLjqB
gAXaFe+5zKrj3NgE0prjyog6Jgi5hjSJTKf5NMK3mCqwYBxOezoz50wMQspl1JL+j+e352Al4wBe
PdZp4O4R4BT1l/scmtffwbIp9vm0uyMvM6kModhTlpfU/jzVwyMXVOi3bTOpErkgFgQC2oTE/rW/
jL2/PO6/j5LeV9j5d4iN6k4oK/nHvLojgNTvWcQ7ECiewUFw6e5eo5yN3YDiF9BaLAulX9D/DLm9
EY+LqAIPVjxbB0AgNiLOcrVomt1bbxKorB1iA+n2QBXIU42L9Ao7FVEV+667dRSN9crbZT/GXN97
DJ51P4L0YVmXnuFBy86APUWq8fjupIVDN3ASzg+6vcVwo0Xi8syvrxwD+WuLftizytL6As8vX9U2
kMt35xgew+Ewy/pPFdYBFvyY4mHS4+w1iOIPsmNS4nRuX+Fe6R5tuO5i+qjOc1siI6aL4QnVdo9w
xqpIXOr2717gJUrimFJmB+wLSBHuRoFvlmUb2z0VbNNGJGDiF8VvO2/jzO/Ma6b9DzmPsaXKbdBQ
FMdX9mFRw2de+xc8aw1uXoPVqRMm+F64NyUTFJkv6oZe9GHWQnwESewJy+z4EDy/1W9Y73+SjqI5
/ea2vVBKT2qkPvZuCYlASmXCA91/G988tcjTovhqEbkW9yWTU+FkAgE88RzMczx5bvWW1RoPn98h
i53U+aF9Gqe9DOyQSIvcNhpdO+mF3cze/qmvXWHVh0fLqOq31FnyX6h+2fYxaJJmZl6kk7qEHEMU
uwpckhqs/9R1f0TesmVHst6JPL47uWZoP2XDEdHIJASySqkQTnzDR0B3OaBCeo9Wux9JYxY0Zn/c
y35Tzrp9LvT5xf4LtQbYJdG+V8uKh3VwVoixS1lIb8bRU5jIQFpuRrgwPJeZbgzvRpbo04XWqVdH
qT2H4H2G8VHD9XXkcI5wKebDDRRq5lpYIVjnXtk/xPgp4qk2FP153ViFwiPFggQMAe95rezaU8d9
y96t8hJ7cE6WC46dyUqy1gp5PalZ7Rw6iRntChlfRypY8ymMylj9XeKpcp4fjBvdHnXNkBMFpYwn
NrIYpfBkVqNPnHT3BUJLUocIs2TQqulDbh7zIsRXUr1Yne9ohTd/cwpNfvuKvB7DxBpQg9GEtHub
z00P5qzGAIg8UEfJ+SO2oK41bC3CzEmFQQOlr4IQnf/xNabd6LM60WCpIRwNNxb2Xw7DQcpRYM8e
LPsgVsu6/pOKoEsVLWJg1ED2Be9cK2Szh4Bo9X5tZO50nsPWxYf6EitBfQHrLGVk4AYvca3yluoh
SNdlDsq1OZcefhkTGaXhU4x/jj+aDumE6m/bi9q+2JP+4hZB22njPVdGAwHUQgzU480czVRccUk2
bQRQpcFmcbno+iEsnRzKgzVb5pHPEHEUJRXrAjAOi2Y43r2jK0uUX7B90R1I0ksC6gYuXZh6GLLN
N4zDf31bIeFLvwWOL8FZmCJYoeZZ0Iz54e1fA7KiM7JKvusMPna1cl/uieWsLdFGeKMds6oHkQ3z
h0c0Ie5Cnn0JXsnuL7KhXFM5R1JQaVzD/mTGyIxLwdKDuQDm6t/DsQXqlpkT++aN7p/p3JxpOdoD
z/Rh046fv+U5PS3/X+UPEGY+ixpoEZdCo45YvFwU5C+A7bJ7dZS1e5k+TmGd3V9cffDCVVc9BNrD
RrT2rxiefohHsm2uPE/ggIhFJfSOuwl9uwdr+/AxNpLteC18cYyf34o6rUvntsaX0mptnTJiNGQP
WfLtS0qHBQuXBJUTO+Li7FXiruDK0JvbbP5G7OjIn76pumPeBmp+OYObzsHbALjXQ5HUNNBkxEhL
AFL4SLBCgXhTdETwao4TJ+syZxwMWTDJh4CXg93+aKnUThGDh3Cbl+XNpUt08XkbCdSNsxilLIV9
SzJQxMBkFgsF+ZgdFvMLpzX/hnMz8IbtrnRZKN2LDTiLlmIrH36Aji6TSIhTHnpqZJBAFdNp76OA
bLY1IhDg0ideoJniG4it0fcQYY5x5toAX/VVKqHlCGXgj+xZ8IA82GfXKphf9h3v3qtm9J8hJ1Sp
x3BvWOqBsjBKo7M+Y9E6h9iLJAZbeVRePSfaf251GU3kK2mH5c3bEi0sr8HTyYCq5G0XFHPvZhsu
rlRitgT4h5gbGK46Tcxy0p5+58Mut6FeNXdYF2TVvf6lMaQWdEgRIqtIB19ICW7GwEkVfC1M4uEF
aeW2hsok7FrGfvi1+F7e7FmW0qiXSuqL+q4i681T/sJuI8WZpI7YRlB+YXz7ntL9mlWlTAvEPaLo
GqnU9/4sn0fF0339VveSjwWtnQOzEQFzDcgWnv7bwtiRs1/hdrKTo1AsxVYBkIU3dHgVqTumm4in
kzQYh+8Xqn6chkCy10fa5Z4EdY4qrbAu0bHNyFDe411QHfRcRM44SztPc8T8W5pGRxAgJEyldn4T
F11yc313ax0F3v57bY8NhBa5hINP+gNWPJccoe1cAq/qzpnYqeQijkeDorBiDwiCrIqztNMMtKEL
j9iwKP2y9BtQAddW2n8aRKEYxtuN6pnI6ljJiweKe9vTOoc4CL79/x0Fp54oaM0sJ+JUf8pVKM2N
YGRdoFFlfRutF2SOsuBokuomksJo8DnlhFQo9o4rFZIFymTpYWBSWX/NCIYHXtYzsJdAr9I08URi
oM/IKJEBUFy6nDZ45+69EBxUsIBJSaqWiTllRVF+YJtYU8DmpEuGYeAwF1H0puRxEIYIEYuXC6O9
tDJ+0SVKB4p4LPRcfonylOfRxrvFH+rD3Jfg4zdmvbSFXBLL5VPJ15VRVU4pyr3kISD6bLejfub7
qhm3ThgOC61CvTCuPRqWFXrmHgDkRroTPANajDvVNIxroTacoJ+Qmou9SKKRHvdeU9m7IEPXTjJl
l3kv1CuYhgt5dfq/8FhgGaHYRi9MzTlAnKOiunmC4dvV/KRcaA2siprFWhBU3sNc/GD0ZFe804Wi
mss7DRHwD0XeQOyeklb9CgAoyWCB9s8UHV+10lkCAsCaQRszd7/s17pUwYF/dioXw2I0BD+XrrFt
e+/03I6lJ5sZ62P8Khen7QR2HHmMLLdNN4GfmedslfKaIjGeNbnFY1G1jZ/mnhBnwns081w8+RWV
IVbLV8xprWOLuB4uRMvxJiVGqWEKS1miu2U+cTPb36uQJkPD4okfBKuHMa0O1OBNaKg9U/4g0Aru
YuUmQuSAFESJ6F36C4U+nHzxNDouM2KsfIH7M+7ueESU6VDQ9zcZNFeWInoMqC5SYqDu/lxr4e+Z
WJQ4do3+gU8f/dVP2Y7izOd4TC3IsSDbrnO246TjZ4tIEOm/CtO2w1cbLdL/Dwnpe6Qi+Vreldwy
XfHBoI3l+VSXy0blpPmtE3YZwsv8d5XfygbzkEu/Nd2CXIjl/QdMmx7UPCBInuk5i4Z/ScefYqMo
1K6fXdOy4xI5CX+IKwF5JxyEoynW2y9nRIUXzKblfdvWPX5c8NNvndlEV23FF5aL9nyIfNArhuu0
c29gxOn0ROxyll8dzB3RMn9RBdKwU5eBZ/yZqwPakRSqeLfPh/r0IvLx1o0pHhgncc9zV44e1hEa
NZU7U+T6KCK5yAUIQR4x4APaA35E3oW5vvVjl/fFQugiItrTLFktdieLmyD9Vkz1en4seloXTQVG
33ZP7MqjwG+UrLMTPzFa5A1fc4lAEV1Yrih8yZSXbKMqWG5ppxTmqX7KSUoMhg2ZrdPoYmIBhT3C
6XgIxEUTw0ZQaCCZEpV82gg2QOQsxkOM1Vf9L2uk+igs1jgiCq++kg1nVtU95rueDJ/1EdCD0TUE
F7LMN9BYU/VeE/ug7pFY+Cn8ww4IiC425Qfr7sFgQrfNdx/Py6gjzMyl+9+qmEbEHLHj+UfMsYKj
fNV1A3dTELP8QRk6s75OFLmDzan5PfVy8gNwm+5WC0F1J8Zv+U6MLkoj9qA+/vQhpxFt5Q4EfVdS
OLTMGYLKeyQtso9oWda2tcXuatG29psqC+ceVEST+93RS1pYcEfMAnnZo/u436VEeVsFyWzYBK7R
Yaf4YvUKbx2ZhufQHWryu0h0KSwgg8VKuOofIrQTlUrARrkryJM+F7y54ZB7gjPzR/g+fgxgYOqK
/7v88aY+2HGXb3/7RWYwgPG9ZBGTvO1Q1GWogIX89AsAWZcXYgSxf7B5Sp1v4Xok2dUUuHH2/sCp
4OWnvfF0h8ot3AA0izlh9zwEq0hJhbRJbGWVapFEOSJ1cKdqm7oTeNhrY+hl4pWGT3n6AIRhiecQ
1s9o1DGzi5YAckmlEQdfDeZozbJxuoCUADTulc2mbc9AI6DbFwjJiDOrWFCsczFSnueBtmxbx3Vl
0MLLv5giFtZfv9UMzWqP/mc2JnrE+I6ojE8LrzG5JhHWXD0rxxxkWTpzcce8rUJQWZEHU5FZZvtk
tPkXGPFGRgSXjG+NFeTdKcj3ksBmSmbMjkgnaCIWpCiZ1ggk858zDcHqxqWFGShbjSkWLJ6qmxhr
/Cto38FeQo1q9wLO3A43Y/cxJnmxGeOK+7/DpRvcpJxQGhBp8CWcK3CAZ5/K3CyrOjgZDBaayyu1
m68/+MDbmi0Bi89wORykdlGn0yfenk1M2EMmjWMhBFWG1AcPPYJ3USMjbyRxUVOlG/6wLyO7wZkK
cHJGeqA8SMZgiNJHjfFUdwZSmUae+viHDefRyuPmKObgE2dgn1spz0ZdUHcc6l6X3WwGtb2yOwPg
H0mSphHpjPxEzkDLWcaf+o7vqY5M93H/kSUfOOtnQmFAuvJPFQn5ypAk0pK+6jDRP2rJxLL62D5U
PwaUzPvAHdNQxsLQIeLGCqir+a7jBt4FzeIaO0ZLsHqWfm2CRh5vUVBqQ7261QFb/HjWbPTJU9Ke
9psPSS5/z2UvJnhBXKOaxm+9z7H+u/7RtFXAu7xDRP9r30NKcvR9u3waFIwwVlkSzEu9F2va4v/o
HX8eqViy0MlQFFDDDKZcstcQHCIamstSYQIYmoZnHjn9Z5sXqFCFgLckziy6Q8lJCSog4KPo58Yq
M9PhjOtcR41/mDGmePGVge7zTPo6EdTvLzYrAyfsuWUYKVPSxF20JPuabdVJpzXg8eCpcQn7LQ8R
ZkvLVV5TI7qcn/JfcQ6lfx3+qQPkLH2opf6tofuZuAO8kzxBEM83XG4PpnpBrr9XEDN0HO3FXKhL
ZHSXJc02IlcSE73ZZ5GVCCJLbUSIoHALogZ+nUGGDXFymNfFWVCXgseRDGaP2XMyTkmfKPvIDc+A
ME3BBCDc2oPyBHbd3e2IqGZefKIDvzbocmbVL/mF3kNLDLY+Ahm/vvm/JTGpUWo7iQZmADtpqbYC
s6oUZYGm49TlZ3FLc9hLhL+OuhFV3Ta2mOvVx5OYyCIdE0JhkFba5o3veS02Lr8Qt47NKFsItumF
11f5+hd+kzg64bRqaSUu2W0WOFCOLJxIM7yneM/hl/bvEwWgRHoTiGmN8K5RVwn0DmlyrWPgWY9T
cCIKLN9cI3wA7tPxf3oeXrBJR6aJSKOgTLdHRkUu4v2POf5vM7pGCT2/g+lA+jtTk87pIQ/Vt7Fz
3ttNPxmZRLd/JlgYMtOgPbLYKgDe/zR9uDWYzzmaE/57i5hHv6AQU03IY7V9tM48kyFm2mLvJ7J6
zDsp6ObyAWOmIdhCdq1/q6Eh7FZLX2y+4Nlp3BDObuaBQ70/REygGa4MJKIOPEY09axkg/xuQ5YM
3ffaSzpoD9Zyr2vf3Dm+XTWh39AA1ydNvmgNjGSkcshdqepdswZGingzkY7IyEdBI5XjOCnx2XoV
F31HGLMCGf7L9k/ZT1XdAmqZVk7H+IkQf83teYsvpjZao9KDdCjYiJ4YCmaK4sntk66VcuGzVH6b
TwwVY22F0lFMGzhCszTNEic9Z9YCrMl409kohnrZEnP5m1rv/6ct/OzzDspwYbqjKhyoSr7nB4dk
d4rXMDS6sVPyWBx28dpJTdKBxRAvbNhw912r1JdRNovP1avBYyoM58Um3sagozA12lN2ZklY/gAF
K7EOkL3+1as+VsSq0BaMwTCQsjoBzzCHyLmeQsFZTVZM8KmywIgPdwQPYx7xCt28NfhoS+rXwJXF
EFp/3395w6q4bnJFN8inNGIVicZOqmq+bhGbq9rNeKyIRGpqp91qVXrk8Y03a8tm9P09CmzqNNIT
gl3UKAGnQ+xnrN/zIvs4S7JouFc1DulPS1xONCWM0e51rbnjVc4AGJjLg8asCuDJuxVy3dy+OFTG
kZ0r1SS8GK9GtUyY8XiS33BJEMHtAC0IYrvKpHg4wHF+0vMfM8slmzm/rv+/N8JOhAATQktAFv3M
vZnFB5TwCLHIm9LWDOCUMCOCEbes38SUmrN9gqWbYP94JB7prsfFKK1KI9hTUvCelBRx2q9DPMs6
KKUGvV0w7kYXwp+YJXQuBL9GcfAhW1ql1oZOsimLc3nOMZ1XbH2dWWxN7uhuqdImDm59sQocZ2w6
/9QnHL7CepZsvIq8lZGgJOLZygmLQ2wedZskuphFEIBHQVKtyhOUVo3FmAtq9pXrQZGb25zJ8RVI
tDajxreCw83HboAmExILcU2J9ibc4vQKBzmmKfbWiU2bnLs8GI3hokMe3Hhc3/9q8lsEmbdLyAWJ
7oQxhpZxPbLSWjWCDMqbS72FHchUd7UWO4uOTbTiBRrvfu6m4RXls5boVTd2WIcvmL64OC+WahuJ
lT8DfxTbsMHVQVDblpDeQo8aKweTKiZPSFS8a9qkqkG6cRmymyYqN0ntw0Z5gyyQQ6Bmz+sengLD
2JGk+qUzcKnA6ZBxXAc3YRE0qBpaWSC1q7QWaSwIxl1Jl4GYCxoiHFiZq0/0cY5/h6T8PXNoQT/i
4H23JPpsl4Ns+OSS9DYHcU8yMNpTPa5DHvTkdb6ju4Y/kpF/ju8fh7s4x/tdQ5/zUxbOBfp4OmSq
8Wrd3nfKDnmxxpm9JL543WAaJUvv/l0j/TqbaFA1oM7dGQR30G5ijZn7+S6m/f+BfBYVrdIErDJ6
pmmUndal67sOiX2TFJsCoeg1ju5+LHdaYPG2f520Mtd3ktCL8h3FUcdARlDXi6/xUGMBEbgW1GCs
LrSjNvru/H7Rhx0AOZbC+WW7WmSl7N8r8cKRhAQqgk/z6KkiJCRIYgYXWJ8dwnmPsqI73VMyPVHs
DOReQ67TFJtMt6/ss0huVkv363WQRBou0tRLpDIpdzC0AilzE5f/RlPG6Whw8cUCzqBik9NLHpj4
aB/Zq5TR2mPa6AMqHp6+47cuThYwHNhNZV5W9q2sv1McwxFQqUkzTxOryXGP4VKNTH1EAi4Xfm1i
R8IXCuuqOQrz8NeUtvnTaSlEyGrRc7yG1Im0WZ0dsyVap1qpZmHigW/JSGDYa4cfo3vyF87Nezo+
tTnpqdG6wGhumpIKd77amaY23VOo77v9jDP12rlIHWuJL8pX9t6BmVzVpDrX3Fb6sX9ULzZc1I/L
/Dlu+Yx149MD19WgyeVEMHwjjwu8teTe+w5pAQb6hnjmKYUK737lxEen+HTFOMsPKyY3/2CsAEOS
o9uq8kjozxLwNfWgWBbLL8j2n9Iwfh5Mbl1u7V9rQM26R7WFdXzQ/hwA8wuLL5SIBkIog4u32lbF
DT8p/nuoK4dm1hhX0asrvYlZ1O6aY02nQJ4rU3Mv7qSHuYauBIWoc5YMCZPSqglqH8pKMTRcdjp5
EYAhouJ6mmhX+LjUt7fUiE3zBCWILauv0qUCfj0ELWfXZhQp5zFFXdzj+DlYDY3f7+zndv5SXza+
MitBoWhkm1E3ISlv2mswZtMe8JUtezHS1gfKmQbW/UlSqhNf6J6IR9ckksyNQeWCBt3i8ikSbuJA
AUB+05h4cVPq+J2bCNY0hUOQaqzFfYRgYT0tgWXVKcTi/8rODs8HrlPQep8um/NzfznBUX6s0ePm
4Q+VyqahzJ/fUBtm7kXdXnNd7pK7v7XDszg3yPOF4I8IpGpv2yc/jPxf6DvSUHAoYtR5zqIa2Za/
/gnM5iBN4u0mSqXPwCp/aRVMnZCo+Sxw0uGt2mzTWTBOIb4srfEZVOcqog6ZOfWbMQAXryiiK1Eb
UZWQGO3Z9L4g25ZQzgUyGpqdEIujKc0zB8FSOcmVPXcr2yTKBjPniwG1JeswqHRhGmsVxdrqFJvf
CptLESlDiplrao+SAJYyAKp2REn4ROMUKJes7j8eMJmYZw8mEGO7R6F4hfMc7HitKLjfFuOHMIN0
GG50pg4Zbaj6J5414x1GO6wZ4w+hOh6PbwUDWlhJUY4dJnxgLlznw39QIZ9JpB9fIBcyC2RhkrCu
jMYakBkf28XLCe9aIZlIDv2IhdYvXrtj+5+b7tnhusBe8lgHJaNi9PN9J38PJzZlW/bYfj2vMZ/+
UYdkyhjHCV8fyx9TPigeA0gAFMnkjgxiVwL3JHBpehjvtQjK7b4g3594uQ9TZ4Y1F6N56CkX6DxY
a6CrNFmsut/lrhP8jwmZSxHA+7m/Jxp/HXegRDypWYn9kJNTTpoMMEXTeUXAfoaXTMNDamF6lSwh
b1bkBRyJzp886OCQuEYJ9Aey2qrsEdL0bKzGuxmCGudmK8SoDkJ8Ha9LpqHndXSXE9RDNyE4Fcwp
IZFuzkhwuJ8N+uO/MRcP2eOBKncIFIV+eJWwZnVN3DnoHyoD2PcCmmZ0pq1AvSiDFeJvjhr7Xuy9
lSbN9pux/cbi+SC5cJb0Etf287D8QR5wzyI9xKDqK3qEUyMXA+93hdKHYoO+MVNxn2lTlMRScBHQ
f3MOQthn1C5tu10/BPx7rtRf55Dpk9ioPFXsC2qiuTXxguHTZOlRoA+9HYOYsZFt3JByprGAPiBk
/fo9AaMxybFHWIbQViWglTXBuKvqq0QfcG8DzX3lt4lTRwAqMBP62y05Cxh9S4/Q+6AVW0X5oQF/
D+yjvm3E1RKVPOGHjBU5YmtdMwpqCEKxTzyPTGlFXM4Lqb3EDACevusJeBIEqHTXZ+d+9eAng4U9
ak7Se63JIBQOGgGu7fVuICR0hZOuVq4e/itGwWs3krSGlNUjtzTgWU1Z8tQ6RzH5siar3BiTVtVM
3TpnKIehoYQqQtQFFb17MRSibgkpF1QOb8Li+TE1YwJ6Q6ioejOIPztofStRgfEY0/K4oMc0KYM2
w2LvB7hK6Mp03K6//VdYF+WFebIkPPHEQ1m7626X74rz1hHQBR0l8eeRijlE2FETL69A/mToPA3i
jb5C2gyFiYrAAc+8NoD/iSMA+zb9IAWTFfawdrLfUrqPblGkJNKzdHJGDrCBhmuMdKGJJVZPXfk/
/HtZEr+Aj5JBK51YkzOgYhLfqePQgEdnMUoVdlMX13tMOHP4DMt5tExA/RtduXVQmQOty0g2qEtZ
LR3ySdGvjQtwC3vd70TWKfOveXpG/IcbpZaETBEYaKfPDL6wmhCzctXeWn6TqjVerOvduhz5B7Vi
bGSqDK5cYcutAUOIwXiUjm3QaIMHxaCLlEo4GJv/GAn0NfqJuJp8qP1s3sRUB7yJYp3s16++lNbx
foN6TJFEgVHMIOi419dxducamPp9wLd7+U+rvRnl2vRD1ciUxc3W5qFUbv8WBTgfeVuYV1ya0vvC
yY3mNn8s9d3w1pxrRIUXEzO5LbKXN1dCsDwUmg0lE6XOshxyKQO+zr+8Sq9xGF9Vuqx8Z1d9Ma1p
1pnikfZDYQMc3Nc/cPHprldKfHE8ZZJemUwJfYkRlP3baEjhTDsivdRIm4lXcCbRbmzLQhlkh721
vvSa/rCPim05lgjsKHULY8iHbsltahyAnBtdMHbm/06BSH7ZJ2+U/p1h9kOP5GuvdQeH7/LhVWyY
3AxYh/N0lqnbXk2qC5ZUZWGGk6zO3G2xTxVuPvTrQQee5eeT/oB/LY9Tt6WO3d5NkOxL0izvEKIp
bclGZaG4YFnHZv7KZisduhB5tz338UYynTqfNKgVKMvdkCV0OvpfZpIRRQ/Wybmtu6IbONCSoEzE
RQmmao1TWm0DYopBTQjO5zqgb74BSTKhIYg5Eyuq2MR5sRN5lnzZSNQ9uNIuTCt/DToQ9AaB6H0G
XDnMlm0m54Y/++oxsi6ZTI5s7lOy6VoP34QoQZTNZhEGIAGPVVdp7EnaM0rB+3KGwawaoyh76OKl
WZb14FuOe+r8chcX0jhoqqNu23Lw7jPlRzlEgVm+ypH1ErXBDQIAdGvdlduDa4rwrlR5tYSZGhh0
4SzQbx8s0mfNbmwB8ZPk00pydd65GxUgFc9/NS/RgZhZD5wyERjI3SvB5pkmoN47gcEYRKojcrtR
hx2KWP/Fi/nHGP22ikETK9B/49sh1ceiR4YadxOyBo1WlsmjS+qeADPSb2UpNhB6QCMNo6c9W+lF
g+7gvuFcPYx2bsj4/aYHY5HiCK/RqmxlZoGT5ZarVVuMZnkDo+pekG2haPLr6mgwx4cHHj/VhOl9
H4r/u1N4VUI7WHF5FUPdtFxPk8R0mXl9fdOp0jwOlzCwwn9OTTLtBr5LU9Lm7MHzuOLLwNBfE93D
r1T2r5F0HJG1rB01aj1W4CX66jVijEIkiSmUuxaN8/izoHVHIbEFFxPYxrLHoKR8Z71LIIFWC8pO
9LriYBAaODVo7Ubn13vWeiHtxn1uITtPJalSQB+lvlBZZ9yfPY9s4UIQ42wHR2uWKbn+p1kY6yEL
8Kujv+FwPRWshODDcQgsP1QNWO1mBw9LDPmd+s1AxAneIXa27Y5k99X+DbxziQc9zb6NHKctYjos
hFyOhDMbf1Qg9sdAX1lkKRD2f7616emINXsxpB5wr/mAfHLAlikE0Jr1qq6uMsSuqWnE5IXhMwdc
HubemOi4UEUFNQ6jWOuoBHqXghBMB4fTIoJwp8erdPYVSfU40J4bR8y4AG2CKmWVa8ZfpTa2JmN4
su/yvTlMXDq17hY6R3ub7wplvLjX9UYHHNDxMKeJBV0ja5MMkwg3MER6OA7dzOEfXtLsPDRSkRKt
kxNgnpSivlN0yEaqjcpDPnbxcrvieAYjE4szB0bwfg3iJbu6GLELE/JqvmIK4v6D/So0JsSFi3Fa
s1JxGME5EZUt9HPcY+mOJg0NEljV/SJptV03TILdTjnKkToiv47mV7zft0+nyk/C6MAWDXCd9Lxw
aNcRaieB1im9D7dF8SdrkeZoft7OrEqjV3xj8dEaE1cB49TnYSb4+wM8eBEtEgjhRZvbhp0xdJLv
XyeCwIGZ5J7ombUrtYG2iGGI/COhqNCsAALnDvb5FmYiTuiX/m3UltOP8UqCan1qHbT1T4XR0Zsm
mAUcC+38/n+ghKxfPNu+vhJwyN0rLd0cOFdROeHTp3+mGmFriybIvK+7lgEqdJ/KJ1bMvqnbKBmX
7T8lfUv1OB84+RQXxpBrvUFTEpIfcYphQUpCD3Ol4hvS0bvSkCGaWDetbJv5qAGNJ+PyKxZtiNdL
6E8WX/xkPyMgqm2IJt6nSQnCQXlt7aH3AIbdKC2Y1nueYRpKCzMwtLiccR6M/hOPdPlBVMzGZNFs
9no1nSA7mPtN/EIxN2613Dz0rW7KknbFQarbNkfTvNHrQ3w22artex/OFGS1QEInojg5ZekosBQR
4rUHQZpRiBrdk0StkEIB4GOUStk+3I7LgRvCTk9jRWZrj6q45juJiJR5zC5KBg1KfNlUDxAgSFYJ
Mt/diArX7XBWfMiNvdN7FF00Eli/Hff2HuY3hyqXx3OiqM5JTH2yN5fGZXk7XzWk2Slx6/kGBDYh
fF4/RX5BhBI+1knXqUJVpfFSNHwD6SEocyXGVSwjlgA2DdEiEF8JSR7/nf7vNsFzVpZpuoJLrnbk
K0jfXcDE238DB1GB4FXHlIdirhhmUDM0qc5a0/IydoemaQQj9ICzictGWw7GaBtQhVIAvL3wQhN/
71bvNkNh2EKwcDt23ECAJNoFg2QNwpojU+QCLcgLyPRc3zeCzIiZgUqr8AtkDF/MD4PZRuk5OUKM
z1+RcNUPLHoaIGdjqmA66s1x1sreTX7krq/HzrQ9ab3lKOBBjsGmurVi2aRopjBXLe6kH890IYN/
LbEVrQvBzOFACjyiwDq80Kaf+uVk8AoaKmNKJ3RxyPe9N0S44D55rqmE20BXtMcAdQyxabPOGpSs
or+AM4mH2s5sseGUg+k0qKMOQ3BA+01ozvn6OR5uk0lUYqRoSrgdBUDkGgYMlFhVOrw1JtajnZ1x
QgS1l8ZSKMWbSuOGLKhSjRmuitv0aVz5FOCAeKPhr7EWsAro2tfJHd7Z9og9fFiuakbTtjL3h0dO
0casob/TwlvOGK5OBCy2u3fua1fpViJjmLr5mEZlah4oux80x8JBlb8SHy6Ep7oZCCgulxrGZGBq
CofXpkhUMtjRbzASREZ/ETrlnIPW1QuxGHrBZJaNqyfeADvQoEsworJg8wPNA30zWIRxC7NgGWiy
koNR3Zja3eN7NXaoBbW+tgtsuxW+jgBTJYaSwSQYw3zU7y5nP7842EROi0R9gS/eOpOnTR5fwpMW
BN20wirFAHNtp1R2nThEwtFFNKyABaRevqaYQE4HfZ/CRFnj9tuAyJopoziLvmvdnZap3p+gzGh6
QVj4veXR8t30OY7Fr3oYOot64yUDJJv+CjE8PRuRN4pu4nZ/xp9pCjDVLcrpZh+haV745sqvebBC
lgl66yOfmJJ9TTmy4FR3tWUVzSNGt0K8Vpro1DdWbp9htyGiepaprdLzHJ/lorDI9TKVqlrGDETo
q0g48sta14HhwfIFoXyyrl8pbsO93hamj8PGnab/3udsI6Uc+ihBtImfmmBC9KzH3VjxACYaXw2K
CHZBhR+K6/xb+K6JwP//57XxwOHeQNrK/4SU+0UbuKKkuZW9cdE3cx2xK140WJ1fhWAKNGHyO3Ve
iWHCK7j2iI4/zEY+q/FG4ULQaeWHVvNKXOQ26nTXIpStqHM2m+Mq7xHYaE0+OIoWzy+zO3OJPqKp
+iqSVqEr0igld3OjInRUTctlu/DX+K605eC2CdrhIaXIGhOwRvt/0HBuobmr+chmnK444jPLV2rU
te0jGw7CdgkPCq7Ritg1smbHUEwvyAwzYgs4JzS8m0z9FalCh6TmF2r0LemArV6JFHHKdsytaxVF
Hp3yF8mse5YRpRnE8MMKlyqqF3W9nqMn148CpToVpEiboZZw04CKAOFhZ6Rbywy2FkiWfJxnScmk
UYbMiXIX2mkxQZIVZmQRpgTpvO1h+JGve6r24yKLxtZquIS8DaqoVgFqNzULbfh3tV/pgYXlYOnu
USb7XEe98IUmo6EPxPMF3s2YfprutH1TVLg+kbVELqKMsmsOhk6tHI5FP7fZlwEkzb9czMZUi2Gp
5Mioc6cY3yoD1iEy3dVZDS1yKTbOrcgSQuaZ5XYtW66jR9ooL5p5qlExjaU5p5Tl9sTfY9UPfKMl
Za0vP7mQ/ooQ25j4M+1Ytz+T1V9PW1m5XnbeebQREvuOoGSKnbP4rWzyJ0JkbQ2EC1leOMadtzbZ
UdyUVzqRMalgrl1aC2amU/rDMv3lhRsJBzjFv2n+8eT+VYVRm6Z68z5kPC4HASk8Cax1AJhTs9h+
o8aD6V/gOe2pqkkfoqOvxw+C4sTym8nDUNQXH8b/wTifh5VGsgfMfNUHThxaIqMGlAVM5RUFR7Qb
umbDR3vquQjCLpL30NF7slj8mOz367ebQg/Dd3AchKMT3+qkVCReDkcqaML4hrLFct5H02U4OuSX
+kHSzZ/S0lJ6fwtG40tMXCM79RFcXQsoY1/1s3B5VmbzTxfwHzUNFvEOE/lI2Xqj/eX2yKDzFJ24
8fyK3MAuHQ8t1An1J7nnSh4MXO/e9h1WH0NRIh3WwP94FbgCm4hgcxVJ6P4DgXiPodbaBZe7yzvA
WT+se7Mwhk60dAQ00bdjnM0OMD+Fx2trPsZR8RRtmOnA7grqJtNZQBG9NDkpZBRbgg7odpqU2P+8
POlkbp3Lto3DnFnPFAxfIzfj29o5c9DmGwPSrCKe0/O3XK9XftrqbXD/OTkvE56s/BpGNbmabDtQ
06iaiBtvMGwZ8xLQ1BY03Ctf6kOFMeCkRY/Vwo967uvwgOYjK7lE8LOAp6Lc6+reekIIpEwedHfC
5Q8Zb2wTH1zAQjrNquH3D36kbTO7QG1Zf6cCPOjNJanoTihFs68BUDSrbuhfjaE6Dc+bG0/GuVo9
hGVtsYDxJFN8xKzaO/G8gaK8homriUrCjYefLtrxIGpKghLzKaEb4GNu5DFNZ0XrIJlfqMcVNgG2
keOiXJK8pwpCkTklDn5PCHj/p8R8lDMt8R+AF5SyDEEFOXlSRy7WguUtObRSLRtwpBS0xkivYIW7
yr1w8gdue/RwSbsXvPzZphvBVJX2rqEPVeMg4aTEAQWsHXKhu9Dm++0UiAilBGpz0xBQo+J0/Uzo
jg0C53L4to2Ir3eZGwS6AHldESa8/2SSPBTTL2XUYVplNnaV5j4DAUf3OOE5EPrvm6VF2jvMHc+o
xPby6tQrOunt0+fCfeksmwlXIfgmGaavpfOhjgGUwMswuChWGerBl1DzD50S+YLW+wgOvPSKIS/T
bbPz3x0S/cn8ZBd/zl7NH1Yyvo7QzsFSZyXpOU+O1cHzTgWcszqDO3xj9xt8v7OwT/mevM2G1JMy
VyOjyvcPa3JDCU0lsAyUYV5c6dKVnpTlvNnZw5CuTcwPvYjMtxrEhWzfaeL5n4JlHQqdtJCt606X
hypDaEcymf7NiLi1yRbWoLoTz1pqMNpIByCMJ17kLWwBlm6Kp9ZGmptHsUhiNTqviz+y7f1I0nlH
9N/7H3lqGVNRoNrvuRlfy2O5+sLa+9Tp1N7BS+P4QeHXl1PKOYAJXBj7Lcr14dbWCvpgAcJkEZyG
ZtXZNG4cMCkKutAsYNMWfkp7jQwqvzrDAfZzQe2R3g4hycSqYqWGORObtXwcI/+0UYj5LsGMKx0g
hDrQyYVTvAAOYY/sUTf0NJJbl9fHnncGD+4LREvterFazEBPpz24ZdgCnDtKoE3pG/UfSo9gJZwv
jPhq7JAFT4ycRtp/ZMSp2IZp0GsYuU2IZAnzCJiR6tEYz866K130HCj19fwV58pw92oH2VWOk/a0
MK345d1JBTWLm6dggin/w3F4l6Ehk2lP8thb2TW38regwkce01TWqlgcv9PC4rjKkH4jjEpE3zom
ScF46eW9zTpQ00YaY2C9/8jhvm53Q2NRtp54XhpfL6ZGL9FW8BVlDnWsdXJShO9+4J+9Hto5G/P0
cqeFGrTO6pXHD4vKYPYzuJZ/3fwkz3iTTLh9Q5pojsmU/NPG4TXMkVP29r+6aoKZLGY6YkAHnkKE
vgXnwKeCrphXTQunNFpokgO+AqKD7Q5M7Yxdj9tBbBK6qRWThCb7AIklgPMNELpisK05ejZ7SmLr
aF13K3HAy2NqIbS4pIqZyjFDvbktmiVl/9UgHYy0eIutDqGGG8nU1N/mdWFXVdOJw/8s75Ne0wq2
JIl8tmSuWRO0lsbDRdJGfsb5+EzSwefSNfxNvRHrYTSZnYnM+0c/bIQO1z3qhcgSGgBQ0JgaoBpp
EIEm4XmHJaobjJZih55S4fYHGO5h/2KP/bWoDlbqHEjruE7fA1Ny/uZUdTxiO1CBLgfHN0qMzElB
Guyk6jXdhA9dhY/4D6lVEB0+P2kRpuY5yheruYqrgEOYZL27ocOsF12TF2M6GuQXKnFgorbXggJH
grrs5SuGUsURn+p3/KTOAYeunUxSZV3nvtR3JW5oosQv5i+Tf3PxMBlehuTR8XFIp8/wDhRV1Chy
zUBvMmQPUcY3zYSxxVWa2Hv2YKZ0WLiRhcqKnaEC7EDZXgMNPmgxxZR7aGVUVIW7JN8O+aDtFKVJ
OZzgasGFL7Jz1hBqEMGd/Tj9EvQ1zcVWxldxJ39vDROi0+SMfLoieS655ud6qCNlCx1EXJEBfEcs
EpH0sl+NBMDNabQmCPhobiqmeab13AmYWEXmKbOYc9qWWJ3/pmrf7tlaeEc1V4I8ITavpxjPuNjC
/kLt3y7dgydWV/t7DiPSk5v6LOl6Y5YHzQEzSXaUJrK0k/5NA/d8N8hvgFNbgvZ4gdbOWpvr1dK3
CNUzULqU9WDFF9X5wxQtqZJdaB9wwi/robkkiPtkTWJvs9Qtdnz+TNpU5vRevLNTBWub1TfaAVBn
k5oQNgAQj0H5T/4yfGnUrTtL79femDy/e8S902AatbNz0MiTq3BpZlVlH97CwqBZdlFTBBltxIt0
a2f489i4+I/Ip07lBKDd0W8KstFCLiUw8/p+eLzitKMjtLwHRw/JMn6X17Pn4P2y7N9wUwrlPXHI
foKqz27U9UffG2oENUBroAkP9w2LeFHy1W8vDEGuRDX4fmgAicNovwHYfX+bfVnMyKa+mMPG5T8W
up1mVG2EPLj956ahDkTUEQ6QBFAlZWCYmliaXz1rq76zz77WQntjUv3b7OX4KycKEEXdcX3f4d/H
ay/vxAWSOmYfxfKBym/Os8f4Ch8XYSTbPnaUvCGAUXwTDnSGifjoZAG1h65IQvnHl3S+D6ifrcyJ
iyEUx9I/bqqPgpsLMtqcHOym4DrU8Z975vYopuFaZeiy65KKrGSczDK7RaaJhFIUkp2A4eg6WahA
0b2RSM5PanRgfOb047ej9qCEjqnPKjvkH/IWv3hMWpf1m13qecxkpk1RFbiQFCv6RuKK/7kHqeKh
0oZ/bsSWz530D4Gcu0Evva9g+nDy52ecS46laBjeFDHWwuQlZoxNdsY7hCh7hDvrhS+qzCWxtre5
9PlzwV2Fmi/J/uH0haxVOT3+PxgKUmrRza3ZMnZDlkRaoz/YwQfidVZQFu3BJBdu93XC6k7AZ2y6
uoVaUMM/momqDEp/OLwMooPTqX4I3NtcIlZqbnu5d8Jml4cllKrkOTOUuZGyr29iFOYnk9s98fiS
hvSVtm3BPeKFKb6ycUc+PGv0BXB09Cywec0eN50LiDZkSUJAufmXU3HDiAjfDAJC+AGujU6nzX53
WfUQIdbHMzwBTiLlOutPpo5iLpOLLFAPvIkDmaxWAVJW4rT/1cC5xatXUBkUPu6t4a8wqJYrt/qS
WPE/rpDfz/Dx5PWALfVC23KWDzN03uw2YmHRYS44WWrYxQc9uhE/mxQKVGbfHwzcaAt21meNX6C7
Oae5kbpGTIxtENZQr5jIoIdOCcoyjHKyWysvWzYNP+3LyZJS2Jhip1qn7rIkR4Ljvo8ZPgRP4dNc
1q+5tzsP2+MGSXId3ioaheB4Sxy/AAtMw4FAneel/dscbDEvqVfKanRXmcbu/QjApDEHVftLh215
QVVYaFtyfWfsx12Xs6z36A2rFQzwdL6v4O7MbScPLubBtpSo9PK7NO+MPq17+7pYPTkn5BUDompb
9wHzOdtriLtniWF0jPbdUdYcO/3nRZvJz6YMTWYjS3xav3qGLy531vo8D4RCrWqSlgA/hzrmiEL2
gelKpz/hf6KKMR5QD3yeGc+HyoNgHRAZaPqrBA7Qrin1Kf6gUx2NLUPHIBTDZi/DjPDIjlD/bhrL
NDNHevckdwy+oweiLG0y514alv//ShjMZlP0KAyfKDdUyQlBOCux43DuIwBc8ZZp5U8HDe50RyR8
/VC0OCECN8Cf7tFR5RZ5rpJHQ295rRRQBZ3n538QpAzUgyH6b3WhugqGQt9LvR6O32z1hfb8UKw8
hiiynut+2IYnfPPtG9xU0AaqCDrBVY5SZdwTU7g0bPwLSeTix2vmuYihVd0+dHyfgLhYvgWA4+b5
AGToYVHzejmMH9e3TJ8SfwzwtU6iaCgDbEK25tr6eTZqcAljA3qiTX2XxNSqTuK6etDEkBFdqhzv
pfLN0mNFJNQCtvIjvj3bBReWa43QiyooyU95XacJLcw1wW6JuDLcyOuubGVbU+KD75T4RGgKRDGH
/uXYquClA0j+duo0YriAcwrEKp/EpAJmYcDS+4LEK6Ericaxx6W9MOKhYU1xbs0weoQzPw1jThfB
/x0FAI0uP6+ckxkxAIE9iwsIzZXaVe7zXKRwEo4GcCKsf3CItidrW8z3l1x0hL5cN+HDE41WOcJv
s4x8AHpX+8wZNc26o+7OundMtlzXbDGIdDKoUh3h6Y+q1GzUfCd/wbDcq9Bdeuo1XqkH8ac0UC4a
WR8emVGOsEGN3GY8waG0F2B1YHORnNAJVtGodRp2vAjqaPsemGHDulc7ii6Zp6g+mWidfZ4CSQgn
ELLbw/iLZCGtlAqLRueqz834rgphONxMLQXViwrHMpRMWEcenxouEEG7WMsyZzeS9vYzBXlB4XcA
ekILLo/V4yhjA+ELkMgnKky5NyitbifMxtL5B7KBuHq8cYe1ksIkyuYiScdaVqaalsIvWHgXkDkl
qPvMjSV3Ok77bWm22uOAsCEVVYMxVEzRjXFBPwmQDmW8A5Kiu/PtsZl2m9LI/eZWzSFvFJce9DQS
I+7G8yAgt9620g2IGjN0Cx0XZI7SG2jFC7rU/B16jHuYgSClyStqZyoyQKCWzsefYHt9GSOKYiNQ
pkV9WqxHFsfqhcyzcTkBn9jsChp+LCr66or3Oz1pJfsX7WlkqRP46VfZnSRVugf/0oWsWf7wqpVR
72VuOS4kdTrw0MTmgPY641qEDgkjTTpQh+slvh7+vTYbhs1qbeMmf6yNgHq+VJqCGJoBCIORSbWM
XP5lcMgDd8cZ4YJmeTjkDHDukDh/8df0Q85ctFT5A+greugaW/rkVpTyJ6VCuiPss0s8GdKtbEBX
ZO7qa08Rt948VvRjTqXnIScfs0awdyQGJBWJeUKxeYXNwnWW7EqknVO/jrlXdGSxAAR2AS5PFWIw
GXpnW+0pTjqxmrTEsWs/9ZX7iHtv1wrnLTFBkEftQzWnsnatgZuim1Zr99XfjLCNRNwZLBZXnVNy
23U2s4N0+aKubuQyUWRTukiExWudc1EhYG0PEN+UDNTNSSNhmR6D92YNKzgBjsO7dhyirzxrsaaK
UkuAc4hnY6cVeku0zGXCGnN865zX5cuyfCmpDq74wN6ZYfZ/oBkLSxgzEtfZPMTlKvlhUcMfP544
rvi3siCr3Btqf/OMGvmCUb3ywcCHt73CVWPSJrmMmBjrFjmfCZwYUVuB2LycexJ8kWBlpOHIFGft
e6S/HwxYtvTVSN0VFBXi8w02jlkgao5lc7EDpg1kv++kwc/ESEV2F5mkVyxO1Sv/rqZHMtxWYTy7
qrQERQHYSYH+Qrxnp0KSq9ybjwLSqIPhTLPK15KydE3xKLNG3c/I3sXPuS0PMEKqXbvpriDC9Ws3
IUOC4+Vq/9HFAsNcPlanO1S/7HWq76FcbPosWCynl2URI8WjxkBtbvNUqpvg6VNTmYSOMe72A3qR
b71pkzIYRXP9SLmjaDNBavUeGNDXZd/CeBFaMS4FDL8gg/AF5sBeokNeCEjtW008Ed6Fln/Ehynr
G7mPAwhszyXY6qaSbtIGNSsZp3udRY8c3cZi4iNk/9jb983aeDjPTeevISNjfHRfCXkgxankpKMt
BDNin4wbj6QkqAcx9FVzU2NUhRhI+RWc4PQcGsrRqt42t70qtatXnL8M4cA2wsvYWrtiE5h3965y
KZZNICAIc+Yubmol5Ll3Sj+cr/lMiXPThrrT4OxauS7oUjqzRSPgPeYyaT/LcDXgDnKmgt9A12oW
VaQqU3W4Xh4n7MSnNGNILPw+dV6cJbkWv3WYqAky8EhNi7uA0MqhSXydp68iz5H/cyW21CvKUaR6
yyE9F5HrerH6nl9LhhBJ1LdVqzQdfoJ0PTMNznKVXmXj6Y2PBNj5s8beXicJEC3W2WLB1UJwoZ+N
obYpY2nzOo4q6nZEx2sT1tSoO/Cs7QjvBvA2G85mqdZhkQcKUBRRRuRGaB4WKpC90w8jteqMEwee
DwxJNFsIgK3K4/DYhii8mb6UXCdWrhuClIXNaCV8uyCLNqWLXO8tesZKPQjN6QEChineqs8pP21g
AyfVvRMM4tcK5fDPXdm85UAYh8nZFFnxZDByc7uj8k5ocf5Eha50KUT4zTPHMj5Qe4LhChCNyqUO
oBGB0C92EQGRTI87YZSN7KhQrdXRSMr+aXuna/5iJZL3FTN4IiDDtwHWGnyT4JFiubTpxFgJbeom
scLLWquBAwOKHnoWVppO9+/ttjaY1so/Q4sNU9lMJscqp3o7p9SdAxiQcm+2B1HACEadxPV+zlEb
BNpkNU89VojBLBRpz7F255DF0fWkLJwB+9+Nb30VqjTLQukDNLemWocztyUHWAoxbbA+34WoDA0O
Hj53gqm2ZEjO7qDUA2Lo9i2bvWemvbhPTO8LRLMNWH+To8GTgQv3NEFxq6mJtWnJU1ixkk5K5VLP
z1P4qydmF9LPOBs0L/KLsGV1qYjX5pJFSufqCm0ibkQrqTN7TA9xd0t55u/rayWrhmqalL/kVUxb
bwvXgy4ntb0FsnSxGJY4grmcyKU85wwGtzSErBs/vmhlQKRgZj7pVKiNHP90in5krKTNOmiVNWI3
TiEQxrWc98IIzvcinOMtKjMFlp6iemF5sm/pdNjhxEHHidHs0bg2+/EwrLuEcn/t5DoMJjLOEg0l
IZiWHaMBVH9lGmy7Xpa+ma0l0W+VWh9Mei1c6p3Q9uBUi/DuS5W0gzuXwJy6Leel3Mv9lOeB54BN
1z2C3rcUjL52n6rSGsTj8lbVGvySBVfqsRsaufMCtaxIWhWNOSkGXulWScL/RKTL0pA37qXes3Vz
F0F7Pz7MYZek7dJ/+BykuVQj/O+7TNFKw1XXcYgwYxb/8tlgW1dx3ub2BtrXXk2D+8YRNq/NKFWc
1e3HjeX1xhhat6ED3FvGXqqLf/guM3MTswC+EpCTlckDMByNyQXnjJZ4O+U2Px0D8iH9XLJlEfH0
vPbaBLUXeAdbBYTQCeAFHa8F4OE/TdkxAq12NZerucua2dAEh2/H9vuZ+3umLPAZbCUBLTMKl6+y
5SzuKZEb2m/lWgrcrqUILnh6GPl1B2LUOF79l6N1q1gcmlejUQsS0ZYmCBRFZbWQtyIAMLJ0wMtg
vEOg/RjUle6pjgdeSAXyEWQknCYOtu8cdP6hdeH5HZUwupWULvkCEXmQlzPORA3TPhIBJWrd6Esa
DrXRNztXDKw1q9+sbdirobiHJfLCyVhCwoxkXIOnyyS48eji8goF8MrEztRhJgqzsMVJ3XXWTQcI
oG6Ws9XfQ7hSNqMgMN0NimNO6B3h0psHEa+gyAmx5yKY/w14icVlOObhfad3NoFvyWPZEjZUEQzN
5ngpSPEdF/JV3q5asvNrPNYbP42H3+FKYrYJu4Pb+Rmzb6VZBRg6Fi7DfH6/v8cTeI021TyaT6J5
srGoD5hjYf29UvdjprVeMz5w474T0bfNVJTCYKU2L5PIGUzpWk1ZIfPoIsYcNeaJllzXARvpe3WL
W1c+R2tqCG/W/c7PTZf5QaJ3xtYujhXC4RPghs7/v4UY/xZiuxux3rUNxvaaAnTLBgyp8iFHcbdT
C0tkkULp7LjeJYIhDsqi+uA3tQ7q7bsNrl95DRlsA/sn28fR5OlC37CGKmsdJ94AkbI6Jc9ItOa3
TB3Y/PSis/2znwfsNjY2oBZXNRCdXE9OhS4RNQmACpMACk0Bp8pc1ySaX63Nnx3La3VkgC/MsEGz
vSWJCUPpDbTzPf9rRz3aO8g3uyfGuRMrl8llZquo4mXNspjEfoVg1dKkv0Y5Byhgd5ani00NxVrr
pnAWk0RrxvqGXzIFRUwgvqIVQyxwiol+IXqkrjHk5vDxoWSQiSAhpY32M1jw+QQDD+OaaQ1zV/jT
Mg/MtEZnEf0YHVEfEL6VroMUmydigWPBli7E5E+bZyveyfOfb8eRPQq+IaA2SAJSo8v0cRuc6NZl
ZLxPeYBnit2phWwpbyEBvfb0XtC9x8/qrZGkJj9iPi1aNzlDxQco73YwLC2pSueCa03ke0YyxfAf
jzhB86+55fD2btBjEEmACY1GKrilpr4ejpxdI5rHwSKUEeGiaaHONyaVDOo74NPJfUa8ldMP3+fY
9QtWLHKPng5ptR6E2d4ET2nH1eeMxdDON67JCRE+RZy6uTSjELUPpi3WxQnDA7mwtRUqvclQwPZ4
B4GjduFGzwBvCNAsEb8/54khi/VKjkFzzoqSPAhthRJFby6dRZo0fUFpeysDxuvzdtB2wnBN+dH4
F9ZBHS4trvMXkklJdUwURCaKVh2F3zKXwVWjwOGjbYExd2AWW0laUuztTz3S+Zqg6VenGUDEVp0/
P/D3TxvxAByGUbBPpRBMQpzJ8IHQPMNI3qAp/ixM7Q0yOwBqRqX+oR8p/0jAxn83aI23gar5yWe5
NKqgFq5QP07u1wvGPsA/dScLReAd4C6JxfGu3q9jIi4vI2bQZ8TNxoEyOzWOy2CUxbYyb204C212
clhylA85aX6dH0jkZfnRW6gObKCWOMBhMqFm1WEXlFrIwMMNNCNCvfg+UtSGS4EYmIn+zpyavZkw
K/T5eA91kvA7EF6yseJ92c+NFKr/pODd4HwS/32Y3OEQwB8VaSHByyG1y7yA/dG45hbPigLGKU4P
kpVLrDLhYmVW0+AtK+FxJR67CSjcSZIuh5EtEZZPCPfuRgP3yFwNa/2U6GIS8Mp2F/JghYFRx/H7
EzYoQ5YVPrKb9IOWZlXTUzjZ29Dr4ggb+j2Cz8q6El0InfkYTd9Jz0WCu+J5pKIIJ6wI5Ja+y/2e
VQ7HPo9Z9PfIrTHs99LP6u8Tg6F+FI14ffwc7U4O0uR5tGY3eB9I3vDO/sfB4tx2Yd09yrBTbXaA
AwMcZPjOIrQjo33ZbF19fcCIQ5ecML9OYYVjNCvOL4lzXe6srDDeWwHqzYFXq9U7iu8Y9XzKnIUb
s6xMiWTHMg3Ch0iIkX51VTRJoL9k0A+7yN+XHxLgdlZoRZQKbV1+kVTMvB6KtKto/yOuPt1ATeRq
Vbr+Ftsj4TawQzK6fcI7MjDB5XwqjPFyyXcQ4Nycm9PfbBRgbooWi82OYkADw1uOdrBSnAcr8jVu
qmpyk+Ex5o2Y26bSo9kdgK7ar7X7c1n1fC1/IKEj+yDQwj7oDbJ72WiPHhsYlTgCczXlrcU9QfAA
Oh1QI8tQUA37Tao2Pdk4mM4aXTvSJ7HoFirtYnw3lO9jxFWFDsn57LGFcM2A1yeZI2lia5Y9dMPx
vArtnHcRsANt3qDQ6GJcMebyMNEhed1e9bl+Ojva6oZVa8cpZ5+raNBetpwGtyjxXVdcbLs89zic
C4/HNUhgVRyWrSdpSLpQyrRgZyHXqjDikgIMf178qnMRuXL05CeqC2DHIHKuZ4UXnZ9mJqXFP9+U
GEPHIwcQ84oPyBJEnMiV++eXlAhhK9Fq8Ee0otqlmO/PCNiHK/bhDkW285VMtUlL7WCYAT8Idly4
EP+7ZdEsFqn+Kk9nI7DCF92X0z2EInML1+MCKI3A2vTZG29zBo7IO2ABv+2rq4SXlNKoOLblf4/I
vLxx+yu2wnFM75fFGXKPDpeouR4DkwqNvDBMcDYL57wABT5rmdc/cBuliLUhm2LZuAinnz8RPQZi
BWBNjyL3uKUF2dGlwGd0gtHrwXziujLWjcP84Zih4AioUi32TUbF6qTpGhjGpA2wdxcKFcrQWCC5
vJt5p1t8aHFdr4pl7UZjY/HU0M2sGzt5Tmb2M/5payFliZTyv6I0KR1qTws490JU23JebkQcSJ7X
rbUP8Zmq8JZT0ZFIEsa6OtR+o6V0JFGNij1giaYgqnLAYKqho0dGy7GBAMHR3297NvaQVaTfSMyl
+PJjQvkvwdGaSF63axkmeP97zYHnyhmbCm+dy1ORgszpRUwOY79NNtVyUKUX8TNADvIG1hLM4rmU
XqHMEm+HHHIoG1Nx/Pbu6TwCQuVMr0Okma7LbTXwRn+adRC7WCbq7IBz1Z161GKe9L7fa7FyRnAN
t7c9XZYgqb82Glv8nYoDrpnrIeSS8hZnxVUCSWanag0a/bMLfS3nyoKwSe10HnXqt9zsd7t8lbUf
QI+T9MRPaZqFoC1F7R9gJjnhMLG159dv7XgPPqSCDqqGL8G65Y7rm70n60rb6FdKFmQoB6Et/aKr
yv3v8aNByFm5lTFSwnHSyRmJ/Vpz0MJU/hgc+gZzb+RfFwTxR9KiR9BGqy7wwyVR7i4Gu9W/Qfw4
/6JwSDDcP4eLCJ1Do75qymEtqW3QRcDhh3kzMLH5NipIRH7ROP7XnoB8WEEtq/DZ/hR5PxAFQrYo
ZN+IR8yj26QlnFETszF2f+RlKwHQvW43FlwN3T9Aq2N/kGAT5S7EXxhDCcy3Ys5uDnpjZuK6gux6
ZJsBwmeS4Pn+2b2oef5frGAO75xjlNXbM9wuqdXluxdX8h9c6mkVieWEGUIA/50NhPLm2255Cp4a
ZDRtV+s8b69htVAYjpHAJ3f3fSE0h+qI6VgL2H99lh2hgQzpIaK2dc+mwWVhOTxsqoW0WrR6Tozj
Qzih/9cmmp+U8sfrAi2oKkc9B8RH0nT0vw993SwKiirYRcBBYv4Mwa7Odj+nAo7TEz2I9zJaCM9X
Ge6bQcvODLnrgH/NGKi5Sm1JPBcAdX/6bFtyKGwKxdZq0wEl5HY7OQGW1HP/gdjtq1HalfQtieZp
VyTv/ggcR5/6F98djY2tnZhWptg5MN0ZJ5AcJTENLZ7RNWEssbQ7Ix+UvbDOkkJ7uDPLCRMdCQ8a
q4GaVlb2304u+OcRL7BZCtWo2P7NkEfJvcZKPwCcFGp0Etv56vnx3KvO8E1Od1vqEzkDHdwRQ5Tv
DDXH5r+eF48di8WFKa9vk2odIy8OQJyb1fu7O4AFcyzmbKEgbTqZ+4nI8nfGiTPRUFA96unUC1yB
Fd40+StUjsE6FpEFhbXEezSRz1O2pMxwbppltiuK0MpFk2mpDmUJbn9ZZi4V+2RSVkNN4OoPnozl
A97cIA+Tx/kA7ozEgVFAjut2mWq9ksSltP/FlFG8nHz0iNTJaPeM1us71VDzQAlzwEEUUZqU/Z0M
LKTBSHCUtwg+Wy6/plC8RkZ0zmKkjJz03mWLAe7WVd9JMFDiaNh1KuJ49/U1aT/xHLPDy26cVX5k
+A+N1P6rJphiTP5PFIBQ67EaYH4R5yaoIf+Wzy++chJWKfvtqgiqSQdbO+SIFCAZOGbvCfAeSTd+
iV8XphNcTL1LAXfon55IeF8onFj0iE9G8Jsw8s0hcxMrCQXL1o+FqgfC2Y7cdo0jtbvGuCdeHxn5
DsMLx1OJEQpRxFEq6hNDhKVP6LtPvmif26EL3o9tHnLKOf0LTsiOUR5zEKdEbJvFEpH6pJCF9qay
2tqNy2RN5c3IVPwHmpC2XFZ/qQ6Y5NeoHaKs/0zlrLMCRH20ZbiIMS3lefeM2WmVlkmEVnlel8sf
FLLRz5OwWEodnK4HIwLHnU50U4VGVNcR0ZZ7e021C0DFAdPnTZeZdjgN1mBxJmCQweFD0TBTZUJU
UEqW3lGjZlZXQJxMcDZ3y6jhTpOa2PibyeC3FRLPO6aI2rvnGs+zZNO48pTNlcMUnmMhq1Ae2Z+4
WyTwR5E4e/it7zFgCwfd3ZeODuCNwjx+oLsWYHPuwwVJwnoSV6YwMkO2uDClEHvmRLzwO7+aM0Kf
SbEAnNnhJCVscmrJqt/r7k7TW5W7tYaEPG6oUYwRNxtcJhyh3O9UaS/ui2qAjMiaANygunxtC2O8
KmZXTk6SOFST3Ckelh5xhZnhhznXMRyb1tMsxY1ZB8KbZkwAV9Vm1+p4HrrU7szxDfmrbFe4IbB1
jWa71WB8Vhr2/9kgC7+I6x3TAX9S0xZ9+Xrk1Dr+AtiDlltu6G83JpSd9PKxAHMkWGnbqU3KuvY2
cI7qQ/aF7eDalovXt7FItQ53yfkXxC/6fqtkjy0rt5XQL/ceFJ6WrpbPipg4BaV6Xhm7vXvlAZ4d
zKUSHbL5DT+0kuvS5K5SH/N4UJL4qXcLypQ2kSx0cw0g89HqQcgLxy/9uLDv8bQ5uqYqY0MYIjDp
4my9sxAZtauM2vNUUFpMXe2JTDuBDN0FmABqvdH5+5pZ/JW+6OxW1LI1IK+ySdF3NF7Qpis/r/SK
1KuRX0ocXO86MWYZ003HvegVOu9kpRA4lrcZiU/8bmaaZuF7JMLZ554biC430e53itJe0qynP1OR
WvigCeNC9QYLe0mwKUkfTySRA6o2c5adh/4LhA6kadnaT18PiHW1+LbD2Y4Exc6q+Bq1Naau1nky
sVe+KSbdHISWv1HufnWGxrfyZMQ8YFAYulaBoAJVe5KBsZZc09O2WdSXUrDRtyujifUhobB6rtEM
uih0ZeGvuU81Jeg3GdC9YhvRQId269bEtDxgrh4QTKQVElH9c9eA9jyH+JQieb9ueOdEdoTCtfwd
SYxD0HtdmonAQg+6KATCMlrmsOSDKUs3reU7HJx1zdaP6eGoGZzqu+kqE1nGqvXsUAhFS1HQVCwM
JA7Apjm4efNr8GCG+OJD4Bx+wEp5kXW6xsIn+ZbmnKVdQiAQo1xw/GW40/Bo98lxIIqt4mAS0KBW
cXARwfXyYjOScx3lSANQV2+AW1JxbGqWd1j4t2tgljPhckSi7FHt+0waXEDV2Q/qT32UY5236HVz
jxgobZIvktwteSgdPd48RG6tCt/wZA8bSTVwNbQK79uJZ/pG7Fi0jF45T1w3Y7hcduRwt0SXD2fU
01+hZtde20TIzzHY0v7wa3gktu6hSR/BYRCwjuOeG/AL+15wkIO+ZA9FLfwa9oqN3geTiIRvhtyo
W2msI9igHW/znQfqVT1+R9JkvhWVzoZfnmjDkHHcj9dDKn/oxdSSqeivnA09RzS8zVh2Y2zO4NUV
EKOoxQURYUarmuwtvN9hZvoc5AutSLICsvXM5Cfp1ZU7N0pxcoUOemwHkibu1fLps1tdCrYJT2ZQ
gGSYd2vcLXpb+tnuYVktSxGPpMmDHBKQgu9hlimp02fGhgdAQ3HobCkcVUJLNStSQDe0tiPEv/5W
yUBY3pcXQZG6LL/hgjFCHzldwWszO6XTS90eVMzwp2bUdZPMd517pDxZO3k1c7BT2jEJxEypwSsq
dzBA6jv6Yp2yZuADmu8S4kqpMM96ho470ltS2TigR99Bg83ZplUjrqQq+Fw74vYffQZGfTy7uieC
ZEkhOmimtm6jlIRZfLM+1kOTQAYTClNZzCdyVMyJE08XhN2/cAUmeD+tZpVwet1LNM8rxfTMJBWv
wIqxOVjkYfglEftm8bj5KPus9FHybAwu0nsgipjd+mR2xUpR07ZYFdmwOOtdfIvDbkCQ+r+5DIPC
ytTkE6E+hXhMow5FgOj4hZWI17DoQD6PlJOlZ2zKldfli/4meulTERdLgObFc5PogQy+EnjuA8Oz
LrdkzPstX1y+id2a/eaXXDCee1ezSvyTZTvaUE2ejVfC/Bu7JlixeWUZbrcTEX2PtIjg+Qly+ydL
P+2o000C+HPm52rCfCwAu63tYdH8jPp0Dh58p+CxAcEIP4hdR2d5yaqQYswndKuYwmAl7lQoBrIF
pBKGGZgBg3ZAaPgg8lUXSiI60e7/PoJOegkm0pLqU/pTOhvlVzw+ISuKy52TphNkVmEQozyMbwXl
ciNGMbwV9MOw/TZe6NmjhiKRyhjK6LZevYxhH6bCWtNSOMiMIDLeiWdYn/TC25EWfY0Bmbl+2jEC
EDE/GQf2DqEQa2RR2irCGDW4VOI9NVFhSr8PbLU8FHHPpd+HzHFyH9mcVMkd8OYt58m9J1nARCmL
etUuHUTkgPuuy6F8i/u22jFhm8SJoDjTY0tRwWbPqOcIm80K2NvuNY3x+bC3UIYwJrP66gAQ6cmC
nVZUv2Z95Lw0OhfMk/bG4RZppjuD/wI426OFOGRiKP9EhpFfr+tYgU+NeZi66Faxynl/ExWdlFNF
2vkroZGneeG3mG0LHjgtQz/DEktmQLvmrEku2Bmt2jfBwfRTXxUtD3ZrN6AlKTKIftvwdsG/8wSo
LPMM3+sNMIxwKXhzSnHkBF6kk9TMXqlmnitROeYlh8Tg4lxSyBgbR/bQ1Ique3uzzbA0uOTV1dcA
EC2JpAkoPoks+9xaA7ADEk5h9SxawPA9aPb9avZE7HuFNG2VaS5Wb/i4bgST837v0C6RUKTp1Aef
nte//R4MLqbl3xWnpRhquSfT3mI+vN1C6vWmuN4zBeJPEk1wGTRgTR07gnFynkiQoUaBieh3XZRD
3UEv9ClIKVGujRmrOrcIUlFuWw0qkNg1AWUUGPLAXoAfPZ1molCSFmT7AIdY73mLaxZSW28yfebJ
QuRSrzlJpfBPrsc9r8tSDj5yAzUrZoiVmU9HZ2mFop0JjkfbvFOZ5f2qznLWs9JrSQR2AifnLEWS
/a2BeBrkGQPvb06hRNk3p2nrQpzIn6M4ac8dcdOw8ls+UP8OxgXG/roJnmYa1wOK39s2ArdoA1Td
nSIZIObBHcWPmM0tIJFwS4T5cSiPC3JP3QxuZRJlkm/wZhoNvFUM/ViIjUb8oerlgz5Dg8JmrqWs
BSmMqDpyDwGvE29faHsi1DFH+/nzAtzGToNCpkRYZebXDBTTRlJmntfHSqIu5L0m0qppOMxMyExL
ttRtEGAqYA1DQsFDqSBpMX8Q+CQX0G2bfInHcH2EUEnDEY9oZHeTw0UAEfYiJAbm3EjIRF/CZIQ6
uZ/ft7cqWVdrKv2JPU0KgdVuyqsU3n254d5M+ovAmnjz5fDRRacNOQPaK+e2BK2kL6ZatE4c0zCz
SHO5x+Fr3TE1HZPiuhPUJotfwd0VekCG2jVWegG8s/64MKN6usYAuesytcmX6dCrjhmzdWpcDygv
HoqLXdvrcChK+wIwk0pwEbhb+b7caxCfeT7/8gowOTaIRYkiwC1E3PUNOQBEG2pZSCQMdA+cHhq9
hIkyMjgnNcgTHIsHLCtEorpzYVwFxUztHTF9wj0K/gOfTuNMGcSGVSzl34xezqRXy9sWITF6hiJI
GVeax4/zvQznFuJiO2tWtk+RDmRRkFhv0TKd29l7uN1HqxRQERXkzTv0VRghSJ9BPJtE5CLVH/tt
W0oJWwpcPlGmtPnkv6LkqD71iFZR31mRxJn3IitI5DfEc0i0HjiAe5ViVgyb5bjmkhUeFlT7CvJn
8XFr2eTDaEGmK1WX3fbCj08Rs7s+R0T/WpDPLrx7SO3mHdXZHDurwK+N9/As5o8sHd8yV577Sleq
TL4/9I9Wc1MJM/6/fHbscPIX0D+wQBt5ujWgK0PcyPa/HwJeeFkAIQ88yB0qZa85idmkCYz3ue6h
f94E+6EXaTtnCYvxTIPuJblHaXAuCsvcN/l9InCgBGNKzs/KsgL0Mb2G2/3ggmFPjwNcNnej+zyJ
NpD4y1+/akioErywuGovUwCZWyo2eMSsDLBSkdUoNbD3q2GnEvo2vsnEH41LkUWuyLlU5/oL6WDZ
dNYHFx1XAGeBPuoh+kAfCIb962epdgMTOqnVKF5NBKKOfx7qOjbgQMiygnIYDuXcE2K+rJdxBXW3
CAcdF+/tXWwMC0fTWeT2xsYsxyf5ZLkLCf3DAPIG8xCBl+2vJEtLeEV+WJcOMTmpiBFWLNxSHDoy
2efmK43XWB4rm2xKRLvSJfdLu9fa/i/Kca4wbpU+damH6qIj0D66kjWLO+OXYPB7J5OJZpgvDf6R
uWEe36vx76YmlTvBXG7rjkDm4VJBV1Zs+BhYB8Js0OaXFKATrE0czY6gx7dpkr8hMyiWokWRor07
4+LGkgAFmtJd+T/5JdhBxqsChkvYc2rhI9uchsY/Gasu0vfjhZv+zxqDaWodUGIAYBn/JvOTNS+l
VZWROI0FIc7FijTq/gwY0WCYBYC06SQcSbVpFfN7ZmpS2qD1pu//AHZAe+hUWtNVBC4vwkl22GyO
SyaIgOxEVoyAV/s2F8OlF4drGfEd9szKKsbxthNexRkaHT33XDUdjKEMi/ZSmhOToBGg0tO0o3pH
a76C0Pmvd4yW3OTE4iaI9i5GchHr+zgr75OWxzukBefHTMFQRWyDxpeeGb8fNQqM4o9ZtJJXGBq6
PVp17VYzoWgDUrQj5JPU0M1d626t1qQLp10ILa/elgJSrbPPHqhHqo4SnybZ1eFeMGqrm6whDV5f
3RbB7mhGy067gZmwpuiOQa3Z6JpEIxOmFz3lUtRESEi0ypnWnLILRZ27ol+JbtvIW/mMAxxrwYsh
BB+wbuo8oXvef5a0d5rSu+6KG+fc6KQroSXS/eHX9lLLF/L+dJsvqVrKKNu4IP4ybyVcsjqMeTSn
N7HuVHUVCxw4xmC/oCAlQNKT5OhKdRJdyMyTT2l484nt5I+ARp5QYMAvARAQbts2/PZpa7EFW+Y9
ORApXD+qMaxf2aeFVmTkYoQQZi1hiiRFYRS6HiulIkHHYG12mzSdVMu6ykzsmruhS133kopAqPrn
Xo7l0UB2JZ7z17q7vzkKEYdKpwWaTvNwDk9yObrNsMG7qaxiTFbYWtVrxQkJNHSSeKmmkIuw4mvT
oE4KOyMbotBGb6GsdsMSXK0Sevbs0ERyV/J+8q62QcL316NjlsAqP8mkjUKt+qpp2uTeOJIlP2Mk
eZwexa+NSgC6MffdZTwYeGL/rA7xvtx6QTmTPp55oU343N+jho1veUBSP95V8UuDfKeUDu1j8DmP
DVoL7qb3yVnkeh1eCZSfqHkdbp1nvQsGsxjUhlmGxsHWffhjAW+/XkSo/visvKKiY/9DuArwTp0A
M3hW8o6basgg1dTPdIm+2i/FOPBHDpmT2BJHqMIAqEFZGIGmTpSOxf+w9rMXGBC05pb3wlGrqkvj
BQ+QG2Wu8RpUmRhA1EyoBkSTJmJqam+A5ej33fNuaSmhtbwq6jdNopTAeDxl01qboanm2e/funrP
TLFMN7H8MKoXArblD5c5PTpsq6HEGG/vT0nW/vW0dGzjreaFmJl42HyHOAO7XsbzVPPdWOJQ8EgL
mJiWds6UdLcD9YHZokNNWXwDFlbiCBXHZt/MsTgLhJR6sUw+UOvsLtOsAI1lutPgA2K8rdWys0xo
KmVnPPCXuXMAhNAWgSUyKsguL4oAO0qP9B9a/Xvjak1IGqWLnrRwWK6PnHHYHOCnKQ8Rp9EcTuGP
kugMcEyofk7Q0pKobzrsQbLOd2xBHh8dd+Ui1iGslClT89UmlleXTj3uN6xOHYLZZzWA/DgZ5msY
zYrdG8/03ASU+EJSwHI4w1ZsEyKTGoOGluPABB9WvQYRJAvYW6k94Ovcd1W9G8/1VoR/aJn+5/rG
o0Xk+wRL2BWQ3mECUWiWF7867L74heBw8RYloUJFK5JaxaR5Ukuse4hqq7XBuk33+ORxfXRgnZfa
5iAgtYqzLy324V0B7lGBC6ht59ZC00lpcszLfObV5LiFOxUZZEo8ZeItTjiRJMzDG5ZT9cH9h2DF
owbZ892jkPRXkSM0my+iJ4epqiWI+JsiJhe1F3kpbEpbgZitFt4d+I8RoZZEel5arSWa7qYlDFSF
fMCzIP+JYEPWt76tAUbSSe2o3FiW6E//i5cHqxIWoZ+Z7RTeFJ8CYuDs0Jrfjetcln2PteEYLvoy
3NXxqhocCCUuF3fWhYNF6ZK9qzXCa1uu6PsVvGWKbuNJf0g3nkFO3seyOPHABlh/0XqZDMjmq/xw
Du5EetS9Z1nhxXyEW2+SASRK3TchUoMBWOHhJ0zo388ra9EmS9zWdd61cCXTyFJ8Xf5Dpb6ttHDs
7WhYGf/k94CWP5aRkCDtdhDtySnXM6ulFUI9rzlrxqSZ3KIvatua8wHmnLwBFEYI5aLWM6HhfY4O
UUrEQ8lu7fA59ZSaJBP32Q5jDDwYxj0G+yWUKaat9LXZh8LOwgBhw6zKESPxdCgv0F0egKTsxdmJ
DGYhEBPVV793gsaDFDeIZ+m1weBd72g0JdBiW1KaUg6H4Imi/63RvnAtxBkiA+Fy9j+KDF8OYkS0
Qqd1K4QnVXkA6HM0+jkICt4akmnEql4IS1XvDtz0sFlhsaAITjPdBWNnznpm42GJdDgazzy5Fj+g
D9Id3mbj+oa/C+AFPkVvgWLQeqLhQ2Mjujs5C/33KSNuBrOu9r1ruHL4lvTr+3Q6jr3/nHrDqStg
wARa1qFsbA8NkGFb8xMXRCMNtOXuD1H3ZhAvBO0X7NiejkU9TWw4tn8Kuf7XxNv3a5b2t5Cv1+N9
4ULKBPx+73EYkCjbl78K43WAYVFrg3Vip+AQpDPkZKWMjINOmnSoG0E5Cy5VvV2CleD/g7U7miiE
BF2RxLRvVBNZGIeSbOJ3SnzbTKUUo3aqsn5ctzn7c4kZzDAZk6vqe97qqQt9oTBihu713ybsqCwk
CEur4Zd+5vGtpY2w1NlKRWisEXnYV2aEUN4g5YTxUF2sMsfMsZPPdd0Cous2rO5xwKxEEfa74sFQ
WiyqGcFetQGE4V9+Bx5yoXQYSfnuuqESeckFJ8IFvflyROdXk6HhmQ6aXfswKYUSq/Bx82A6lQIl
ej0gOwcZs9yi7Q+ugwcpgPo/9zJlnBoWFumBQAr4F/9Cn1c5wTuQsdFuufIvBmxwh1oQpkVlhUpN
K9jJqSeYBPVsZY+MxBQloC6y09HF2JAJc77kxqimqZjXYshCZHRd6BvPHyKogBwB40tT1uH8Lm45
ZyOJIgKZ4v/RqUVDZUXwjwKMGoW9yYAu02mUyThvGNLU/5fUVlHSmk0jvgYAiVXMG+qrPWjmNbjs
GLBetQ/HuRxhu42Gzvle50prrMMDoFeyDfofddQf7BNdlLDBY7q6MsKy7K8bIRuNeZZlQZAUuBjr
pOMNZ9P6l2JJ1coQLJ74/Bom16HeEbuFMjMNJFlRkN2d8I5BoNbmHk6fQ0Lswuf2OEQw/TWSovBw
EqRDGKAsjsQ2Qvs2GdLz8/cwBWpEsJqIEkDIM0eYfHPSMqJq3dn83bTkdDKPRUTI3EOYwmMOHI9L
Md3gg++MnOJmw9eUuv39/DL5LKMaAYOUiqZH4bh4TY5MybbHeNWFywR19+b3EVXMkVfY02De9KnH
cO+ysuEwky9pkCB3Mh9GUd0MnrSv75cbERrRaAmG6R6zf4/kMsi0jDkA5bYIwbG9XwBFWymQtq7b
BciJ63wpRPgJnpbOl4nctpkF0aHFPQEZoxRxaLkrvEkfljn9cn7HKHINTp4/UotjNZy5DN23PiVy
w1qha8IJKkC51l4dGbahyNrkHUcJWJTvhRi3is5WEYsq3l6Out4eI0a3unGFiUiZgbKZj4uhsetP
3Limdj078jMn+u1Syr8rCQXB9CcNgZpMt56gsbtob2Ld+iaPYJ8PJINQcEEBw0P50EmPOf1fAwex
9rz7nhr2lpO4XxswCnd8xp0FSPjueXT3x9B4mnUV7/YehqWYZVz0lmkg7uwgfAbPm6f2jpHGhgWZ
W0xeWIWW3Pw8a0RDrUgG0yMtNMRP0sLGPYN35Z/jxxB7ePHPVO4aCnjkKJUqrMRaw1SX/B7s2DSy
YM2kpRZ3fVq8KT1IiTUkSXEWezkxEMDzlxlPgFB+F2Rk1RI++f9WAYdAzhHWQi5Qq4t9KYJxdnwG
1JuBvdlWoR51qUJjUnBp7cR6saZc0GlBXdsELnjbE+0Ij3XmV9daW4b05/9EclgNQStaNKKlOZ2y
ZwVAFoUvSLzo7upwfD66armVHPTUxFls92dmdMgWFPcS9CLRhasd5a5c0ErjbjUm4ZiXUSs6IViP
5Nn6tJ+3iIr6EZCccb64WgZkVXIMgN538jVCOPtSoySvZ6W/8aYD+QltRpYpSmrdEubvbLRDOmWb
DOlWNUcRgW1mLEwR+S0RbH04CG6XaX51sl4VHCr2c617v54AtjITpayQvjHbcSWdxzu5cCElT63j
lgdpg7LLEuAq28sg7eIox6LdZRAVcZzLFrcOsSguPDXwvewvcJ2SYrZetbnyHXv/r8VC+pMKbJkc
0GkxQbXOHDaGY/bsnNtndQASKhV0j0jBnkGQZtTa4dwQ5RtBkpx7IllDs29iXcBH5+r6gYFPAPkE
i1vVrlSWUO/iLRfFdfVOHar3MJo/9y19jObYevuGH8T8s58N9t07VIQTGt2w8HWPbdPBJDqiNeYl
Po50fB8PskvTAjM2UO43U8OM7C7MqeqHCl5yjV8dKyq/uFUBI07IkVl3lNLQ0cVWm8gFq4oyOzu3
oRORXnc14e7j6aFCbkxc/udZUsXW4jBgvBofhsnPgw/9cRhGhgc2HmkS2j0a4nEjTnDnXEUzi71l
yX3FSN1HNNwQp5iDhTZ204uoiUhiuo1cYf9EZiaWniq3hiqIX9/xH+iq3e2jRUAAoVgH7FLqbojn
Oez3lDUBeUxUP8YmbsPFM+y0oF1WFp4sbVa2S6ktkFUaHcSkK6vK5KD958H0CTxt9MAIzceVIjZ1
JjJtKkR37943M1wG2KHUTg9NJm8WgYsIp71+KmsO/YmMJx/hnYeu3fQBNfddYpaixFrMJNJRRP5O
GkuaCxD/TSqRHRq0Ri8FWSB2B994hlB0/+OYqy05u5n6DPvDh6shY779UKozMIBWVfDFTDwKN6Kq
NOzXDBHzFuOku9Tsivt6hdUbkEm/DI2Ase2jC8LUFpj2SCD7j/VuIlnx0Vz8+Atz2LOaezXhBoiZ
JzDp0a1KKW1LtQ3Q8eiUvmCXi5jwJKJwMgBjWSO3ZGWmK4oesNv3Uny+V8oS6wsnjA6veAu7wdqp
W+XHGR72FWAazGo24m/UChQWb5zJMISGhfLFzOFPRUmGfugtcETAovUXBFbZlYwc6gxWKRjzgV6K
OUFlItnYR2bY0+PVyYB11PCbFArQmybODbrI9gKQnVDqHcKTYLwkNPaaM5Ia0rDMPWE1ziv17++O
Runo33ufOxr8NmGx3O9z1T4eOjOG69cts7N9Q6KhxFdLmM9Pkw21j2QsBAHh/GpiGXuUJiaUV5Cu
zC7AYzEwUaAh14Ep8HXImCJtVBx9BA9nINF/EuZD57+tKg/cvOXlvLmiKF4UK6QczOajVKjOkw/q
brYMIc7kInBiR8A20hgZ26f1eqYd/bZo+Ol0KhiZEVGYeDplk+/+v4XvKW2O1AFrPpI1Udgi5Ayc
c4mSG+I8XG8SMzTXXYMRla7RQ6iEjPMUPSlITVUJwU1kMtyT/bMqMyQdYUdWnFMl2sEQAzcobOJM
x6wZ7+heCYDyUdw/P2phWot7q/qOM0Tf8zOoIxYkbnt8csPgeklCThVtNwmEarJ52utL8yPA0wsC
qTzpYTL9dxJs3/jCjBPpxWwExtB3x3YloRvBJTTJmGCp/Ue96niyJs0gBTHxg9L2Av54bpPh286f
98TPQIyBLqHMGPnIVuTuiuA9RfxBlpdXQfck6mBv2JDnaDZJIGa/P1PO8z6VzWwLRWm1oEvGIjc+
k9QPyDlhLxlDyxVzpjw7YGYhnVr7SGslGl2gbnLR2sLlLT3xl9U2OtjCW/2kOABUzB055dtQRmyg
+e38D8taQzyBCCqc+CDL8IwhWov8EeqjWvvl01MSsmx+M3xG9l34lUwxCxYXG2A8qDYrNikGWt8J
UV1HExMyPGMtpa0iCGq0Ky22zkzSpwySMrEVuR0oGoy5iXSYW+KTT9ufPSvPEEulc4/YVueJZnBa
Rwr8bJ3c/H9f5qXUdbHiaV+ir3Rh5WcqS7eh5wykDBX9G115d1WSiSth5PXjuaVYRuAfi9a1riEh
mwmpx0wqBq50e7w+jBNV9Xv3QMXAzaXZoNRHzXdMPxZDcAxiZB1etqT1cki9mGYGCVTCQChUXKNT
2vNTLSgs0wU6ip+sN/+2bFaVkyuM+tlTl4inB8SiXvwEZZYEIRfnBKK5cXGzo/nmcLXHtDJksZMd
D9TxsRJiCucJB+jOLBfVPRmsTFOfum4rY/So7epxxFdtpr3B7cZ0QtVQs/TfOzxHRbEVP0dZRFhp
XUIo81xkAce0oZfwWJbTBMxG/OIsLvT2/FEl+fr9fwpnMnFmi63X+DZRwYqrxJ236vmIG0GLX3+4
VEYym1EB4JdKpyMmdmd601E1Nd+m4spUoYaUv/BqdtgpkExutRfCsuX1CrUaP5aFsM/ybpGb3M2t
KfFOD71GegDi/3yS5If+XuLT5WMSVTxusDNjRK5xW4jX0+zTIRr4AUzkpa2TPBApGeLyzCNiDD6H
/z6vEfRH6JgU0ieL+rbtWE9+BBZWBbLGK3WLUySqNBekyuKx8su/vK/8Ffi3s+UUv4tVZ+S1cE+k
bYw4tJrfCVYE3J0wQ0M6vc2JPgZTPs16egjzcUx1MeL6RaeF23vCT8WZsI9gbHpe6XwIXK4BKBxM
3AXiX7Qeen3upiBQ8a1SlWGoYkeJYE4OxrdIE7LBs+GEPeqagVwEhon9RoK1z9fttVL3SG0xZCTh
onMMDOrbQ3ZQsRX/lsUbSZLQL+DW/kqC0Q+vLz4yLCNqrs2LPDoei5CZdqdRgus5nZVohyttFwNY
1/zf53A2AeuPpHOJebxLs8ATUJMJOSrNkhd+UIfbsWu4Xfim+WcBNPD4ZAQ8vDwYcWMPEmgWgqX2
T8yD7R2QTk9eQsHblQteRUBnXOYFqT9BsTkM0DSNxbKIiO1+eL3bJMGWs5jHH5qELuneSPozFnUY
CWlhRelA2s67j2F2DOmt0loyDhtUz3F0U7zPnJhjNbuG/wnUfB13JBNu9XoautcYUNFrS0dpmezl
DHuNGWUDZOMeHkHugDpdTNDpO37ztEcS3F2b2aYvYKem7tDvdfkk82mk9Lb+/5iWqR/NDdlVRpXk
1KLzqTRelWsfwT+KeEQcXEfR8fP7ORj1MhzEbHzgTfmkZMHVh8aQ2UssqzwHuGg9fz7SCN3rWmtj
WwG0FPxGOmcplBSnmbiYTU9Glk68vLnAmhYRsHcK17Ol/WSgB6L/UuUEv5Soqrn4+QlqBNiwwDat
eVqFWIO3jznl5anFTHoLlWqIvdnMa9ZrHgEYn5R6+27uDheRAhVwDwROH1AA1iU7Rlu4CzqrdvHN
F4GV/oJK4tw8Z1YndpAYBa7FdUglaTfRNBPJX97UHGIRsp3C03Z07g+P4abqgEWcHjJP5k/XBdiG
ovfdBhWykA/NE5m97geqIdvGZs1TgB7a4WtEJ0f5M6u8TbMXzkkW7f0z4pimI6o4XO6F68Hz2DyK
aqTAItraiWnqAbo8duhgOjGb3eUfFPHp696pyXSz9GsdBinHlwM4f5+kE+B6oy5Xl+oFVqf5OoCs
yhGNliBEuVR2gESYQ6kplvNbm9zL7vTBMB7aGCLIw7a+CmrZBuLA0xkmXjYhB/gz7Oz9qRBWH/JP
ivvkEEt0+uhpIYt1+iJz99T5GiOYLw+h8P1EbartYTcrbyq/ORu6zw1QS8sksuAF1a5418lqVciJ
6KMbhXXFBDXwasCyhD56Yu6DYIGsr+PTUHkdbIHDRTYsGmaDN4xY7Zkde7o4ACp+G7q6/xSNDEOB
6aekZJcDxlDZZiF9N1flSOjPwcz6garOfCoeqDq6JdvygzmsgcI2XwXV0B2f4rObXqUdVJw0StQH
eYFlGmk29T7IjBOca1+kB9X+A1nKFdlJnbM87D4H8beFiTMEdYGx9OCF6FCCb8aWBPx/5fUZ6Y1w
vsToY402HKIMB1KAkWlpOqeeAbC9pgtenZ2A032jfrMfNg7sep7mD/U4iPq1PyPhWQjGQG79O1N1
EkzE+su2QXmnOdvM8dY+6vRjA87iiF59kcboXKYwHz/ovXVJpYC6Yh/Knje+dFGcqp72eQfsPhBa
tAfGUMKf05d2pheordCMkLyRnh+FVS6ZCVXPKCFAhpS/Cb7Xq7N36hdr88w5wYCKENk1catlrvng
LEyg/nkc2HlSB0V+85QJc/Ev19RtJjCQInrF6SZNsGYh4kAu18KD5APFNBQS74Ecp/VBlxD6CKcS
CVYpP3a1hfUSlAbvYnYZIbtef7T3w4jPDOwAncOZEj90SPZOAiGvtqcg7sZotkhR53B2KT/otihE
hOmxYN4dEac9ny6F4J95U08KWr4QH3g/Vy91MZTSjCHdRlQMkAxq0Fhs/QoQ1sBeY/gb2JUrk4cJ
2Hb3nef5d3Ccu2mfyMPRw9Okn9vFkrqcezbQiLS0Rf/n9uUEU9M7zhTGdDZRnrx5Xo0sl0AVScM1
IvezNa4WBzL4Gt5bwaxVBBmFqT/fbC/A1M/aKKKV/gNt0IwxWGfdaJg5ubhEU3v/Iq0Ipty08hbH
xuaDBf98so2gpkD3Au/2nBiNBjD7uHBtdI8xNjE6LuSb3orkhIVdelDTimC6DcqAkqxQ+4NHcBV3
Q7oj8V9y5SeYahCgfpvjb4PeOhhF1mkFAzyJbXTZSt4soa39FYooTBpt2TirmVTbzuOlcVMqO05j
ZrIRrhews8oOZJj5a63d9GB4yUjHL3kILXlm4OrUrAWwOQZcKqey5zvaH1D7qilSNzn1xRA+PuQj
bFjArY/pFmAD6rWarrrzrlOA0MZxoaU7YfWpvQGx58CQgkwiZeXecTr/eVwU4z7eQ2CJRWugsvoB
9RA5z2R6xnoFrZABoI6cQQb12gYWsUewHCyO0izrdFgjdYJpx3QYZX/QHnINV+s3zYTyuZZ20YCg
o+t+8q2nmIJYg1tCCxCBWDa+yKs6K+406JoZ6aDB8k6RXYnZPez3+8qrEfR87vMYSK6LMvgNP1jf
Ol0enYiUpzs1E3wRvYxaknXdJki94f1ctQgcHj7iUXNrdPUO/Tk5L3E3GtVxVg0CGXVgARIlcE9K
WFS+2V5hiastUUJGj1nSepH8DZvBePbCwhpAViaZ+K2Tc/cIAgB8f68ZH2NczGeQTLDrPOBt8QHJ
BWOcmK0Yw3VvRemhsayFJqw6Zfi6s1+QBZbjNeGRQZgT1EJp8GxxaDxiMv+tjux9ng1qaBd3sl9F
if47d+VKszxWJV3HisVTmezeV9EMceGDF2YMfo6Pd0rhMsfnH2z+MFPPymUOPAY5Av1plyX3+pDE
ye9WwmpcOHGHGLArIvi5gbWnobgmlaazVbjNhLcZg1fMYn1sDXXnngn7GXGYfVdOuDXQCBiMbQth
R70gHKrpVYUxKAhRmO8poFZeGNiqnlX8m637S3K/YDiorjVlzwBPr7jVLxxyb/u/vP0xaDNU4v+m
HjxhEsc83Y9L4Sp+ojE0vfe7DseiRIXfpahkGcU7w+e++NZ4fku50aVmMoIK5U1gJ5EbXkwYEDus
IauKLgmKWR0ZnKxFcjqCh02JCxzCQ7d30OI6sy6A/e8JdrvKIZQd3u1VE9wx13aT+ZWR17Sm0AeQ
FwakqsAY1R94SnWo0Pw0o9aQytZD3FO4l69eAGCDXzrN4Y9n+zFgFk9J+gdpGZWLvBfyWXwwsHr6
kJCl55MBdMWAMaZISOCqi4DM+l87TZONqsaAaC60tC8hcCB0f3/RSlTbie3LixW8fgQWXXekLp5u
z4LNs1f3QWSLkzejVsrTkArzBFfCq2+avNTtVu13h6esS2Ov6j2/XKONCs4fFoHYj8pI83SKyjEZ
08LOTJsAcF6wdOh3UonpCKfusRaV325iQiv/Y1gfMhJN10GC/kdVbr9+56TdUowUK/4Kx+xx4xTA
9czUkxl4c9VHv74Q7P/5pTG/+yhjmJYJoOKd2p83OrDCll6Y6qdWuG9BxIV8Oba7la/J30Ln3shf
66mdjz+I/wOIPohkzCoTyPVXiBlJA6V59CDnWTY+SHDjZuJRe7nAu5/JuKaktPyGBMQvPGEjOXBw
rYxmbQYElt3MR4HcYaVsfqILTe0nie/EyYKsEybn3RkY26AaKibSWRSNWWPvPBBsts2LuodUMpts
ShJenCQRJ+EZc/FVXc9u1nkYHLsmh5rv0KrAOgT0tj/DIQykguZJweG2uh6hA9WtO1j9ocWxgCEx
2BSS8SABmg/0SYaT8VcylTuptJzbVUWNR7LpcqUlo/Gm36NgsM2lEfKfa7ARddXcf6F89+TNycpR
jUJ9uY3KlCB9tf27/NVMslIqb7crXVePXSRT7MsqyAEwCFqtXA2/BXxAQ0cKCKJVcWvEVA06pmmL
E7ypm46lgcXv0Vbl9BHGXR2mLqT+ZRNDYNaIvBSlXv2YPlrIqu47JhcpOZyRYxWzJAEtexNnKL7u
D8GY7fqO+eqkBEBKOsX8Y6Gvg6EfvkgQGXlB6xYflCH1kRt7cQDy22J7x2MbVitiPJjqJUch5Jaz
ho99BqnGylGu5fD55+Cej41NN11qukIUoL/jlcdO5sHY6K9qLw9BNeYFg4l4wuU06Qkjac1ZPwBA
QUQmGAjeJ4b1gzDfS13aobC+ALuaok6ZYj/zKUpuwtA8uUhghwJY9yFMqMkqhHPbIQOd1pt0Fu8b
RhEzI4Tk4G0POpaInMkxe2C4X2OfGisGLxWmnm1lEY4cykG4tVE//fJDju0Cd+5IOtY6SSYtvppp
OTHrUhLq3GPKLsPuIIieoeSmV7J1ossrK+3RLDmyX7ALNCuT30BZOsMXW4tbAIL2ScCJtijQ/vhv
QjZn52cyM/yeR9poMbUTqxdwdMT/hw8Bo+gL9zcig3NH6E7+9NFdG64Vka0H8+/wCmRupjuuRdCL
WfeWN5Rf92niIDQpB9Dj2Zywiq+AGBg+ig/UVJh6DoQSZeXMjIF2zf174QrQsTAlcA1MkqijD32N
Hphf91mFPQwAaHjzqucMAUzSIietyssoJpQjtLotFH1n2dFfA1rHGxoMGbpNZ4/vSNqVXxUVRcMZ
8nWLz4I6ouQg3o+SUTZlj9Vzn3hqNX/uNHDgH8/o4HCsp35oVd/i8q5Pfq5Of0gMtJ8Skl5sXq+J
CB40eu7opV+YlP4nJ0q9ypoEgMXEDEdcsw4VJyRcd+/UkB9MgEjapsRZPgZl2qLr+s6sTA+qhSWp
HCXtvIRiJz7GXQOWZZQF9VnsFk1kvmoiaBSp/K8S8Hb638S/w51Dj4JbgXtTjmRI7O7u3jNs21FZ
8Ww7Qs6pmmtctOaz8bwHG80kLhOI1vArQvqNW2IjNxnfUNqLWBaIhgFLyE3AfIJq+g1ObhaK3iCr
EnA1JelsWosJS+5r2l9cmcRviOqd8yimRl7dzgTTa7y3Pp24WNL/zZkS9+5n+br+MO2iUTJP2Iqv
irYoeBPp0T4nIiT0dFbvgLVhSFb2rklYqsrEbvQoLqC9MVJN0oGjnwpYweJK71cQZ9P3WJ6g0PCs
+IxwYJCLP4W0tmLIsQhQQrytdVMO/YqiX9M3CbqsV0/e5pe80zQX4XdkZxG7pTr+tWVofm7BBQj0
RNxl+pCigrMleq5KToj0kqcmFmYgNQowt0SqgSFZ2xfZW6ivLOgnTB/EvEPvo2LRAl9kwVtfGqDG
o4dE46KyKLId/AuWxnboMXpkDvDddI9XWtv+xnpM/EEntN9q4hOqOPnow4L8DGWM8Ffzvy2+GqNU
GRCip5gVSTlIjqEvqc/3PunYz70xJU/n9fV6ypqFGAxaRL5aD9zs2xWao5md0I+LVwmNvqPTEfOF
n30GCKqXYCVW/AQkXPpd+ymwj5cjLVJ6GsyrRAwdabirwlwc0zhFSVGjkc/dM7YK6BIGbuu6l11z
eGWS+rz2FfLbNpufBTInhR4WzeCiqZhlNckb6cpEv1PZ1a8QYXfTb4YMCNBvs0UpWV23V+vHXfgE
hLxWZgfpBBkKngmdmPNJYTCMC3+09PkDSDx3VG+teuLMfmUAiIE01YhmFCRSnwD39pxLQ22RtPwC
QTbENbZJG02M48IUlm+36RM90zfX+tnUrs+RU8mxHHw/pKUrqDG0AaXVV5qQ/hAdm+Xmg12ao0KA
kZU1c8lZRgPA0I3xEZApJUoP68gRX29rFSPM3p+MjRdywx/ulB1V3OtEAxj9UgJwp3XpfkZpfGco
ti3LGI43nGYk8awh6CQzkU7lVz2JchxfCghghJumlRh7LhVYf3lJakPll2p/HYN9b6hZppuIcsds
63KuWa3toU+K0JjSbFGHIc5gBentUKxLMVYokJOSXTa0y9Nfm09e1a/qyMnQML3FJRLADqYAETCx
+Ey7eBXEfSBenMQNeBNLoqpZLvVFY10uQ+t9lJttf0bcW2A9SAi6gJB19TwwhZJsHrGbqmeeNv5Z
+LS8JbDXOeXxp0Tl4rJaYgqXGVj9wketTA5ZIuKzzzyXgbIQf0ypxW3D1a89bLAcbkn1lb2OLzRZ
CQGhKqi6V8TqVq8yWB+Qf27v3SxwizqkUyKq0+jhaQCtoxlQjmL4GI8dYWO4XeLEIXPAgNFN3EBN
tzd0GIopXIG4r5vFpuyX2lJ/G1mJDZI3BmZsL3EzmyAPX2RfeJRcsW7q6gu6KVDbzXyy0tPENlIf
cqNtmyWgkMf5U6ZY0hHdx1rISB09hgSukDrayf3Pngq9QY9772VS/86LiTw5xdR8HoG/tu9xNXaH
DpdgzDM1SDVlzBFytxIZroGm0f06avf8tmo5LKDHwueH3PNfhm0El4XbchQedNiAJwsTlrcSnSsR
4irsspbpzqHnfY5rPjdnGlPTOgj/eZY/2zKpc+0ZvHvdUfi01jJDHtIwjqYqTMtAlrbCb69rps9W
dhX1mpvN1rAEG7NEm/lxCH80w6/sqJltcLWHNVxI7yz9F7/i5GlQd5Lxmpr5rZnTfgFAwfTpjhBh
+SzIz7JrpS3Z0VY4qha7bXE4ZEccnuZDDqGU6gQrZ6HeiHRQJgzD409C8en338bXLxOS0Keq8pGD
3bVdUyqDbdF6VOgNFgwn7JZ8fk8wfZI+pPYtcGOHEpHfmQjv1RcAn/ig+TZNLP45XtmYWuabjFUp
rrt+f+LqyQf/oUkOQ7o7iUefJ+DANwozgZVZXyfygiqJYm7/5QlPMPHom72rBfiaxwRa/lCKhJa4
9+40EylxBRfNeNXw6GM+zecbPiBTR54i3l850TCfJBMU17hSqoXQiXHtZUUqlG24jS9jPSpxE/L4
rxJ3NlD/ZEg+pnm7fVCS5upqv9KD223sg2qrWie8UVZiqZ9YWT3+7G+ijTYHBGrfPTFf3nCYUVJx
RT6VoUr1F9ikrBOn757XoXVArkTw+UzS1I/YihgBsUznCyiLHHV7IyctvYEYKmbenVo0UQ0leFgn
17b2BSAMjALJpHStaX9yRZAffk+XrNBbxsyLh/ckB1/lDsYRtWGofYXBSlvu4UkPYQWpOGUtqjAg
jIP5gINkLf6CFoQHG5X3FMDVqQTTTjrA3EiQmgcVeIWj4AwkmUwLTc8cg7T8Gqyn3OT/WKaSZSs1
r/mXgtcY51I/ZMb8AO1wAW7kvPOybyKBS6KN0apX3OqydyP9Ya3MdrAljh602b7FwQLRGCneXkl8
v+lnRTFfbq/DaD5O/bXnUh8j86F1uTK3RzbuQPY+wJGZzfbrMNMZgKI3DQndj9+MzDtfQZDBv23D
awc3nj1knfAmciHdZHgyltsFiFcI4edTsAHcmAnlALfirYpe4kmzby5sN334xDO/dg8sjQkwNbIg
W7TGg5AIsSS4fIVitIZ7i+1UxQcoAj84nF73riXdHdbcNDzkPWQ7m+m6FcHGW+0lH2aLnos7ZtJ3
fAcpYFffP/RFkrYpYH2z3u+jiQlIVLcyGS/WgNeEouDxinsF3S7CMWuo9521wCcDRgNx6tBsal9s
wWUymbf+F/wdU97TIsO5/TBxLlb4+DeQlZpkYD6LGz9RTTaxfoJWJKPZ0zHxZrWxffWMbrtPAh3i
OQLv2a0KqutJEZxp210veB+wHYUzIoQKaibPzgy1UgJRXSTxUnhLc5AQzwR5Th/yNktkkSF8VemU
BsUhgRZh6CAWRqbhQyYMcDPjC7iPBmp1HJBAVbjD2/TKkaODsiwnE1qNEp/uluuwDxHPD63X4bIl
yJ27YCc6zGcr3AMqyHDQcu++qsdW42qOorBkDh636Qaaq6KCFPHqdlEoA1VMTpIm5KD9tOfsHWlv
utQ2Fe7KGe225/qTNcVPQafcTn0PgwCfzcMjk/8aoSjsBJNwdbl91u+UZygthHkYdNNyYzLeqRx5
rZT8sbMekyNhsWOoXODFwkvOMlA8/5le4PYQg9XibC4Mn+CHLMnLq2PNV372xRsudoPTDGKzIG9Q
ipZOm4m0PDEHg7hmqEhK0ulcI4dl7Usl6bijPHWEi32O32Yjyb9RIXlmznmawpGWNDG3Ei3y77CT
U99tRCgg2LfCyNcbjm8B0qUnAdonWuFDyvdO49OYKcAETh3Hsq5fKto59tk6jk/mABC3vgLdVmxh
rQ3czb7x9K8pAWahEJQUdpDaoxkC7BYdlEk/du0JPflq8aCkXKyGj+tmvqkncmGHzIDr5spEdnaQ
RJIiIPGRfHXClxArKGNsIMM5lij+gbqJUXeW8NRPNu/VNxz8+NM+2gm3JowZv7cT0aJka0PhZCro
911aUjW/XfqGa/BfQRo9SH5pQ1OTxPUUJGDVxr1ZdY36Rp9lW8Za/YHS6UhQedD9bb4cpxne9Yb0
sng8TqBarWeF7r2d3lszBW4IWlTXFG8jCOiBZKA7q3edZ+h+bmg9hrrR92ltN/4WPfbdGWar4U0C
GrVmvVLajXZWxFr50UEgeAJ846j/Is4hueh1q+AMVFQbUOwB4/L2aQQx0GL9FDdt5HDIc0dqpz0X
B6d4KG0w5xB45h347+FmdgM1lKoQee7FwCOsegn9NiaHQLy1b4z2nEsQrLYClG7m1dAkhzUT+kQR
owjfcE5ydxsyY/kDQz2mSZ+m8ltwb2j7faj1YRS3M+I8TYYai2nSDHrHEjUAYviRMgvVQ7KeH4o/
Xx5FA9GxnhHAATceHKm5IykkpTUunGLQoH56Xr4BMf2TGPkTjcMEw92VZb0hJM+a6zRntWHgMHHA
b7F2J0VtAsNgDmxZSv34cXM69TV9Jt5Oks/zqBz0yMwy6XdZc12JtIWs8tnyN3oA0rmGrjziVCo+
UsRgGBVqvFErTl2fno6U53vIPX9zAhFPpYsTyrGjlTus10Xh5dVJXh64RzhG51vstyUo9LShGHir
TbgCCwaqad/NON9kK/VWS3AaQGsAwNtIdYkXNk3/vLtluBVHC5mseAb+36CMTw7FfjfTqXbFxd3E
olMPgVBGzuWtAvUiCfE/ECo1U4BS6kbuvcRNUbrPicF79848UEsH1+wwhw1YsPuOomIH2oG0cIqJ
f1nkwJWyVDhdLanoM420ac6kN3cz7GKRhv+PK3umtEX07gkS51XjCx9gh4QTm+V9PU3fjlTfoYeM
O2lUJEObme/wJ+rTVS47Fj8tmYily+WQpAVWx7lXVw388YeOmgRq0lJYaNFd0IEXjfjXSB+ggJGi
XFFdFDjfKLVQ080/YTyynTVBHNhFcdkah4/MOmS9qfRrceMjF+K7uxDLbgfUgk/TKzpUorXpVMI1
P7u4ewVGoYxp5Yhj6pb2/NW29GNg6GRhmK1rY/Tnh7d0wLg2pewthST/2knVdqzRv9snjTKhAIJp
24ouFBihBcjv2L3IrQkI2jdcYTm3lvKtrtdUlmAvNkAMlhhLOmsdMj1tyBU1h/lqtWDo7RDeEWB4
A6xz65HfO1RNMLhpaJpabUgcsAl1H0d4Wzi6gcJ7aGZY4MKE57rfiDsDrABEpKuBzHXBZ5IDnvd5
ZzxbAOecqyNoJSkokW36SH6EfJZ//tnIPPrSADe6irigSqxwS1lYoGN88WdI4zSwivmwVe/MMaXV
VCMScpf7CwaeB6ZB/J2tGtYftLCpkA4cN9ySIdyJAs/tlqsalaf0r4w3QRlDXIMfJVI6ZdOSX2sP
Fcf9RMVCUNi+Lewuk897EIi3LQW96OwOphGsmCFLFKJ7Zd4KINi34U+LI9Kjr+voH7yudHoF4XN0
UGN2WT1DZyJNLNXGCaTozditxDOU42JaSes/cBUwp1PQ+MXB6pu0vc/1FEFpJFNI2XCga7ufRjb6
VfouVGMRMqQjv3WEP3EZuXabKCXNsTnStuPmworUy5Y7alNPz/87DrphQ08wobDCSA9n5M+W/yCZ
iApx6FrKdXxhaFI3+Wlsc2tCH7xlD2FfPKpaEJpAUiOnomWTHeLBtdShTxrge4jl/mKu2MfmAK7V
p+ZngPFYetTFxxzgheWzkLYJDSzl1mLyZKhEuohliqkt5OdxHE1BNXhNsIJlUjU396fn+tKlB5CN
4o7jf9lXiGXzQrLVSY7xkrHMCaGXLUUezIQrMGnB7aD1RR9ZL3+3eiJjqpss2t92u4GS+CPhBvOK
mZp0pDXgyKAOdn1qIeOCmXrksnC2tdTFv4kAi1V25D9hT9w84lVkYy8rqx9u8wud1JqCU4YcLnQ8
SqMAxe04AJIkr0JIEHHgKqmIUvEILxtRFf1UokrW+VersxIkG4Mp5HuplCm6HJyZKszweA5c7Pd7
tU3Ig0OuJZ1SPbJ83QNHMCe2DkOdI9GeIGi3MI+uiSKKREurDqG7A9eCvqv2ig6F0XXc4NQAL+4/
K4V7PFr8r/XvMh+khJILzSB+gaq3bjvyiatmYoHFrmSsZy6bNGG2wbYDe8fW1nIKOAyjT7+72CeM
LuTCUa8SzzCtLnklu7f4SHLpIzx0vBXcM0pVqVC/mECyUsN5qDYR5zi44blMN0I1iRzIRGA+2ZZi
AEutnUZsBWRAO0HytZ8Ijg+p61ctHyCfy+ArfXlK6EJKp93LHHihPwm2ucARFmCUw95XnANHr4j/
GviCI4ZaFTW9VZ9p+GF76UpKUjtTJ+dlAt90l56+s2AY+LTVtQYEaMNwe2DzOWH9/lVPns1q3kcf
dXcJZ4aMIWkEF8qxmA9DabGtLfJgSjmFGL5yQg4idTVnefNLyz6IwhkiHbIWJyJAIOY3A1inHylU
j4il8JtGZsklc/5/Q1ClXGkF6QNU1BDxVxZJgHdEdHtmpeV7gB3qR9clycz+W302I8z8LjYkZxl7
QoIDthOx2YDeSirxd1G4U26W3RRCpJ1f/cSAIUPhsXTUdMFNRhEhVMQOShdq4pP9N2IUv6Ra+8il
AczRZ0EYX5R+xuoyNSOF63QciIKApoSQg/qCW22OyvnMvtPjAvezBweHkv0jjcLSLg14t0T0g7Cp
22vFNacwJih/mp2i7nCrLZ0qYJlOjoJhQSs6VRyIzxqZNlkYhJMqhjDTLu+n2nInG8F5IIBp2J7o
V6qy+Qz0jWFfCNQHpWAardudqgMbby5/nngpmjXkWy/MmDG+rTmREv56d1KIL2O/hZ/Wf9tIzSsL
InXtEGW5geMbQDNIvXIWbkYucvJwJllm1zMOId/cY0KqZ79LoRBNYYJTl7FOZszCTb/aXr2woVOX
wrVXhMakDID3ztU1UF7iXyLRLF0eKrsq7aBuqav4PtU//LuNohOcJRTOUBiNSU1diBp5GLaYzmic
UvcqIyjJwMj21cZwD6xoEDIYrp/enYIiEbPtg+fziOBQFXxF/cLuYzHpoiXvgZ/gmmoGwagguslY
rUwzMW5bpkoGEgMIjo7xYytd1D4dSkaRbNqkaGVisJBoYcdBKeI1gsN47nLzF8LJI8zxCspAuHis
N4WyZM4rgp1vJRImXF9+KYulsEtiV2HCGAarn1cU+PCeq0F8o1gySxSJSIgqxcXQjHsEnrnV1vTr
VwJTEwI3Ls+B+WSY1hjhDqAU2s46FVzOjskQ/5+i0pCbqpyXUDzSrnSDg2t/hNqilpVWyMg8nlW3
FQxa0YxxUvFxLvxhWmSI3ia9yYx3BA+Rfl+xkH+cpJDbPYHgI0QzC+Oym3oxzWpQJDGpBdLbLYYl
z1NYC3NGEjfuZF9v+C6E3sCp/kMxUcXKyXYM8XilEYz0BGET8YdrD2YtI6/6K1qWv+c3hBCC3QKk
MUNNxaqMP4z3n8r1htITFolZ7VeP75tTURpRZqUTS73LP5yp+zjtzsLpXY1tf4S+fzee3A4sN+gx
R0JD6z6ycw1sxJHt3h9F3on5sN3rrFrpcfLQtxppwakCrz6Y9NahMhNosrwRMsO51SXOmtMPl96a
LkdZaqp1mEPlycR0kf59Or46+STyEaK8fIsfXAR9EFxiMjkWd3+1frVCwO7LIfdGwXq2kfbPh7Za
+D8unABTsrCCm1QcQxtnFADf/ULgRmTgEiIl5zrKnusMw26rl4GYQsvFC4TQzj+9HqiSj6dbUmTs
QdO5fAXt6LbZtEAmW7or8apqm2FwQMkycMcXKICgibbwfLev6QsYwc/Wx5itxTbpWEeEmraF1h2q
cO0t+K2ygCZ+4rCHIbVt1tC59rQljQbmRrPRRkAtISBjOy/ly3eKqt3sLkz3RfO0DP7thmMLIan1
WaN7JG3fRINLzePgWYE7co9h2bMAomEhjN1X9BmaEpHsHgkmGggVQEoocPkL/MPZiYX+WjsdFDhe
WLdUHAIAv2sCqhfFYnbSvb4/Mbz/AaqyVlYvRoXAIeGn9tD/UzjLxDjI2Xp/m5mTQZMMfdO1CZz2
y7vtdiGHFSfIEKFjLORARD8zNzlTsB/ie1icO8e93fq/pMb94ookrHbr+5XsMymzoibX/79dZ2e+
bUyUXl9/OQaIwzIww5hVPnLOa1nQXSpVlC9C+L77/Tggj/AWVbWIFXnDyTPMLU+Sn56h3HQyeXms
8Jmz7vsTApQpHZjzOfc4yt3F8xPF81CmFcIsC3Z0tEYKpJQZT4pfuqfBqjQozU6jkXVrQGJoA5t3
2tHL7pR2tJH4zTzx87g2yaMouJEaUUbrloMv6LcxgPp0dGpTUX0LdpOuEp7Swnf7TFSIRTD2Nt/R
iOCnyAUgGo7LAGzxZdI9yUPBGzpH864Gh6noKNk5331dMPfisAwfFJlUdsBtoJXR4KmCCRhjlAGi
6RKXLLpSlReSbwTFSx84MOz0X9GCBxRwPqdD8hfybzW2zfoaQDB0/AVhBjflxQPrT8lco44dwXud
OI5M/KVUUz+V5IdPogjCw1ruNy9VNMMQpZtwxyqizeq1zhQiJOl2VzAT6KbKPASVFl+VJ3t+ty14
PJtQjmUaqoCoGbPWxnSCXVT6h+/n0FEQ8C6G7jSMJoFQtSPmBALHcSQp97TLCTbgGG2UiVdKY43j
9D6VOCo/NifuI4yNqfeFIoFU45QosJJwVt88TwX1U56WDiJfkWcDClOLsnusLph5Ru3SEoJGb36b
mBx0iT/2gRPLss2a22V4tFQJd4BQNpKMjbSe8tqjJwULBBdKGBk4Fon6FjU5DjwyjJrY7jALf92s
lvjP7UgsiWT8uvaqAl4NYknusCtTzvS9JIzdWP27XhAOs/7WhBlaHxQlgI+WqAvD0vhrsGB/SWDZ
F2rmQEfQ8lWaBLyUl6/v8BIk0vUKZbuQfdZhd0bOWyBhHRAUj9I/HYBsflPIl1lmafiPhDlY6dBI
P1LDZbxYdHSR9iILfGq1sduNs32jICGXbSJw8576Oe4HKRKDgIB3WfYkvQfAE1eO9f3fEttUZd7r
paSRzQtSS5BMbvf79vU+fF0jit3QQPfqPQZw4E8bjCMRZQ1ogTOFSEOI2zT/YUe359TGp1yhOXVG
ks+Z/cNO9TAhyvPyVrM8tUPlmrZKVSU3JqJAB5SZ4KJOSryiT8QJEHniTO5I8oI4FMw7gbDoBZmz
MzsLtH/DSWRP7y4DmGrvFHKZyb8j6vPk4OMVK5SFcagLpEk3IAOUQw2kG5DA5Na/MAZEIA8Qc7za
GoWfNzSrE1IjHprq2f4xP8SkFLFut93ayrIaGbZUiZbJFJaBKVt991IaUlamoz0K3wQ31jm3PtBE
vhUuzVEBavBhmBpXPYUuJaOwl1OSuAzdnJbf8BaM1WzrCUKmW4NCYqfSkgeKMjUhlJ0B8R+kxxeL
s3uhA/wfkd4Cbf+zo1oS9+Recti9R3a+eY970/nga/OB5xg/c51lBFcDzj/bhUBbCZah2cQ9GPFm
+1DfP2qp8Zct0yomb7ZggrPV1mwkHhzDK/4YVsGm3cTKqCcgbsqnkAeFf1cMRY4Hp1CmyypppD5u
Siz18S5rkc4m0Ffnbc72U+oFZlHNxSsh63wnoGjKc8ab55SZklTlK9+8pDWtnITZn16WjBCx0iY0
0lEZly5Ame7DE72CZBhKvCcVvJp1TW7hducxLdXIEVGpfECshyLefLjLYDZl1h7GXVadTB3HXtH8
Nx7i3JuDj725Ix7tiorL/4OIjtUDKVD9AfoNwN5Wkeh3+GBAOHHADqEpM5AIweJa8aZSdTZKEB7W
Dq11Jg5ZegVx4guobda+m6kQZluHtHF2Ka8ouJtKGOEzdKauv25DFVKPOoQinOEbybvqat3T0HV6
8jJyUMYHyhtXedqxfdkY5oFSNwNW/5ENcn9j3aCFF7p+WlQd4j40OwsUe/zRVfZdiiOHERaslE22
1NeTwj0HOxmjZilQbwcQXKfB4dZ7csJe05dkIsww3X6V6G3hWtodzEmdWSosTPp/TIe3K8jVKKdH
iW3Bi7eIIxZJ5Ewor5mXcCEG+238+3yB0XXqIVsCbcPXnidDqvZuwUtha0TI2SybweC5gLK2ZDc0
bsl3mvV7ZJ4LtAv841Yh46Aq9ID8ywg/TTo4QeX+vHE7SoH3JoawQ4s5WDc6UrDrppQYAHAQBfmS
XaDIqLRUFd7ApsIPr5eZzz6Pc1d7/j1U8ZWDB3sE7pqFnIqOOMJCENDNzKXoFZ0Lt1ESCE60WTho
NB0p4FagrC8+abggJgdkdYBzfjTBGn1Qmqko55KEs+9Yva9dkYxNhF4L8rTF1NaVbHfx2DODajvD
mflTCrc6m4ecmuaOxJQq8m0NWJwzs0eqR4kafQyxlz0zb1FggVu79Xejfs1qNPgWEUGbmQxRfZ7e
8z/j7g7MuQ7o8It8I+PsGNkJ70msNx7paqMUG5PzNSyClRJKyt6MPmDK5mJgP6XtCdyT4pJiZgAQ
PqUaRmfi1/Kksemkr9+DtqKQktUIQEXbwvnfa5HyUZjzTnIVy0GmIZeqedY9tGCQkA+q/cbbICf6
GgTisUk5WhVJr13VGEuAGkYBjMP8Wg/2m72O6WaCINLI46sk1oYiIlQv1WjJzCorNYPhPR8g7mc3
JACY4GDpr/dY4VWruslP/IwiHug91lLZh2iYZMCfU6HIj1BYQoYBfN0xq1IpgNaLpZA5VfXQWh3N
/dvqUZnTYp48BkmrI2hPQIifHXXlFdOXVNrm3rOPIBmNTppJU5OAAPloeY0SoVV/SxaJNrvUCn5i
dD5171Hj+ApcR9BB4E1i8Eo1I/l95qq5rmXd+w9Dn4WWkBycBPtdeNkSe3neOC3zW1ETHSNctvil
ZIw1RL0BY/kMxpnFMz9htLH82DdP0OTh8QL8PNZuQloWEhHMwFOdVQPQgi8E2NYejW+jJG3XidCk
9SNN5jHW0aD8K9iBY249hHYLneVbCmnKY+D5bOZcEkN87VzMpvhFYNPaTfEnJpzuD9LTMNLqHzfx
Va0oanVNa6Ebv1zvMsvh/O+yRCK+DIgUHHRPmRewaCiZRRBtSiKugF+cLr9CADtUvQ2aqllMJNm9
oY88aP7zi42rFv1VlWDQ8jE90e2tXFaj5GvAOXBG6KwDaLcIqtgLsGtxXHQDB76t/43O7dQ3RNzc
cXP4AgUANWa8N/HClAVFQdiBgiNqW/mFknW8ykGf0kVikYf8nnj6XcUW2TAZRPnvXGBhGSP+Vpac
WUDT3FHG/2F4i1jA7KCInF442exBMcVx6N54ikftxHewAJmyrhme6nLtmgUJ1QyxTPPy6Uq/33g3
JYw6NiTd9CgpkbPOqgiEufTZw1lrZv8jVvxMCQcbJJJndKOXUYnM+LkEahE2BkCakqlmAsR/aLO/
cajmbUpQOuxGUBWlsGQ4FcD2y7lZrblSKfRLlxQL6IrZLHhXyTJBlwWQm/+XLSQbz4BSFaZR/BVx
7BxbKzHb3JtBx+g2hstswHdlr+Hbn8IgKUpaPlK8YRHOOBFN9Xp+Fv/DEWL46eG1Ijk8enSTCd0+
JOdUF8ven8IQirZvGpUvnG4j8QeCAkQBPsqeTLZRa0v5ZFgKr1dV3cx3IXap1nleM7MzhnqNkA+G
q/bCGAEqE0fiR8oDjbhv7r8HZ30Kt8k4QVPoiqtIPsh8qqnjKD4wrazBMkHikzQNBliTEcA/vw4g
efHS94p80Zff3ksOSn+BzmilPlLMMlQkMzJZTfyEbIsQ6WZli90gzXFzRlgkqGMIVgOrNA5qZKCZ
o8uq4JKWFGfnCN13GaH1+AMb+6gjm2+/SoOzkl3HffLglE8zhrPCdKSOuqAKUzqkoBAl85IeMEVQ
oFeaMfxH3DtoJnHIl7nkCKtqBWAsTXVUY+ZXj9HZoeqmc+n68TUCkUXHq+cr2pVjkYUrqD/DFXFJ
IbEVMxWKaaZ07PGbsr+lqAZidpCCtYnQYuSXeWeEur94CSKHTakIdrgOOGzyGmlZ9FCbMqRc8JL5
ZbFCjSt81aJgZC6ButrEBQu2pDGBOtDgbx//3Nwx6u39uLjsSy2HG7aY0dNY4bV/a+JNGor2l0YH
7sOLjPGPMlGAdGU7muI77lVW8YjXCEpMUPGVGn+TGPViz/xmmpOWaWtwC2ahwQ3RdvxnXDJgbTGp
xHg+IC+2KJ+GCEaoE9Tf5Z/E+By9PTEZEaBCWmt40d/Yeo6VohSZ3F36dXXAmhhJR5ePPgEQGHA6
jJpQbWHiSPYflHypMVA7/feOsQ5j3qWdTr1wMzPQucAPUCfxl/w+o167v+yqSOB2M9vpG4MZ5pwz
kmqOgsOdMjKL+sSHmEiq97cx4WlN+rwoE8FYxo8Red5xugTVJa7XRyV/NyQfTak0kUUydgRUdD6X
npa21401pk0+L+LcP1076XXv10gVH6nWehYQ62SaJN9TJ5uS7WEAdH7JaZ+9qr1ZWZh3cbjI+L7O
YyTmmu6/Xt3lWdYkzNBlpwNhsqNAI3gTW8LaGw9qhiCFFGSnwtuYNXE76eGLOGLqA/NJIcL6DNgz
6pDzAVzakpnO/VAaKfIlASNnEM0PUZhEBGi1O2rCUlIZGWgBZktNWsqBvoau7R6wYZd4hU4HDk4d
JQOtPZ49aqEKKD7mLVIYo7PSyCdK8pdw2eC0zPYUUz82yV1AQT8iVXIOVdy+maVoAzTCCbBw+WZo
sm/gg5SwV5+LbNrgchw5hNS1DSMz7ujAmevXidYjTo2jL817bsjGfknOVdqoA/5brHLg753J0Yt/
hRLe6sEN6O8bubBqzVJrmoNZu1izfYciJGmBJ9TuyXY8ioHjetfi+od+l6UlQFxwJkoA3O9kLFJ+
T0m3pnk9YJbEpoaEmnzYKkmSRn/dInL4NMU0f3FWtKxSW37gxm6yaiaxnqlQq+ebNjMLBulPQrn7
74ait8TJ6ixlod+IKXgfeyZJtJ4sDui1PxFevV8xBZpQYzvhMXM48yrSw7mZ38iZuGhg93qObDTd
aDbJb8etxPU8u77glG9AFUMDDmyBk4KPEbAS+LhI3jmEX6FAg+pgFF6dufnM4Sat/aeIjCeqEmTC
Me38ZWDW48+Dac841ZdEqMw5Kcr0yGguPVT8qqGyeTjjEoiZ4po0LMfwfEl97aP2wZLgymIfer5Q
ubfzzSM7pnTu5dlOT6BqEV0l/Dczbbo/AP+xA4e8Szc34rLLn5H7O0GywektfSSVvUr2/9RtczXy
heFD7VpSTQB1PED0T7stcWRzlhVYmXlKUR/ep/1OxwBhTwo4qcSfrosSFGgykw+fhH5EvC9tVPOy
OIM23g5xXak9TlFVYwuso1nIZn/Oouy/UnwWJw7MLw+EUg9MXo3KBQmPNXqCAGwXPGnNmyo0CXI2
0XQZxpU7Lgq5VLtAkUaLRvZS4N1WxjZDpSpIv9wJLUfcf2VWhwIz9zZnaJpop470nQCy2n6EtdHj
BjwmFm/sHsPaJact3TT9qNicA0iw2SYKw186yIiSZFPsV2+YMbagf5wSMeR1UltIVbHeTMWqiYXU
qqiUGKEhpuW+AalIzceJEY97XXGBMzQx5rNfkC0xosECZFzFmywng7hWYkl0iUishBlHQ65nqy56
9PqCQLcaQe+Beh71KN0x/DWYyEuqtLzFzmktVVoeyWH7dsk4+RenDeA8NE8pUoems/0GdIcfidSb
+7Ge6/HVkSwjg3sGcNGgJOqAFAsSdF8rI3FV6n9bJZ+8cb+BG9FdExcQP8fjB2t9hokjR7CC9JoQ
ER6KIG6QeaGKOeuh9L3rg/oe4S4LfLu+qBm0zckepoGY5DQ87/Hew/HouWJT2fNVRQJ22cQzquKu
NSY4SiCiQwWs0uu8wdLy1HoprEKZWy29QAhmKYocCjZL6D4GdwDgGJ8v6F8o3uzOsxTMtHTHnY5d
+Uas/FxpkUO2WpWJ19DfsWyIInFOLWoYMFikIBrk+J4bYYlFiraaNzHDmUzoiaGPIB+07u/JESQ1
s/WR/PgOelgVeL0wauVdnQHVy8Kf2vvVhQEOddp0W5sq665F/V0C7TguRe8DLXcPsC02TM4DskRH
HRVd9rM6aHfRJCCr/HTScLUQK+uo6ShMgWxnLfD9KDM/xXZqcP+/H6eYY12hghpgsQFPA/YaXJTe
wY1Lcjqpb/6kXDjsWjrVWsqkmoIXEa3xkUMCOzBY/T02FBtYGNinH5ud1DFY5tScNUg7w+X+9J8L
AUm3/u6j4P6I/Pdze0QOzm5AfoVEHa8A1bICVnT+4DSdx9Ni0E//ToJslC9ScrnSjFa98CxGlRR8
F5NLyxS6BImrmMwWpzTZDxyS5U2g6+LJXLZGTqrH8UhqC4ndOCbtUWNSp3dIJVsd0GzRgpRvTC0t
DJvcq4ZZjFV1XvgGctOHA0fV2kCZY5LDx6qbeBIExxZZYs6wowdQkF4OuM9ezkYuzlDCI7OjJ6a/
JojGE/5ycBg36eS7JVtwIS8EeTXIPY7dJvTPylhCoA4K0U7kU2xoprB8pSmlWvQY1iUm/GJ04Di+
uqr4+lKQtrfCCudjtQ4X7tWDCuBvpJY8YMw4+zN6KszIGNAJ2KY4X+1JwXphiCpQQUrcPd1jhb7+
3bO3Dy0GkRdLMFllxhWaji1KkxalsFjTL7qsUE1fOgP2iQKLTf0lQRL6Eamcyc7cAC7Sm5IkMMXw
FH6ds9mdSLz15LJmOjwtJLZKeJeP7eo9NInogiiV1HHl5jDgBP4mOZ0+f8UWWS2x2nOJOowtx6L6
PqqLbLHzr41ToSvTFZTt+uKrNOL85p39Ze6lB49tyz9OpePrPBOCEFu2ATQRrLH7iz6hlcBJjUd0
k5f5sKQoMJyYzaLoicFEKtwWCoO5ccoQlWkVIli0LUBLBnGBZtRGzbp4J4tdyxNu9X842IrkkXQV
Jm6jq0b1ZfgRi/sBjhmXB8NH9bZ2lTYNyFWyUyZPVukQfTrOo01TTiIQQEpI4MnVTy4XrEvxiixH
Jb3WExJZsDnZ6StNt/YaNM/G5O7mBbFT2itklNXaLUcGKP217PZltTVfT3KIOj+tAai3X39HwSQC
0BkeNVWDmTi6D7pyWU/Fu5TTpuoSVTQU7To8omIUsZzWsf0L3L1uE/D1CAe4XI0fAt1gPC0RhQsC
px/le0KWu4nQD1w85hxcUiDmmRF1IE5EcsuToy6DJ54CQt/Aymm51SG+3fp8/fosXSzGfR0e4xpr
xHkAYdl02nQf0esovKBx/pz/X04THKx+HyemXR+8xue5sTKxXlvaLbHh9KOjRqOWBxiiKMz4JsEj
BkgAtUIzeuyytXNB9Jy1ct2gDzatqHjeGKYkY07vZsfZh1wN5oUM6pq3/0vbJ8IEPtrAvW483NaU
udP723F7lRC1MUdPSmSNHDF3rn0EB2LJB4KPISckKkXTtzUAuYHb1bIvSQwPLPT6ya7qDYhS4pzD
+2I2dkqDnCdq3rUlaoDipEsLu4B5pl1upVOm2uQkGaEarKQkAmyUXXzDE85krA2shZ/8xjC2WjQK
GRxsYr8EkAut2beewL7snl7XE3YEHw34ytIwHRlUTrJP8I9aFMaWGj76kyJfm4kmcm099ybRApXy
EDPQ30F8rMFy7DAKfw4drIWhvCJMF5BbCNQlHo1jWrTsY6L71AeEh0xrEujzOQpP9/WHW6z1Hb4z
VekmbM7Ux/tNwUewOaAmSANcAZ4ch7mGqcRLs/XbZN/x4thcUlsXtJXpzWFeCes0ABwPsA1pi7ZX
ur/VpD7DvskjWLCLNeukdvNzP9ttak1lg1A2n0dK8EnwpATGsxwfy8dqkZU3LudiNTfStzGzH3y9
RsElm7XHKzjcZvF/W48Y2lOsVY8x7hy43OWOQsDLATXh8aRTXQMiwQWSfC+2Kb1+GRNThkSr/Cn0
D0Eu8bzxqQADSZMxyyLPDO2hcMgZUK2Xos/zxppeuALYrkK4Vn2lFOKxn798J/DaWspRonkjiA5s
pCChy+ayhP8Eb7yHkD1xvsOtwggVIc4mzN8joTFM6ujByuZJUm6K5jNUtXrJ6Zq1DxIeyuDNbc67
yLWI+mH5HR2m/TcUiZAjCX6jABOOyDQ3sSpuShaF2NJVowAUMQTT4Jm4ANwbhYNHz6t69LcJwHZq
WpeSJbnQ9JfoPY3gcmfkpmEDSCEapA5ISIGkLdigs3zvNL1BhDxFzme5Nvm11+JGn4lejkN+tC9B
m9l3kBNYTx+pWGf64W0D6Fo71Tl0sygChKLG2mhTfe5JZV3BU4b60aUVf/8hU5OfCWMqzv8CxXeX
BLCnXRwne2cg4CrWm5rw3NU++TjrvkDTAbu3DWzu2mtPrcGyfj8fzHDnwmBBGl4Ep37vnzSg/NDl
HcQqQDESZtDqw8NlB5O50dnW9BngJ2DMlj/GYGz+2OR6B/Mx9zPR57QXH5sQL7iH2h+YGWiHfVNt
kFZEj4zrPxIbE+X/hYg3HNwp0PR3cnBaBWKo/Q+zxWo+lnzdWmoiPqdaP8+EW9R9qmvbowyI1i3O
pZ0cw2t7VXq4YSwvvzZb8aW/AJIFXfqVV/tUn7/zwcOf4dpb9Uwg3VjoBOUBMggnL7KSDEk9puwO
59egStJc1wYOagPCf/4YcmJ/OTj5SBMnfJS6GkpieifKhJpXnXNVL5HEhOkouxXa0GIgVVqGBKXY
SQadiV+Y+CrItZSND+h90KJHWgvQA5Ns2tzSOD4Sv3OERQfEhdo8FJ2GH077oSgFZIQwqFRaCn1T
sCvgqrcKZXrwtISs6US20qcgYZjh43PLrQTZhc4PRcnE3sfGte7W83qOzy1RoPkJWWMD79sS0wNS
Px4gq5lnMMfXmxPkPy7/18fQ85JwqqZle2z08sjfTw50ECt1KN3LhGFg0kFoV3Gwj1FUef9vUeq2
aH35kUbSfKZzSuAdDsqM4r0Q88wg/CE5ln4FtuDVN2mzuxaZlg6gEVtYX+eGDAKVrmqyyvRfxcJx
uPOvak0k9/0SiqaaKEqhOv+6XEnG57nd4B+fz6g9iAa8CTxD5rsmJMCQaqKLqwN3MA+NYiHl5l9b
ppQbnEjOTcPJ3sadGs9lgjTZsT6B2kcmFC/6gLdXFadPP+++8rU00SJRNuLxhEAG2FIh6l+6JoNs
ReMq7mBIZSCgHXuIVB8LDtw47qN++yAoCVBJsAenQFMv5nDYSudZtkzUGr82DGcSVhW3GaVbBOgM
QNG6SkTr24XxmyxQiccPOUsUNUxoI67izJiqAA2kik2gPTSShVY/J5NfR+g2fnhzKyTlpcTD2cBX
t+/k1yNFlCyN85X0kKH6k3a3vIv+XTLdFq5J9OLBshf9ZDlHoYiB6rU1uNjf4IgBIGzNglh4kIdY
IGG/KGIgJonHSUOIYLIjf5OpWs/MpIALr7AvtlH04oOTFPWbd4xXfnokU+F2NGpgIyfXkU0i69LU
VoM2HqgcKh+VZ7YBTsV0DbwhXGZ+vggiFCXqB8g1XgmTxT3zqozPzFjdUAFM38rVSOhkWifF5RWW
bFJjbuBMHZSuyJzjP9EXmpKg9b0AYrv94mYvmo18efdLL3bvS5SIt59kWX6Epf1d58H6NrBHXTgV
O15ibvVHpbzUfXEYA7st4LgcqkrukhxEetS7afA74DJlmJNHxkvD8lVw0xkyfBpphrZjKON0lFWh
4NNnwWlAOVyfvfdN/tvQepo0FLhd592dSaaZ7XOSoPGfgHc3YNd8iMnJYm+D4zhdnM0Lu4ER9mdP
64V68QzCVUYXq6HW17I4oQI1wM+lc5k7Rwl1Bg3sY82KqJ8Uq7kViNCOm+6mKqCxAbwhUt7rPxuC
UZweid+78XFwOEyQNOUK0kaMq6F4FhiHzgSyEyHuBSN/QqPJEXZ/Kuvf3OZOf7fuE8BtheEuwMwT
APqUlhil52KP6bWW1BcMCGHr7KfDkMOKXfmmfiEdaC8h6Qa4RZRSDoxJMTKj1NVVCn4d1s1r+hfw
JjrSsW29CmOH3sK4sWPSqR4m8LrNj6gDyfAmO+w6DGr9NvLYT1EmE1JbO3ds2u2+yIpQCxTrZMuS
ec/SPOv/Gpty51U9qmCpv21uw39tjnrNXjFBSfBuAfy9JU2iiokNj5Q7+Bpa06yKRqXqNlKOeWHI
8e/2iSFkICqIJqD1PBu/ad5K8PXjYkpRa1wZ/wT6N9QURRpY3WTkJzdtlsGRDxuWfb4IrjFSHncU
s77pc8alniAl/bEwwCkpElIBls4S90gK8W9VumkV6bAKrpnm1+5ZEva8ADO5dF7uLYKtHG0KemBe
2/Me3OVxAbXsJwsziJy0gucXXqsLxF66/iBZ647DJJybOWHa+/MT9lAzPfpj99+aRplpy1uBuLmg
EsO1nrn5dvN7paoXNl7YjIfEYlU6+IH+GxRU45Mr7kvCAPW8ozWV4edW4u6OzZmE5oFTMED7CPQA
kq4TuaBQ9T17xZ3fqBXyxQYywHnAREr4SDXsplXb6Dz3Mn8blFoPvC+GYenHEgULM8PJjo9ywlJ3
BZ8L+YtC4hlDJjm0oCsYEanlJJCjLDxNGrDPpTtCwkHjwCUz3xlUu2hNWfPwZnk17i2y30OIpBYd
2VuDP+IFjzoMHHC0cst/5jQI07hkcXAhxXkGZ39BVRVG+9+WFgX2T5q8xKnSDJ6UJYTEmmcEshT9
0KgRmj4D7LBow8VnRvmOsT7F/nCH6OeS5OwdWcVdMiNBsBDTaU0ubB/K3KfwTjTbr9cYZJtja5M7
9phifG5MVQCIj7TUYv8nwYKq3zWHA4lYZ9+CD0V6yX+azrRTyO7zO7AAGy6o/G0TVhRqu6ouLWyW
5geaNDEm7znOlR/UFBaNG08UYUb4NLbLJDvGAHfxkaXWaDkNF1dU4D6UlbUOzEE0H9kqMXAxGavl
C9qfkttjcl1CuB2WOggJvLvyvujfhANaZdwg2OXk7MsNj34jGSE3dl1PYqRnSK38pkLkojhBPbEL
wJoamcmlWMWDoksuWswg4vkD2SS1TpNpfGZk4hrT8+kcQBcgjSzMykRHLxi9fZbyaFEn4HIvJMbj
5i9oE6zTnqwqWYUeR1uNCjkksQqZ4Z8jJRQbwAzQqv4l4Rj1+zk++ZZw9Pcd0WH46g88/aHzChQG
zyVnws3m2Y93U4iU9nTXbKX2cY2DCNS/Q3ri17UASKBWQ+3eOCGUf+AB37K4WxLsHdgIlwLfBjx5
C6qDgJF9aIsguRNrCwF6B+moNkFxFAV3gx9PpQa9FNU2CezXYt7lCeqZ31uWizpwstfrnaBwmBy5
m3h3vg4YTFnJFxakua8Sg+goFHTCBx9LtBqndgDsLsYdCWp/J7UJmWlbYKLWmluMuOvUsaHb/CJP
xehIBV1j2Nb2PPplNuKLFWu8a/2ANGBB/t+tYChzfF3y7BOPy+VZXIvrHHvmd89Ym6oBsIGG5edc
xooDjIlI5dP5uDo5hjA30G/+U2dceUH7gIJPz0HV4zJ0RyJqPQXWko5SfHNGZqBaZFgWjL9i4PuD
9jEUvvlbePZnDlB8f6dBlog63HWVNPvnLr8BFo8DMh1MGVmDYVAQFbggRC9XyR2vHSvW1EGPF7eR
CU1pMfLUJ5tESiH15FEGi7N3ADt0nLdrO9UqSIJVH7JIfbHCriuCmQfKblCQ+u92dW9FrZ5q/Mv3
A/t2SdhcI6O13e5Zs4rcsgwVb9UyhmIXIdVVMaMSgrUSURFpePrL8N2bH3wjnIqrFNZYe/T7PvO6
UlUiG9mnK7TobT59FAIl8Ru3qrFKTd+JGgW3iRrpg28rL61WW8GAxe8CE3V0R+t8b50BG8FF4YYG
uPPu0iSffftF7e0BE5zhmA6dPqWqNPhIXvvnEOSfBoVu98kDYKZF3efFSlKMdlQ5pOXkC3svd6xy
QJ+Ccll2tjUZVbiva4P95pnlV23jDL2Kr6pwRzArrjgUXp0JPXnyQfj27upHrFf2OHdrIC1+eEpF
x3/oPUx8nEP6wX4kO+T6nVSRxND6ggaeTqDU+lijCHP1RbQWdJwcWcQJeVeWddMhTP2KpuX8QaGF
HfAMcNI/QDIi2glJccv0pnQbWuhiy7VWn3NJjeMIHbrr17GP8Hza/dJLBtgtMcDwoBndZItSsPRA
BsNxrqi11H4MRQigkK5zT0dX2bl36mNewJg7lcw7o/iWSN1VjnzsE61gEqTHTh+ssSF+ZDGMWLIK
MvgQJ7SMNPVzjbLCNmpLfpA83xZu39t3A2a7re4VvExCsCXEZqasuFBls7yk8JdDjMpRrCJJZhk4
gPYraCJQSZi2yYHkG0ryavw6EavCDkGrxSWKGtxMw4LoiEs9dO/v7npWKGnDDORAQ48VJLk6kJKb
VT3O34nl/ET4oAeyWEQBja/2S0KKFlqb05s33RwoFTBjrbQPpLALQEisb+ttT0pqei/ALZrzO84i
q+K0yjPqcfRBU4E8DPD9zvdHsBnGYAAXohkju0CacT+dL/FFh0npXdXZTSF9VwkiWfIt0rIdX0B8
G+vWs8iuA2ufhckv4b6K17rVNGXjhLJny7s1p6uByC+aKYMeV4/WzrCp8Y+scYkwMWg1xipvz4Z9
gg8EoJKWmUsGbGjvJkmBloApzv+euO2M8eXlsT9O/5GUr7ie/IUGL5AB2rsoV3uuZdIYlkemhu5d
/smvX1s9LATpiRCD+fMFb0G+0mOjmIDSsozZycGFxYOHgvUDiF8EWLw18tTjXGcSVltN+9G2sjBK
2KUjQeJ/yEhe+qk89X3JS52WbtJbJuZOUT75ID9PpK+QpSU26DNOqCp7G/7qGGWONnvrU4aGHH31
BXdPqogssOW5o7KGNvR6awzoBOabrqLpBn6YiOQFqL8VigE9Ep3MB5SwkZMFbHrSCSXvfdvNiJnC
w8WhyR2FIJ4amTBokGip2cMyLIVaCkxrN3GseH9jpwq/Kaxew4llDlbFSt4muT0mOY2fZu1n3WTQ
L6CDzbg8njXOSC/nhylCrDcJs67Iw9AsetEfhgYO9ois73uzHq1vwXGE4MkmOZAwRHK/NVkQSmah
AthmCYdQckNp7GgjsOKKfu3YZ5TBdY5BR+++9+epgjP6cNAvV1zk5FmK58e/7ll8EZo66gUlTvTc
DSemR49okVdY1G/39T7pfr0lXJ45TOQoIgtanozwLJV4vjDiAPSqXc/oFQukQUZHUanbE7aUvuDX
E63c67hu8+HNT1AyaBzgY5hvItyoLfK+suADz9eA0iTze8EsDEmuGrSCm197TGTywIjzWmN3VSgl
3dGDDejQFEKasPiDox/SkMoCso/6437cBZWvZXuyaogvmNl1Caj6UgnGU3sBpTzin55Mr3MNxvon
uA0oMbJIPVFVqEm850c1CJah7qUFXba2s8W0NXtiCSvnURZPgPzcl4Rj5y+QjDmpbaxPh+/hxRQz
q0ESa8Ev/vpCKET1gShUVNiWRuX/7Wu8J30ZHbANxot9NxKW9uu/P74dm5/6mXpUernXw+VbNSIY
CJz6VdsTxrV7IpB+J7USsLREvURSwmmGHJw7c+jruuF8OzWFkXvnRmSvaaEC44M1iUBQbjgTXNTz
55hyWBXKKrNYyUe/BgO26858hYfJGdjknFnavPM3Qrg4yfcF9nZFCXeXTqqs5e6oCwVO4Rzdei1k
ccACBoDvA9/+a2bbpIhwNHfOtteU1pE9SJf9TNcqRXXgNAYZOLN4VKZmI7Vp+Bnw95xYDHThvFWL
sSGWWN3R9NAXmkxR1TGwuzSRAAYPFfbS39M+FtwG3hBTGNSA1V4ZBYg6mRhZ+ZiTHJQoydCwEnKQ
C4hqzLGqUlm1IMCMa+YiqLZXjSmT7XcvAnhfdrElJJKyiIcgqWjC3DgDIApugMgP0TQt47xhq+ib
kuJxyTKQou4GV6R5GIH5VafXMRhD/xSneh9FDkIc2/qTevbvqPrJKK47UXgKKN2xsry3ezBQy1vA
DLcKWg5OZ2njd9Dw4tmPwdIdKyGp/bzPDNQyapvR9cJ8HPbzcyjuNEnu3AWq0hhzaPUdgdyJDJBq
71bpkVt4BaUAFa8ggKvVI0fPUzsxaZ1WdwHA5ur0f/c3TaQnrCHonw/kQjDsNCkJ+MIsC33ba88k
kSg1qQypRqQmzBQxC3xEBZiaOBA+9xP4NJ4gxF4uNFApFdhjZWJyVo2neODjoCtmp+OowrU7UsVV
FeWX2tGaVpVqqVC0Wd7FeC+8LuMleZymi6Gg6cbSYIky6wC9//ISPm0c3pNt5MSJ2GJFyn37bVf4
xjOEAcavyxhhgqUrW1p+NjUW9Hld0+W7ozcA0trBLaZPW5ZI3SbY4vOaiKy0XXH4oF09j4DnBHgT
XDkn0lwKMwiRH6J8FbKjP9l0uPZD41TT9TgBG9vLHBxSswS6q8VJAPGzoxcuDfiGjYM7u45Rlg+/
AUYYlSSdq2jwn8izP/0cLuVfuRe+g6rRdn7r1+Euq7esPlSkbxkc0X6xkNmVOSCgi0NwBVYtVjIR
P6xZwtVskPmvFaDKGt83BgZ9lURLLSFzha+2xemuYSKz1O/pvi6KU0S/ywyX0Mfc6UchRc/DTRuA
v1OI5MsD/Z/5Krum2PAlZtatrytlmOJ5JeswPiNDNgQb/hrda4kLuvVDrqRg5qzm3O3XQSzP2Js3
LlxT0+UCmamZ9rnT00IagzTxHSjbwpPVe7jf63G8sZH/uZcEDyrdDq9j5rUi1Vzyr84ro/9pxXlh
iW+GCIY05ksMZZvdFuZsORJSCwHj4nSabwbFW6vHon79A3rxTQSI8MrlEcypA1111XiXQMIzeDuk
BWz5t3NIY9Ss+8TpaxkAicIps46eP1w9RzA6Nrh6j37TMH2E1hVvkKqqn0dGqI2klhEsPZXPl9rk
6h9hL+EIMFSpS4bHwdTFrvo09v771y1DEykcRXTcSCttcUyw7XULF4cWarudsmbmlzDsakxufHI/
ixE5isnD5EWl+o1tTl1/ryuHfGVi4MMpl59GOfTorfeoo8lIne21s78YbWXZ7TRhx5wbDJgVGv5J
jfxkES2abdOt0u27sGyEvI/STveEVJGenBezQb2jLjD5TC4sGCZElrVXChv+6m0nMb53wV3czZMG
glWRCZfIvFcv0sOyve15GKnzJ3ja0ePBAdRFw9n2TKaFa2ZkpbfMu8M+/1MdxjnWGzRXls6TrMA5
CzA1YWx4MEXMBELdSFpMPpiUaF9UmYcLqCdhCPIGsTavtM7vTJdnhnSZ7I36jwvh5zrlsglSAVCq
yufZGce5Xg9cWbwc8zDWpK93B0B4xi/ygIs9NcXdxh9FpVFKSi1eLRNgmT4wwtv37cHpSuDlN32P
SKrlW6fZ1eAqgDBZgwrnWL5mM3Gcb3c+5S+Z/BVYNl7Zw4ESo0AdWGpqXdGYJsXBb9X4E+zIqRs1
C+qWz05DqscpbACIbh1WdPbwO9yBQcnpu6cgen+AnK7aKrqBsei1hEe1EybXOL4bkAQcmKCnWdUE
XjpWy0/dJJmFwpMSQjQuq1yCx8vpvgww0505g/Drxe2YZzfyJROqUq9k4gUWR6LL/GYO2nFFPPcD
j2IC9YUEUmGCkoaGg2SA1L1ufgIrxmqVz4jiZyP32m5n/2KlJgTEntcFG2e3jTyZdNI7U09ct5up
9fpYsIlE3iFqmrYcLdoCBg+q+N3GcKBPMUEvTNyJ/jrjlaUZlayoVkEcbMvE8fLKpBQG9eht8Twg
wa0/npnNxvOUA66TImtZNdh7amYnEWDKqSwETUJbNs+RKw0iUejP/izsOrySxbew3ICTyuQG6rMg
N/ZMhKzrc0Ge6NpqvyIr97yMawxVotmROse79NtWKzUEOTEFGjAnE3moPYqkqfYRMB9Yb753/ptg
l2apvsltYJT2F+VdvlYgz41t8N1ehbJ3n0Qj2AaH7yJS27j8ysw+s8Y4Y9J5LsztidujuXLRWKnm
BYFRc1luiOwRLBsBBTuAZC6gNutEzSpgRazf2jSZSfrT5iF82azrQZgdOEk1X2HVa8o2TIrtWhsM
a+m8/MxejD5q1vlyGu/0Cv66Yz6xCr0WEABRlU7gmUtDvMHuGCwypHoRtiL/J+eLC/bdn89uj9Gn
vu/5I5LorBXPHiw/FOaQcgdmuuysWDk8FCzttUgy5zgfvV3EmaPS/0ladZUMS9Iq3QTc1mE6dTf0
QCTQu+KRj3tCDrKWyFpGDp7tNFL17sopGvUbqJWvm3CtfKpiNJkp48/ASXzQYntLqqULRdM0kzxm
BRCHjQ+2VZFg/CvjgiaiXlViQleoE3j5ARewdGX0gfh77ZwzYNbIy4i/RZ71Gb9tmfoStdw2/1gv
9fC7at8zkPxPWqBw6azL7AmILomh/R89XfWEhc3k3vXRsPvj4miFPdrDELk//TxOTysAR74CYUhM
QhhEMDcUNPBOPl1W52F8aKoUcYG4Fa4hkwzoGxpbJBtMoGeadOtI2k6WxETStJvTseNVjkU78ZH0
DLreM48KaoAc2lt3wECwzX/8tsRai9gaa7ANyg4haquRj8skmSbVvDR62hjJaPYXocXEy0z1GadY
x753eshCUIT+SRl2pQX8GmV6qrEKJwQf/wMG4KpZWfzOzYKGSq2k3qiDBM5ziGB3ub8Rx2KzFGtk
oZDaJ+lNEXTDcynwOatm2m30Tvr0gw1patOOmcVY7l38tYNMWSTcbEnRU14karK1p1nRk8xhqQMD
Ko87OZnatn7HEHCBTdN4C4UlDLc0c8xbNX/9QLkKpbfxmvVncVh1tN98JTQ5B6aI0C7lJYBKTkpw
J6Jc8OU68q7mT2g7rH+2d5fRuA+LW5GwBl5KwsTOfznWzfNv6fH2DgNzJL2MUnd6KrIfFJWZYjVM
WTiZLy6aV+mh0s6yTB3xkmipRMPUrF10pAi7uh8Hix2WiQolnGqb6anhig+h+gh+8HBOFTFHA1a0
35X64us9FMlLbV23DFKFHsnK3MEvMzomgYC0h4ZHVSIObafnpfiFQWChlq8lK8kj6+LSUez/BiPN
fwcn2lbRUNAY1EGxMcwgIjm7+Vi6A9OwU5vE6sO439/875v92y/sJCjrW0DueBt7WsWal7xoIVpG
tt0+nodxjRivN3gxqZ4tJAdCmlHzpNR/aevksMZWc8ousvyilM2dBGcTHH0k9OV3SDQ+izKrO7v4
zk2Z7NnmisR8F38Xd/PWmY2ql5RWeNyRyIYYXCqIqdETZMzkOalcI4IXm1XBd/U3gGVuMjhz2l7J
vzRYhoJpKWCldB2UaYx79cC1UwVr7jB+R3loDxHavpfIzAiRlDSEiif260QNu2UqQlA4X+3T4yhE
wrOHcixaoHz9AoZlLLJTgaT9kZQeUjct3zcTNxEBTc2EkghfvQKrtKOVcMFlZhut/M8fAnH1rluz
I3D4neRKjcSZyZZc1JzjrfTa3KDnLgi0drLs74KXN2EgmUvlP1UvTJ7aiz8W5qslgym1uG5NGxOB
+huF9IO3VLYDiOHmERMdZ6bNnxU9FWVnetwu+nga/1Bh3REIK3L8FRu/SVSSQSmE0kjNBTYJu+Dj
IxCl8489cHNBJnXtOpYmFgTftac5pmVpwkaR55vyTvz9TSwn8IVhoTi1voAck6buSMM6No0xCL0g
NyXKX7pvDS3oIP8iqDRaXZw0mzkyOX0a6JD55v0NIQRCZMl1GJLxsG3qn9MwYJzwzqkCrz8UZ8WL
k+hU5mGqDmt0Jh/qccRqojAKNLtOkLkPUqmbUg/4+nKVupKU0fJdtNxnG4dsYSW1Gq2WT7ycf990
7l/uDrO/ik6JCbfDSyF1uFHDeChEU4RQ0sG2xqAlO6MMOb+NgqtRDtB/Nxu/Ga9G0mdUis+9dpmo
StaaSXdbIbCBx+8HBh/JIS2lydTNo9NXn9bpN6hDF7+GHEG98Ncs5TT9//AC+jx3etF8gwgv8Zs5
l9v51gRZIUzgM5IXcRCXLhQrh3SNPK8of79QMugrioua4Jwm3B6JYOzUhckyLxHcSUVlTfGuLPiO
jsGLV2hh0jqMO00G3HFEoUUW0VLOEzYW+0EPwLKN5OS6+OAee0mZldEX732DYvp9LqmYchFsiCBk
/pHVP3Rvya1MNw1+s5BpS6Zi4W/qM5Alw/deZFsUgIKAyyfMcaLnxvI8RqwpH36JqG27Y1yVVhzZ
jCOLFg5ZGQ3cwrafqcyHv8c/kMVJ4BB6TInE4MuQvGMV3fepc0vux4fxYdr82ytdXSkpU11sLoD0
RTdIF8/BOkOUI/ROZtDSK8rVG1kqag94UamQaj2Eeb8VTXkn0ebp87ZbV2Xz2V3GZNesMJuBCyUW
C7pI5bUiI4GqYrxEI5+Enk9lHCLY+TP8AmDsSGc1MzoJYYefy6Q+C+Ls43LzIu8GHKWQ7rEisAch
Ei9liqxV+2Kysfx9wTy/fxrGJtYoBSArZAQCByMeUXyfB89HKUsOiBHS+Yv/IyPtvtAB4jPqwI29
+x45+VnbNvZz8FLeUAHEv0HKHbkB26OvkPbCm4Pa77Z2piEII7WhEzZHfWiBf0s9LbWO99gIiocE
arefSW7uZLfShBS5apU4nSlO6e1pOCvWWc8P6G3/R9JZZuJ+1cck1aA5SpkajIPxLdSIAwtYBqKO
NniIC5x/YMYO/9hrLCurFcUoUzSV64YQOD5tQG4LaVX4sb5VTW++rLprmWmIM05l6WgYX/1i2JTP
OviPu3GWfHxV3sxAT2J1212QZ7u29R1ExamK9Cp5hsyr86nlaTuXH6kefNlVs7/7XAt2bnfBQ2Vs
TR3VAkKDe+IriHFeDjRY4G7XCDw3rA9dsf7oCRkmlJYpwbiRc5sz7oKDS6MgMIAcVQe4uqEJHc9v
XVoroHcK2bTqO1elIYUNquEI75JYjAmAjz0uqluGwizskFTsXpz5S2i8J0ujg+KS9eeltXbop/kN
wVe5aVKPhCsTwpjnjp0hX2N/AJ+Ca55sTkcz1mkNYiwwvVRyUkLCRikYOK5BIzWgW8TgKdHO0DO1
4JxfJdACi+JyQlaot01vU4w7QjqZtrpOFDPW71Qh6PZUGdZP4oLAyK4RSGTZEksQSTm0ZdLQ87Vb
nfmfMbyEx0ihoRAtYLSlpNBYsuwyh9qGAT/8AuLdMAAWbsNJl1RA5FIdpIohPy2Qa02N2aYq7dlU
gt2SCI15BQm3ezFTL4Rze119eVrrA2cC12Z6jy1sS/HU7+XWroA7uHYauR9V4cXG2s2OC5tW4cVB
5MkoaWKXDyevH1RYdDJXVF4tyJvJUvGvigLN+2k3aqgOoCAypKvmnYMAILXYjR+1G6qoqcfFfFoU
wJJOALQh3G6bOqCjetsrIPaMNfJqn5cxy0FmokWm6GicRyI3LGID7dcgKSs3JUIkjvIUnVTsz+xv
hdD09eE+txwa43q1/G2yIRlpLKy0FWSoPuwDrIOucyg2IjPc5xt7qhmmbrPe9pnDp5LQqJ60WjSH
1tGU/dbv/NxXX89n2stF1Zw5n5oZEUbqEPVlTbilRbl3hXklFEM4s10wGPj+anA0LUh8nDIAHzyU
ngWOvzOdV+FbH132PL4ma/6L0gHD/wZqYJffznjY5E/W9PQtEiqc/wlOpJ1RtlKFuLaxdud9ddhc
u3K2RCAL6xbI87zpsVtrBR3r8U7Jrs+J6fJu6SgG3x5SMXLbNazAAo6OKCcTAKUz8FRNy5yhPjcG
mEswEGmtSeblIlAma+czCES318w91NQeZE/0a+CROVbXPgbvbyOYNO/OQtEr1cjhPsl5oFlnRWRh
HT3BCYNN0nHk6IijGz9Y/JTjEePMU1YcdU0ZuH20cYa76DeXMRnb5mviOp2qSO63jnRf5Jl7/OOu
D1jWjE+9zIDawSUiDcVrsldkUgbsNNiqaBD8jhGW3npuYQhuPdPG1Cj9n6bEtpNM110usP2apsdP
67hbj5KnVMwyLua1qlHqbMS7nrdMcMC6RW1oRnAc0tKBjW2zvVEDMuyDAVG2FuroUJqAu2fl4ayJ
xdTbXKoJa7FgvZ4kuBeUZmtuVRwJo6V6V6ugxcpiPrz7Qs6Ry7spGl+TjBqX9k9U7jTrIQW9+hRB
EHBC1LfwrZANM74oG0/5Ts5VIO3eUWfAfyPnqUNus2MBH8qTuPcwhrugakBtvZboysRpsnm6JyJf
RI6SdIf6OZti07G9VP2oNtdaRrhLYvmfSZu5KpcY+75/+msJgr2yWT3Q5+nzyMgA7FdRZCuka63a
/dN2aoogO/hFaRnIjwLQv53NgPMVGt/0hDM3hJIN8Z7ZMoAlXNKDF9fCX5+fL0sAsKx35lG6I54g
RlEQ2UDHtq4SvjvGKDIOEIxJbIKW/D8HM22G0/XXSqWer6viHt7t+FURwDG/6ar3MXhsDYbKg3dh
4/9KJHHfmna5hRZEIbbXXog+qRRs+f0SoEj40VPWwawjxH/fSwZhz5jaM1mfz+hRD9ZH6Go2Dcj0
RGMae1fFvC2xtooUYGg6+FabeeRokD/gWKwWGnfDuTK/waAgJ6B1AfOvly/LOqcYPoib6HILHNRR
JDjyszPRYU4XltLG3SCFPsXeMlqfaCpBze0O6e/N6IObAeAmBu+nXG7N13mjsYMdDmjvp/dv732R
CHUNJr2UOSYf6mnXU5JcY13Rj507xGbObiMdpDaFq62WTZEC8BFV5SWYlwYf1cmcuzxlCPC/OBIw
m7bQa/QrTTV2LDcZgAUnXE8+hwpUlKPww3uMSVZfywzM0kOZxjrLKPdnNCPLLIOeCmPVPwDo6Jzt
23ck2Zdhw2qW1QBp7huaIQnGfh0KnM935NqLg0cCWeRCO9rjB/qW5DNVQtNBKtNHde2ZjI7RHreq
f4oZPKWxTWMPNREjP/Rv6jMxcWB9lkJSZ38G+OZwNd17gB95CP2WnsryQS8iveTC/7FMozFQAHKh
dNWQzHwGpIv2Y1y2q/XghNei5m9M2Vi6dBrSt9Vx3joUti+N7+tFnuDUIk4tWIKNp5/VJOzD8KEA
KvMXs7a233hwDffXkxjaQE3fOJhBurJ6cAB76GSS0Mj1aITPLlelE7ThAkELNVUIBt8sI9BRQY9o
5AQkGmgjn716cNdJoL5zKYDpfHi7VW44VD87d6g66et+aAjj61Mbm3c8aN8zfhnmve7fcPeF6kAX
zuhFiEwQsCp0oNjJ2vz77rvI6wNHeakVSKc6wbDQ0DDSS0zSLT1N/m1GgOZlmP7kbY89UWvldwKC
EgcHFQ22gj2kt3YeK9Jk6rnH4aWd23YoSVDIyPACLNiHJjk6a7Yi8p9C6dBV1WcvL8F0Hpkrr9Ec
yW6Bmg6lrTb1Xu6FAN51/9rOMlmNoCmdXj58tjLGuGiAuQQpCaFCmzyspvoJ7TESr5KfNx7ebB1U
aLnZvp5r2RFFpKTvSrM8ttuJ/UgXaHwZ1DAqmUIdQ3QB1ocwLfVYe+ROLGP5IzgwvEtmwTy2ZCMI
1GvrJl6cXuMiIQ2kljuuRopLdxE8UB613vh0F0YQqFsEeXqAUuMHNOXUnHvvBGssw6IS/UTLAPvd
IjkEXEoW/LmyfzBZxwO90lnScwsVEys4yyb2MHSYsgIOAQJWBAdHj19np6HKIJ+JEVH7hn0gMI5D
zlvIJFWoDRAHfXFdNNSISR2MJx7ZjToZIphQRb4VEMhl+XHs7wYGzkDFPmuv7EZhJqbcr9dYzhLg
zLYYVdvBp6zqbg4nvFtKe4LkOdlOeOtseFy0/Toq+GUj+/XKg9fTbq9Rc/OWcYgEGO4oK390rFXp
f5dqpTX3BSZNcJozHoe8cag+xfBezTYdm0v/WKcBDqFp0hG+pE7sIhoEpq7wK9rNPnJldD2xQB0u
7uG6Mxky7uv5/q5OmBJ/cgQWzSObltYd25G/dMXdoPqZtT4Sx6Bsfd6PhRoiWs0d9xuVzbhB9YS3
Oy2+nzrfbnWy8h6IukFa4wgJQJFFV/hq/fGuuzHU3zr0bp35RCS7eqwuUZtv3jeJNyKfLeb4NnlR
vGjWliOo73kbqstuup3cZIULeWUO7ilB0+f/IOQAikcx2w9xm4S9bhf+nqpW3HRnvV3OCm1Q09ki
LoncTJwqmJ3X6rS3v5QkIb7WWOChjxdft9heEDRFws7IJa9/aa5ZBl5jv7kCbUZvbjnPg1D/iJu4
1YO9lkskouTTxhmNscGQwiRe1BL4F4OPwE1gXmR2RwPewK5y7ZT5ryGzR38hamC9wAQZdqqspCP6
JyQ73vDQHRXJONezdGE/AqiTOcbxv0L60hYnWeo/LVPdDCbkztuD3A5zwIdjct7mCXqZN2CxgaoW
H7KF5BAjidzrOapyRpyyfnE0b36qJpf3ZSSN5XHKbgVk8Rz3cnE+lOr/iAtEXdLcvhL4iH2bH14M
txfW7wY/0H5HGFnGP3RfQFsPajl0mk+4A9ZBDLRvLhGoM3Edndwort1DezMPkh4hZmipc2Gesm20
pee+ijCHglSGZ715/ZhCd2l30o6hiLBNhR+dhxYFy/Y9m6ZjCcCGybY8Z/fttfLlZ++RRFmnRHlh
7UPGw1REcG0vuQ7t2wfe7OutQHq22+qZF8OcOUzlA7LbTGz+u4sD5kUpVgXhZjr44rbWTRX0AUJZ
ll7D7wmAFhIMYyjWznWNb0X6noc1jK81JmKL8nHYoj1vzSDu74geoHSKd9BOZ+6Ue4YZlvJBm6zS
ZbaGzcXvOmaCjwVmlK71XYOzTAcboeayH1vGygLMHSIA7D8IXHJZLc2e/PzX/zqXRPk4pW07nzE6
Utl4DB1+VTtHvOaQue/fkJlLYvtmyQApdSvDNLOZy6M9snPIPLU6ljzQW4zC4keQ36AU22v+vIPj
mZVZatlh2iQbzmzNSCpaXhTHvnWI+j8YPy1fA627NNZstLoq6nNAnvJBEYBDiGDZfLmzEj79R1J1
9OBnfiUkrcjSqirrUrZ+ShigPulgbdpCaXGALcUh7pZJrRtGCG2+Kwo9KzWGHJUI6psBcvvQfaBL
cZwAcjkQWNkLjBUoOXdCUsSPTUigOhm3vDPFbW8tt0F2x2+tS/k6gbvePyYsyodmLSXqKT8X7HlR
EgA5ya2YK5MWmKQSsMbkFuuezLJppak3NqvBc32btVqSqllBLHWU07CKamcPX8I8oOGuAJaBPDcz
Wkoxp+KYkzzJQ1nUkY8QJ/h+vK28vmu4g+p6pepy+Gx0yViLe0GFVhw+IiSYZGZgw7Fu5ZBN2d/1
o7504S9UHOaqXfXCPdNYlxP/ZUXz8WlMspRdlwizUFparrt0KFtuNA407WGChnGFXqc5HtnAtQsD
vX8J00b4J7Pn4NED+1utWbCoUcWMZC3KQkxSUr5ThW+JtLivwoWnRmD+zuTGIuBnjYrQX4KW9G9O
vDudflJXzQ3MtLNnUnYMWAayCUCkuZGi7RpOa8Njj/tn5/krNcQ6mdrfCszYyC4yPRf7fZPudO7b
z82OK1MzTMyaW8LSS35FM6Ym0/1KNOYRW6ZffaJ5QoWwm6LC79PsK7ukZjQA6IQLcgqFakwrnXb6
o4N5/EEVcQkBQ+be765+37cel0czKtBwMQu1tTIDbcQm7wMjaMUuNuJMQ9Qq29G2oJCAEA95Qx0q
6L1LPC2ElWOpUHRnoGVmdKc0kHIEQ2D3WPnAXZOZ1soKsgp24Hst4Vs57PcdHrcKbPArbFirKcQQ
kXbQ7ZF41CDmyUNDV22wgTm0l4JQSdP0eMeluwdRJAfMXQLZxdfEfZbZvrvbS1YblIfFFeSzzrA8
mvWSoLeN7K3SzBZAtbz222SEK3sZJDru9GF+b40ETTjRQlRAGp6tamVOiUu5qh75KDdIj/SeVFDn
Jujk5q4VB6yuiDnLgIIkiaw4sKw1OOF/PinXq1xq5895hd9XSnA/CKdWxiXjrkwf1pwrEFHbsNpB
iDkbkezyMqoLbkkd8/Ja1KrgDrVs70n0y+Fn4clZrI9fWUWU41+gcHOmmS6kSMLI42ig7gKdyM0V
dIIvnRut2o94fno/Fp8Dxp+nYc5HKo8T5U1W+V99AE/wErHTEG9W38lFO67GO6cmW9tN6BQ8JKQ8
H3u4uWY0jWLPgrn90gTcMB18ykaboee1+zCqIgUPAEa2PI5xv6nN7Tgo5EUg7hJKfxgA3/wDm4pO
sbC723MD5ZsuxneFOTZrqZnKswaN0oC8CHVtswDOWxFRl16t9/BME+AF6mem9AbRz7jrVLdNoLPZ
KLvhikzWWh7v6X2t7P1Wm7MIykCxGbYaS0XQdiVyggmWfLDVeJPsBp/xhvpc1pEVTa+WnaSNSliE
Q/F4vlMhTb6tYR8QSM9hUnxqcMoTsOLkmmfn61sg/bytjz1XLEzqGSWoqmDpfREKPoVyD7GTYiNU
9uI+9yFYc9RjrFuZsFw+0O9hd/FBPdyq4t7W8ldJB55hXmLBEnyR6hOklYH75t8AUKY43SSO/mL/
FbOJsxUhTFQkSB0v7Es9GGByKmlQSQRnzOeeoqsIK4THhAcF0k26SNdxvwu1xEXlW/MwOs5kOti5
/G50XzzNAirXFIVf1i6WV3Ex4ZVTOpB88bY5b6fW1hV2bT04wtspJ36s7rS1twwrGqs9w+ULDvPM
0MXV9QtavZs+FZpxbKuNIAp75S7/mQPoORbOw6PeFDK6myNKmlDlV6MZuciYwa+HQyxr1XYDs8cs
gDOrXKV8PQiF5CuavtJZBFzB+NX193bXNjHgkwk3sf1AiFpppAFSKJA6gZIk58nS6DGmNNlLvEdh
7IqT5dL3QM3RlOGjHK6Ku4OKi9G+zAJZ/y4wPkvVKwU0LQXhakZIu5WDqstJAv2KPXDyUQ/qbVx7
RpQ/THZhSRYsCCEeczqndw5GdCYZOW03DWq2GPH572JHjbTNHfQWIIVxEheJEOWuMBkeaR43CKOz
FQXu/Q5i8iULbeRXLjeIIindPcgfvPFflK6QPBK5KgBKqEeFpXgxIJR0jVDNVZbYteydoEUinm9P
S/eiX1nHS5m/qpncRf68uqUiiXommYY0Xiut8W439RUIuDgKDXPdm90/+vSWJZyG8CiXDA2QYROn
vWhApKTQbEOkZvijVp8JTQGDmtfN0hOpfDmX8o7NdkBZ9aj2vCPAqjD1nbOkj/LsDVNYbqUDH4Ey
/ujFbuCsR+nUTl1jJuVDosCL0QgEyvYNP/UD1K8KIxhbUekxj1qnYqUo3zlCBGq4tLxWGkU/pRvB
psq/7ebmNVLMGJw09epOlQxJuOmEiApoMrmdyPpIV+yIaXaCbBuIV6l1R0Oreo/RGRGvpQu2K6ER
+3W7+HXCPJMkjAYagfAyIYjG6p43l0ZKgG5Rwolym6WE/XjLmKcpeDUzlxXKYB+oaNvCma40epP2
Rcnsos4Q+k84Bq5MMvZEqc90fcJjwKaie7yY8iPN4mR/a6vJvlcPzpjg18RHMOgHo7sPX5jClJem
WWrQNGj+W1mZHbGmVaDuAKJHUobmiKX66IQTk0jUKKPosiSZjzwW5H+Xo4wrp7iWokIA6GWHkHa4
85FJyJ0zGnUGvEuruWj9DQSsRs7FYeWcfTUm1BgB8ovONbXS8BYk/ZMS06CmLp1xBFZGz28sF0z3
/F1v5V/eN9ZVcQ1b8iKX6QaxufrDju8OozBxC0qD0gA/aSR+JpQrb/vp+ys3yb7grbFr5VXHGjaq
Bo6kw44X2DVbv5e16owNDEqXsMR5Q9kzAby8TgNm9PjvddqAWfTjTkZ5CIIXLzQxjEPGYQ+x3LKA
yxTHU+Qv1AfzjYJuCIg9Ddz0vdH7AeQ8VnRW+h84a6OYjGtNrMZ4ZvKFJxDJMmtle32Y910PN69J
wZ7TeEkYukAa7heDvgaqaxC1ox0eJym6B0vnXQuZ2gQZ/jaZHihTOHNW7oTIbhVb9TmTuBsBGwKT
LRYjZwSV3g8HE33N7GVrtOrDBchh6QZYtUspcqapmNIUYXx74SMbMh4WcOruPZ8idilNZ9CxU8/N
1qW0bWuL+HoQVGjiGnjpKapYV3sJ5klDQkR+Ack4KuhYDaGS91af5pkzlbN7Q09vb9MT5AUjI/tB
lS7EUYr/o/zociynnLpcaOr+WrMuTUEPYaqgTLhOfDslRvWeyHbqdeWP/tdBU6IEvXYhKjCkCErR
yepUz8OowmFXeFF7r033boZyU/Ga4loOBlA5Nq6solPoB9n6J5tbewmY+WjWlWhG8x4FmMlEfKCy
0+LHO4taDhLawuasukWlKJqLTJGQnDsG+kN/d4DQwGz+ys00jhfTb1cKShbFsKNY5yDTw8fbHPzr
C6B1dIgMvtYJ7/defgTxeC6GW7WQ0r+2UVd+4tO0YDpAFd824f2O/GP+hiUU2F6iWdNtXJy0Cb8Z
S7v0mz2jcWtlTfVR2SvOMbTYKUvK0d+UY1rNOwl9pJXxcAmKXsmVNmTR38bNh/d7T0VrOEMNqmQK
pbJfxQMi4LN/FsYc1wjT15wi7C9SgutpHC+DhH+eMZwNuFHiOyJMYRoERcB8v394q0m7AtUj7JXe
f4yuA5/MTq+ycdgeVYZGpGQtp2Jaf58z7FNtGjNDPhMNbtwcyQMGm9hgj1W9Kbc9fkw2ms2ZZa79
1Vw4+ZpYXwU6EVq6UAFcJVZoFS3uKG61bDqX44ro18QC6VrzxUjOEIQThtCWOwRGhgAsxEbls259
C7aSObORWveNTdlvsy104mOTsjPzc2tTZPc16XnAQUmLxduC96/QZ8OIAzYCJzYHfYrQXshkQyc0
uCUx0q8iYzGknnCmzos9kOTxbDbdGSDI9WgxWlmXaZ0zMHk6rEVDFT6Q9O7jdrCSEX+O1LU3iFTI
2mVsh75a2dZ5HeAdSNUpunjcS/pvbur3cZHedmm3Qboy7hmfWTZUTs+oWMcIHz8QQhfusnN8aaWK
d4a9ZDunYZwdIiBwr6e7qXDESKLF9nEYsRaBqrJH++5EfksfCrCHCr0i2l05E9kjSwRnW8GDP8+i
8jcB7zHF8WzaqD2bWU79V9N4ZrbDiRrh9qhjsHJ00638dTimVuk5kV2Mobt39npKyh0NRtkbBsVs
x2YNEfL2PAm6CUN23XPjF99x/TP++vRGwn+9IJMoTgeSSdFdw4h0Xh7vPBQVc7kWvuQ7R5W8TOyq
/zsW9W670NQXhOfctdN2a9dfzNXRal5zbGvXD7S0gvGJBC3WKN7yQBRCpJ6WlTo9fXJCw9uUUb9G
uX/Mgkcz+SdtlqNXFmqO0UIrdOFzPn464fNGfcAoQvkAj6TyBogmVdEWBVAes3SpkDxPG5TWqWaa
pOCydt9NdOtkwPq3PMQ6fT0J91G2TzGPiDTWKihrwea6tdSydX+pXN8irVAwQJlt0+sQ8I1e40io
8XRSqViqKgmCjukXZziHD3rqMsIVECIzIxuxKAzc7ii5/W+fyCawI+6QL+cJ6UU7newJp3svfdjX
LvUYchHPHp6IFJbVK7wyNv3VNdFtCz+nDW0y+NczIOgQp3xVRC2hOY/8Rcc9JuheKyX7gLE41LpR
P6Hf1Os3ixMFglhN1O5W9yVDFI5IdRFHWdrvHMheMuVwmWZfaRGZ4ie4twJpELW4RvcBFQrwCsdQ
5X8ymsacM+7CvYdbab26WJe0jMIP0bw4Vyh9d+/e7ypDFxFpvhxu25o28ULBU5djybnJT3d/mVWI
O7m1PIu7t0MLcUtQnGi88sEuLyArMpA9d/ITN2RiZhgVwdQ8xDj2vqezvDnrozOLPZMvfTWysIt7
9DgTF9qWM3QR8db4QK10mQLEEOXLjunagFJEZWMTJgT8UzTUGaG067pkQ46C9ZlpPKPCmLnxBuFQ
3ZUuXO/wmeOG2H+bUIsEsikgIF4fmy6sFJWFEeuZ8DQyV8a79triLZkVYF3M64XOtrIkhA31h+fl
YnCd7+9auRLaxU+gO7MD5p/FhbXmbYtkMxcN3V7kPTtTp0F5dr7JKKKZ24NLVOejTx1yvL9TLc/b
u0cJNzm+4P4CehR8BdMKVEE6fDeOwbul//oUer4GM4Ij/oZkJ3fUTKbASWggfA/n92Ri9kFiPnUZ
T4b6l6k/zUXN/lNvLouTPeg3TvAkyuXE+YT13eqArCw0/VzZpAVRf3Ax63/Fug1XhUYv9JrKkiNa
ICPo5bHJw4E7o1YHc6Yb7HJ/G5lvyb9r44tMp/zPUZ0i7KfXNSFV4AsIJP6s6W3DOe9n/N/dXgQY
4niPF9cpWwDMeKarYPio2q31VYwkON2u6onXu+dDCXJpfr84IneCSc/xBqUFh2UlXELLYk7jJ1+b
pLzOGOWP22RhKLYjkLdv3l5vxAbsJuNzpgMvEFOc7VAkCQNBMbiBFkwlh/JcePNFA8JQCWA8Fh9u
i/7VVYIQy7yu+9h3O7BNjdG+xrD8KZlANSXL21JCnIZw8O1FsMHB5TsugyuXsXiV91GPG9XzTdi+
DViXYwBDFLHwBEqko3QjG38GEh5w9HX/uR12P+Vcfq171ERYi9XBGTejPoy088kIj5IclIA+dxwy
nVK5wBxo4gFWQsc4lMW4nz55HIEFrycycCuPaPH51L89bkfadAkaiYmxjtba2IS/GGntDsSW/Xp7
vcp8BUNb+t7KmvB4EpyvKgLFtOFhWE+uEnVpJktyl/UKqYR0MgOHAYNhpHvyC3U1M4DY9U4sNOhz
RZF3OTwjnHvMk/l9L3m8dlvwEDO1Ja60/fYHybtvovlKZUMUY7dQzyF3tnFmCpoVF9scQK3dfb5z
5e0qiQH0mDX20TtBjGj9jZ6krNxbJ7yS2JjTQnSBgPKeUak/s2rpYDrMFIOsy5d9rDhx4YfIKu7e
BtUzKnUM9vy4Dw5tvWgvx/ldlGNceDYeYHn1SZnZubCii4g0aakls9jvcNLx0cbnl8nyGm5iwbRu
xI5OmDw8AOsMkTe6DEQJQGeq2i2kC684vzFBKwalwVZ3T14ZnrH04gZy1H5yk79iqeYT0i8qg0ps
utvccuqK+Z0igm8O1u+vCii0/UAwC4ZAjGkURq0a3cRmdS22QgkqLn3s/bSsWtbJR+4fQVszRWgw
sT8eAQjjiPsWb9JGHzInW1BVETvFD3IOjxzt87d3IqWwdhxWqEDA22GF/G8tYrQguAO92UKL7G+5
DLAf0SkPojTQ3Pq4JHF1ciMkG13VlM4NH6Qg40lKCf4ZYEF2xVHqhsdWYAb8Y8BI8M2RpVpy8ZEI
UdTgKwAJ7fnMPHIZ99etWHPu9sjnvl3eUSH1ez6tsiiMWXu5jPDYOAcRAMPbZ27X9QMjF8LAnJdY
UGSQWDihZ3k3KQ3gwYU9bk3I5eJgkIk0ZNPE1bHrtUS2GKSGwlhXyS/shLLxCishz8F8UNQEthln
fJUJqT3nRSM1CcqakkxURhVwmwqe3Nv/uwnwwx/xFVv2YMkTz3mT5lEUVB4rK44A7OLKCwCO/Fa/
DKR82HD1+jClImafWOLyh3r50lr8WFQu2clrYNWhycdbBVrYU+htmLZbCQo4SJxPSp3GbceFQIQp
NDvSBhRM/ZILteOQCKgIxOVwRwS9kbwi2ggdl9tx1vjm2MJSKs83q1Z6NTfy+Wj4ckclLEjPoKIM
UVr3VvE+q0i1IDYnnjC/RxX4e4cqiET/w6bpj0ZR+n2h0DrwwQqfuj2nti+W942lVo+CeHfJwm8q
xj02kW1juVi0bL2rCv9DG7uzGZsTwGpDGlGQhQQYZKOp70F4ACs0DwKzQzD+Fm3WfZO4cBwc6zje
yfpYmqLAmoYsaygPxtmo1RMDuCtBCH3z8KEGf+TVxz/3BkkUl6HCSKntTSeMJbukplJCrX0kCn3K
D02gQL8MaOqxm/CIyYMv1FXictIxSY3dY4FmcDPoKEyVuZHAPF4nuAhDHEx2hmlsfkr6xCnkRQT7
YHn9e/VrWEOt47bXczFZsJ9IgEkrrUsXJhFfg8Th+VIcYLP0sSDogTr6oPjCNbj4CNjnAdDCfEP1
ZPuXzgJFU4PNphkZ615YMGHH3JXfPh5sZtya6T5LFQHEfSp/nz3A0WR6FOt4RnGsFchaCScaKVaL
8p8z/iG1K/ShefFISRfup3PIsgia9v9UrMI9/CpoDUv4HeEn9/xX1KyC/ryAx9PVoSTGbVSm3UFL
lSCCXCKbSkrjmC06r/fKY1PetPZact2aZjMkueDT2Xx6QcvqNoS2TlKoMGiKy0s83QuTe+z5MIIl
oeFBkTtTpj1I6XPC9whWYYD31ujBEasAMo4sgLQN39Okj6/Ra+3Zcp5fj+pP63+6VoEQeDb+3lKS
A1U142Ma/oGV36lvKHp/y2ZNQJ1i5cwfTqHq+GzbLJWySBDVYeZmJnYKzdfQdps2njNZW3Ixqmg0
34ioz+Xw16EtPx+RtNq4lu1rJWq8fAzRTlgCtU6IiP68vfH9QXQpUzYa5MHmSS4rgNnws17lyhOb
Vkndj72WTGuZHOx5Cqd7bNLiEDs9BP3i0zpQvGOg8mCI4yeuLgB+0R32LUu2qG8fptGq89KC+84L
ihqKnNGHf1zwHaWvEF9yfOwK9wJInuLYIOSCv+Jo5lxiuArD+OPZtw6RB5DhKVX+WmV3tAEZAvR3
O0Kz+hOseUxmHDXGJYZ4hXH3MiIDBgKNcSCQ+bvuCu6JPXcfYelNEyio41LnUYEdquOzScZwa6jG
1mR+b3NzTtJ62lg44n1NSDDCkwJXwM3clS3dK3kt8roYmxtJFkwtRBprxXGwsjsQn/UEwCKDGnm4
1SwvW1Ztx3wzabunygop/hzSL+VfuQBaJgW8CSgagoiSSBVfR2kiluDdcWG6Jf/PhIukozcSbDmb
RbvS/PLQS/TLHAK29NwtQeQjAWkr+pfYyElsj1IB+7Zw+xJLmo2c0FCjeIaIJfqSD5gmk3jL72qf
M2K1LdsZ2N7Jqn1SaU8uPDa344mgRQn3FrZVHYgY4IVQ4DzEtw9om029hxi/ur91ZtH8yHMC3hs9
CmVosPP7PfKDA1twNEQBEJJ/BaaHc1S0v5ZzfXvCKAimQ5OMnGj7g47+iB9ris3HkA00UFIjELuX
3haN6h7n64gT/CYJE/8Yax2bwPwRbJ1wvC9X1By+PM0tqfb9Yo4+qwK+hhzfjgZ9ig1eRYKgClTc
m2U6gog42sD5snxzlYbi1wBDqBaw3IWD5h5Ggk/JdVzB4VIqy8h6v8OH0uFBvAveZgfLPPdEmxgU
5Nf0aFUTRN95bzP08XQEc6AoLMM9js5Orv9ZxifYi4SbvUzodnONVu9WU2ureUwMQrYuRrfNLXfL
s2AkAhwEjJKL5Zn5yTAC6LBNQ9ldTh+xnS0Cov+5w8la+hqfFJsRH2d6lGtPRNC/yawRN8p/qV9I
2K9KuP8LXgwZXxo/AFxOuTGIfaKChzzj6ZWWNUxnoml/UtObY3ZCCN7RQG3Hz/3jFLkuf+SvzziK
9K94Wwn352pKLrpZulOVoVHgm5tXVcc4DevZZK39gKWbDwE6SDlwGkGZLPTtcZqYJ5Z1VnyNc36R
0OJgNEvz2bBxmsAUmSYa3ltA0wsIOaAanOv7iNmTAtRhp7Ww6Wx5Wl4OoJIlUjO9KqrjdmHLRdRH
axCjaiPwhanrwBptmop5nuNp+G3YZNoYfKpnItAZTR4vYMl8ddAKN8WhyGiSOHWMAGLumL9LdN0q
zQDTmqhHLhegQUgyl97I55srAEspBmitln0rUKzUV288lUED2tp6GjYlybu4iIbvs9PvVoJQtLrY
J+RBSgdGftVHj6+2py+Q7rHZ6sjNS2w673SqLaPXx0JcY9nH3WQSz0ZsTCQKD0uUhPe+cAbVLpRS
imp081VD5GFOdcdv6679kn2YJnqNF5hKdNGyfzfENbcRpYUnLU7dLc1yG0wuyb+NQ5xvYkrMV3Hz
cDGgD9mmP2zVb/t+pI2XN11bPm79BY94jm8aWOymmRdQrZS7iGdvRsgTrV1kZKTDF8TR7tf/KC69
WEE8JstXz3jNX7h9y/+jsRk3qs6tC+cwZUy0QGXc1DC6QTB8PItGWYcXEC5ZXMYZY0bAyWGm4ufF
1EQ6PBLPTiVPkOjwcMtk+sPayhcPVfx/+mGdA7pjf9iiJnRSvm2/O8gA4zT2+KzhIr3cTsCu2J/z
A5KtU5wAck7mo9SVvztFEjBQuS83EK4LzlG4KMWOAvnBHmBIGwzEumtOh/TXVnqkQSH3z5IOrc68
xsCVgvBlvJyyDfph0JRB9q4vqeCIP2FP/LMEMQLrvivy+mvcfSfV6KmOXqXrQcn91/kxSnSKKYRo
oN7APdReQo69dDbY+XccPjhuWVJz77vAeK0y0VXYqabeYJYMzb19cYwu/FUwZppVsyXmLLn53/u/
nvyw70A2O3PKr+FNyg2VcKvINAY+lYDt/Hqb/FkkTz8PQTGwnS4X8qY5jU9WXT5jaZXcCM5AE75k
RXOO51PjhUApye7YQHltNmccah618FR05bS59FE8+nT5wlFIBcsncUyZVrehzcSka+4HTpOngOEf
JgxVDH3RwpXABGU8doTUq70BNk3+okjtypQmb1aSNY7gHX8PeUkeehSczmegTVqGj67NJ6kEIT21
aYI2cxps5xXJxEwCvlJSV7t6h9HWtLMp5KZ7TTeltjGJB68SbdsKZg5JWKpjaLLmwzV1pC/GMXcz
C9xHmJ6d6PJZbvMYdD/ZlBCChLFFgeAnXrEy11WOdLo4SW/HIDDZ0EY0an5BICG2gcv4NzTZWyIV
3va9JMNnhBFOfX3MWvZhhX0SEApipKFJcCFblfPqlQII7jdcAr0dDzFd+nTTcB5TDyuugHdIEkdv
Z+XYEaC0906lPW9v3fhKnjAeJCx/3SPytFsLAsMomT2Rqs2n/1tEAOOKc0lJAtkDOoLo2yAfX0h4
SMbVwJfUUuEvSKiXTkDK7vpL1OqerZSvxE4/En6XbNNOkxyFNjZSsZajkjwVqYtzbIHx23XDYEz8
AHzSQjwHJLnyM5WPPpqjZPKvzMAiVAM58i/PqDb3qym1cX2YM7+a6wHSjp76Dx35z8z8OABAfR7p
lmg+rrJPpNLFHD3DaXgf9sBkps+LwQkt349PlYfiTcXPd3YOzvm/hdvuz4ZCi2yBUckEBrX7x6s2
OfALXJr7DazMuaeLAytjd+4wZja6CCfybjMNkR8pbOodlt/HW/Skt0E9IlPSGctpMdB20ZL9de7C
rcCTAC687gMUW5JEepmw/mKOolnBOP+xP3QEmrpdR4aTFC2AdSZSWBgXBlWAaLDw6NrmukIQeM1I
KAC/ll8giXS+6QunsATa+/gHCBcnEjWzQigkzP2m5730+uoSDKoMq6VtNrDa22tL+G3zYJWqhVEE
bo5Uta/OHFvkGx0IDtTozLjUWTXBoimslqYjvx8LlyryResDD41t8MBiaXTuXbGTCwLnO84yeNKC
gbHX8w1SQZWGDTsANjXqR/zqJoR7FDLzWBw9gBkZjmyyBTjd8yGpajTedJhZRuP1utXo7AZt+rgG
eQPL+NQ45Wj1AiIMyMI68yqQxbvIztUtCUfEUPDPHwpCHism1MdqkeADmHNBmXKpu8ByTVAz0TgA
CyRzT8h5uAeM67mvmE6L6a2HAYJWZaF+H4DyD5FJOGwfDELqGmE2A6t+3YtnYZXmT8L6A3MY73Dz
IiBkfVMl22br6wE6Wpx9AavCsFzna1QNNUwEMTy9xbGu+KTG2+0maq7WzAQtJ58h8ca6j0B7QLry
kOw8wphH3Y6Tw1Ld/IK1WA2exys3rR5CAs13V4S9mJ0hzs82QAg/cdImyloqtFY+HdKi6TaAnI0o
kelHx6S22oy55RrIpQARLpIdcGnHkwxTaHck/LeeWSVv7H3ckAEE9B3pYRLNHomuwV4pwRYlozBO
nUyvOCQZewBTJrNT4VVgwjxOho+yveBUtcXz4497hK7g2AfI9FC8Qly94+gG5bKRK6bjigcF2eUU
ijfeQ3hF5OjKdMPT9f2EpzxlYinrjcE77UVMFYh2vGOT9FgWqFr0oDbGEda9dgVhq186vIWEnbCf
HL7XoNGNPnSCMe/BpIN5AUXOHORIlPeMdAFZY7NzX/BbxQTdUnqdLMlZlILi4DUeQ2mjXron+FF1
KIw/6zWWiiFfrZxfvcE9wnGbUeW0J7p/qz5oHfyMQSlZIesGb6UHLkz9OCYj7J2VF3myCF49kTwp
BrXXzqLZRdTzp2wZ726Tr4n2pD8oFk83SXZPGTjStKZRTWftGkLyi75h/SIcVSNnIiikvHdcChew
v9+sCPyUs9OzH+nkcmOwtdmZBCx3R3vkIxumOhGm7amQxelYI7tjbrBJra5N7NsqVUIwabo3bP8K
kiBxxWDk7CLTxzpLT43nRZCh0gSTrZhTPJSOWjlKgGTbolTsIa4pjLDYG6JXHvGJAT3mFriBbiIA
ixJsG/hF001lfql/lZcUgMMfeaMJuuqADbvSr33RSXd51tiZnPJh4cwD7OFpsE26HA8t4N6vDEZr
SeiAUybTgqcjvvRu4Nyy3Lzbzw7JgKVxxHzhl+UjJkpQWNx6mjucGjsVZ0keZZQo45Z1pK/vbQ1P
PM1Mxl9AylgLnI88aJlTCYmkVJkSPsDZr8hrVk7gQMH2djIr/zTdop9y+pvwfJnyxHPvjh+Tnaee
BqS/Xiwr6CGjxUKG/P5hHRGSV+o70r18LdWViEEWk+FGykN7I+QHVAt+ofEn4yW127yrypE2ajPl
pVTrCVEISyoHaInUJmkOBSwoTtaYaLUev2nbMWKqqOzMxRxg6IOI7FOtnkkhHU+UmP/D7QEgm6Z6
tP1dOf9q6/s/w/lW798zP8hN0TCjBX+B2Brm+OJBjfpDwg8q4FAhZ88ko1ui2CMlq6NzbSGGneu1
lxA3gU+qUipwz9rVl9nsj/tD7DiDerbPJLD5UDesPYXFkFrj6w72QkB8Kv7TqHD/D5fXR7qfC3l9
vU+dPpEGw2XxxKdO4Z1MXW9vE66yxfsgahSwxLYyfh3GBpk4MN2ddOlEo5Cy27hwBT9fqxH3gtMF
eo0IFYBiNoDv58XBC/v4X/yBmbUck1Xj4GzLJXDxqmpcRZSC+FtOT3U9sZEPHX2n3nwAMmv4gbeH
TrsfIyq9Hi9+IUNq7lWGt/FAVGXBYXZJWxDypZ7F560G7+yKcmfGtEcY/62o2T9HBbid+1o46l7F
shIzEKCz5pcEdUVMjhBOtaBoJQKpqq07lhuWwMFlXCHZ1YuDofpWY8flcjUiBnTk1vJtgM4UoDCf
3abNNhRbKwXXPNIq0IJnf9YE9zTqEfMchVXE9p8rqZEmtQNOUMDYe0lwlO2wr/+gO+y4lWkfl5Wy
qlwPmwFDbBBSIefhx4HNLZxwysv1SKBYER6TXbPiCuTQrr02m1Jsrl7yQBPURlVWGSBeaQUSSdac
mL7qwzl2eTkDYBhqRayDFF9XnpG6GCNA5FplNbaG5Z4j0UCs5Pg4S2DPUPuVAepieqrBgsZ+rh0W
v9ZtaIjHEoQvEyiqXCnXZcpugaaf69nD0dMnL/H6lg7FUo84UXX142InBSphEcnAlR3wD1EBlZy5
sLtq00ttItzk3A96A5kKkNpdLoUUmlqAczIVZ6gll1BJB9+JLZByr575roaf0gwC8m+aFHe1zdTX
hZ6EfdazhtIev0HB3eissvgoINAKuLvEMbXeKwgjP+BUo7wazr9kIRnnlLptBMPgpyVunjncERsa
yBUS3P5VFdY9+H3ChYzYRpB+y+srfzWErXy0EpxMXNO6Jf0qLO5e0hf8YnJV2EhUxuf+ESIpzNzZ
XiXm0fbaHfYetiWNYsx2Xhmm8of4WTqJKm26Ir/GWeizVZK/rkcNTPpOvbDZ1tmOMjPdsvHVvzjp
gLniGAkeK4xXCtDDIxg6dJH2MltBM7egRVUCex15EGEcW3O4+ER1FxKQv5XmKzAsCyKccPbsE1y5
BgXRxajHK/ARSYdgJUB/3+Wv25n6fP+6RfhbA2xo9PMtLQokhkIm93CWOMfCO7rfngMIPKuitCGD
dL/3cm6p4TZuUS9f9Us0z3u9KrfQsNADUTAaQBSQRY4MUKtmuNDXOqRXzWuQ7pCSBkKLYWsienYe
WHnnTDor5Y231386Ax2RLQO4JulllK2qVnP6q01QT91VLA+1bzQZW4DxSdiZDpNSxrBOj1erDuJk
LWIODOUobvfn4iqZF1OTwlLJ7JgWaa5uA9Agg4GAfYgY2eIwglfkb4CXWgBom600zMmVbGazwA9m
9t0ENQ/nKl8BGsmZvLSpS1/fsVyP7Mg98yji3bMjqYUVvBrvJXsg3GyzrYB6Fy1CBmyXzvQB5kOY
SoMpYm3y8YKM1vcOoODbGcDAzn0uHwrev+8Vy3DA64BelbOgwndNGmNFF0aWpju9+mZl4UCCJB3y
7V8c3YDhDaS1+UMR2n/aYlHvHcReLZZV5zB6g45OLh2e6YME37GZzyBovQIo47IRKeJYa+sFrAfX
Wnx7GfUWV6uzhbau/KYY3aowkipIiE/UqLnguo36JdhDtqDjrjmZt2Sp9i5nDzYq72Z9D4LUoT/X
YR6+WpvmbK5PuddWeijyrmsrGSYQUdxKGdqDHk9b3VsRnPl8H7ZhYjrA/eXOvKZV5Uftv5Sf1Xpc
L65YdX3yUStBZMQFZdgXt8CZ8TDT4D2xKcmoCqWoA7QSNrV96n8/bCT+Ilx0ZpA3t3FmbD12P79t
NHm7Cs+CfmvDpvQgazvDirWwVn6ge5SatLabHaKstJUW26NP+1+OYW0tsDp/pL7xDlRSZ5S2wDgh
vQe9cTCVn9XAoGIkGUX/n4I9nMGH22EJV1otpvI/cFdaXg1D1dJYEajEBWjXhaY679W8PVMBgayw
eMRVSH+E+1rd1AOtfzt/gtzCU4hHiZzQfFejd+OvL7BoQ78vikNDzApVNbG67ywwnfv6Y1xrObA6
yogXIORaXp8/lYBKanHEuxadcx0PF6FrxTQ68Aq3q4kz/WX1GolfRyeAfPOyAD3SZ4ttrxt2l9d3
OHZoTvZsx0dg+MzhcQXKeeI/JL907hHRPrajM4Kmd/uJhVWfO71p/VZ8cNCOk3Hz1XdcM4FyJ+P9
LbiqliRYoqPwrHfA0BGC8P+yqvge9DD/drdEBSSKLtaHv/9YMO/UUd6IWPIymgW5CQckuJPFi9tV
8iAFLx6NqdvIwxrp4DZnwiOjFcmtMYjq9mPK+ZnxnF+dPjhqrSeQ66BxixHAUqWu+9fie2+MRCOj
1SrbemDcmXgO8VTdO7IARzC0YuRBOuXod/SvqPW00WaMhPBg5td9IGCMQ0GeG8k/w+oCdIb2rkBA
4EOcj03K7/eo1GbKfimSUhSMHcQQ9IQlcB6/JKTyM4hlFF1n4ZEA8W13GoNeZQ1QQ4M6DEzKux9i
nl6gx/YKuKOWnqZUeL1WpaMUeJs0+tlG6qeH370K2FbM2T92daQoPtv1zBMtajb5TRb1fVyyjqPD
zWopd2LTm1+rch+gwFrePRtqsaDYPmvpaWKdLXwmfKnAECdNShhsD/gN6FuQlhx+J2Qgw7LG5Fw8
rw1besrKIxG1dPDru+H/+WmMbuLl7D3nFYtn2jEjKMhtVcfNyS4qzZhecDvZ2okV/KjcLWs1l3tR
G5uuyzhLFGH7KhGWMhU/XHExc+9WdrC8wQphqneTnjsmt58b94cFGGcd+0YWWBjCsFScXQ+5HeCS
HCK78v+dtO7vvczoGw1GppjQHE42UlxnVkmtAzXVy9fXlA8KOq+1Y5ZR7eC5spark3cIUfD6fLxm
dvH5dHcGDE2n+15oImbRVLkLmVHMjkvmmpeapXj8owpugEzn7NiqB0ovL7k0N4Yn8oBAhL/pmA8m
tq7su3OIKKNiSak568X96UnH4u4dsArEfDESXkSoYv/zFn4TOenvsJABiauEUBddglF6rfp3ppyd
A81MbTfU5c5A3hIsDb75f4BXlE/abNw2q2N1/YM17qA9SC+5JVh2gm2enum8aQg2PSCTFPgVwBtl
dlioYVTP/kn1an09uwjFexmnYNiqlJwnuEG1UDKhMNO95UdzbdmUuED1/2ZR1lbfSiwkOTAJyeds
yjanMetPwVdFzxrHon10GJied3qKdIpOpLijkN8dCa3g+vuFo5WhDgD7g0yGCLco5lOoM0qNhWEZ
g0ZeHNoa3Lodao51L6SdE2nfVyAkWVaHU1qsev0zrXBnXfoa4KMPDvwkUnc1kCpJg5BsDLBBDOvS
4tscd9K5tm6BYK2HpQaqE9lm/TBx396QehCSj6vaajVG3w2bFVsxZ1uppk803PdsdgZ1GFYITqTg
Y1P2p9BudnMj0UwcBDYvtgQ897/NwKu1yt6U8RyGINoNRAfbPz88qKuLCQLX2pHiow4noq/3YTeJ
CfYM9QJki2v0C7y2zU988X3K2qkHmC1CRLkIFnfFPjiH1tNLmJSjgNUxxvbHVHmNtLUZQBmFBcQ0
D0+8jx/6CB1m3OJqYHHNjRsSEPXathNpNOxs+vn+I9mmSzmTqp6LHnhA286K4PyZClscQNXmMO/u
3sSt+9a0fxr87HSZ/f+MTMaA3ETbh1ojSKh1LzrYU4pURszuOOcb58+wpO1Xtobn+GunoemAGpaZ
15/t3iazqwJOG4DrE405lChI573MP+6Cxn/w0rVQNdUGKuCrWlTNZDezks16w2yPH3IEtV0oqVxe
Y4kCEZOTNc2KIhZVerOT9XE3yssV1Yuf5ZggPWb4f/tM+tl+hzkczNKvziPaUKA2jAM0jYXEcRvK
dCXX2IGvS5wbYNkYI4WhYE+ezaoJ5Bm5Z9VwoJw0l+NWlgoOT2WpCIY8eIpHe3+LxbZL8BnNVwFg
+V2RSEOXyqlQONJaULYZKweLx4DSAzOmiKWhXgW+youF14Il5baq+nePSZdYIFDN5w0mV3mQSUgN
IzuqE287ygeXKgBBG9Ud04UpezQuWfh1FMUjCM1xMFJyeDBfFTwRRu+/NN0GFNrjR2ykix0zgEJ0
BK8vV066ODyk+0Zr6VVFssvnFXSHuDj1PlF5DNf9Pvh6k3f/UZilX4NaSEQu9sfsvYDBIWRLhOvD
cQOTfQSsuJ2JQGaWiTzb3NHLz3x6unUYtZX61G8mDdsjH3CGQzxSu/2nD++Pih/9uabYscZZaKE8
E60Xbn238z934QJiO6rVQglVwsMfRYZ0suuxlus90UyIEYodS3Vw7y8CgBJvigha54tifhCTzu6B
iTBK1Uc4F8IK59kBC1CeBoTgIjnOO2mBQ5fWPtxyE30Yy+z4uVGqe5aSGR1BODPfIqw1fZtMl8lJ
TIdp8JyRIUMZsTzs3tvxpXoZRnMQioHbSusBW5T/2wPDvXvnlppkLB1BQ/CThajk4QOL4S5TpR74
h8Uyjj8BdUqt2mRHIVdoY6brXxlhedYp1sWElyZIAK3USTibJHQE+eTlOqPl8LzWD6Nw/iWHuLC/
DeSo+L/MSjeTYxvsP+iSJV5GR6R4c2JCe4sOAohkfxpY6vbp0PdRYPKzkAzprlF1SB69OcPe8UiF
VSI9Fp71pdIPsfaWaBkP0JyEIB9vX8E32AnXaG3pcXnkuP7kquym26/lMbt/HHIPcch6xLX7JpH1
hPPENqGWO04LCh3i2r/11UoXYtgR+/N5jRPeW4NA1eRE54PnnF6H+zn0RsMrTnPi9Ugr31/4uHsH
PE4DPjSVQR55Lb0sREcUU/+eu29HdVrHbEAA8DHyL4RlkKnzZgeJTSCjIKrz+CpaAjiH4f1rdTxr
3huFxaaFE5VOUMundw7Kr1zaNn2HVxKjuTK6ibNo8w26TQqb5kri27SQrW1AnUtaYDNHmceIBCIK
LV51R8KcMBxGELnnQOrUYfl9FHiWUiRZiq+IeO8VJLKn4Th838Fz0ymJrleiL0F94ZqUl9DPxpGU
v61qHEK/MjeUvHbIWXEPj/VDL6ZxbG7+JXheSwwL/AJOHK8GJMgkiwwq2OvDcs08p7Aq+yo4HmQx
Qj5s/rJyayYaG0M8E7gZlN/jUwMZz0K0J9F5iPo6+OKTIxRlJaKW/PdNYnzwyOYsxe9Jg0q+19xn
hUuzYPbmNE9Jf6zDLq0H5NA7dT9/LOj77L7OrshGBSghfc0TKH9IQlcBKhlcmZYFarkzY+cl8vbf
pzvM5jr5YpD1ftOBb+AybAxKvdB3LCygC92QgnSB6zRdvDkhVHJ1g/KRV2uZP8dkAxNhuRR/T7vx
0GbKN5NK2nuRZt8Ksk9wbU9RJmgDBi+dF40BlhjJ4Q/eHUhH0yx7VRCyJCIxxvDZRvA3k0xUNBh7
Mskkl0nExysEE6IYZ9OpSGMtU7mbpjsK02sYxnI6ARDLMLM+oSHXa4FXi/7x75MMSXORoBFFDjFf
/es61SyTuZFftP+jtHrQNKeSd/ibrB0qOM4a+8YZTp5OWbYTX7T2T+/LyepDtOFJnZjDFj8Mb++M
PKxI3OLTL77OgnELMDQs+osNAIfSyIavvTyljZ3Gb2I4Dp60CWZFVUF4Ryxp8WHO8Czh5BsEn1jO
zvKt61M/Vp/jT7K3Rf2zYTdeUWElBODXuvTDW01N69pSu0ary3Vo4FbHFHujuahZfvwU680efTsK
R+wzdJYktpobmz92UmeC8jVVweOp7kEb6Y26Qr7PnAdxqWeI+EiwuzLDD0gnl6LSu2mxNBc+nTdd
C1V16Zw+TVYk+F22yOe1Jj+kMGPriwUZR8e6dObRSmwh3rIylbfRCxmuM86OtELsoxY6SE8PRDcK
oG+Ov1ItTb12NOmHUNEKz/q7lwaRIzFPbyGZ8AQFe5HBmYnoapWj2Po/Mzs4VgJWSwjsMfQNK7WF
lK9IAPGIvhFjTqVGdvEmLj1ImQlZRmWKb6Dqn3zRbNMUZPAdwVwWMiLK28p9zpAZ8slTbKxr97v6
ywyd5hEW7DV9nzwegxL4fETBLqalQlCek24DvvjLLnysOBcREh2CHD/wm0NEbyQxIIwvvVEwYjZB
N1ir0W65DS+2sLoAg4VOg8/mOROuQlDt6bgK9ggJPyqVedOkPptOKBVxXt8g5RYtm66cu21t2qGk
eBZTS9yp1j1qDJ+4Djn/IbKN88SUlUl7K5LD9KD9O0OdNo0agDOrXuqu/YKF0u1Rj5G/KvR5yXi3
VM60Ft3EW90abdupshQwLId7B2DqBflzsNT+I6wAl33FYJT29nC+VNaUI7MtnLcOPmYKkCl/xMzz
PlqxO7dD2o9ErJy3eV0kW6I1Lehc6vsSYR+emTT6zdfHHOKv8noV1KXKgXMU/eq5kncCXMH6LG8T
5GepIXmhI3BQPZ2rE+n8Wguz6QHAbWEptCMgBctBdw/ZGM/ckkwNJflL3xAjFWwlsGK/7auJHFpO
vuo0tbaUhBOIpZt8dF173O/9t9CvtggzZN4+flLT9ydJMwZOvf+nfA4bQaMDTRV33IuFJngbuabW
9BkfQ94XaEsK3M+PTDji7Xu1f0SgVKomT8sPtHlw9gYc2/lSX8w6AdO85iEUTg+OWFfr0/OlJcK/
vrYdEOltPzMK5i2hJB/lnwpbw/J1hbXOaLHS9M8lDCE8bbUdrN4/DcUdSjnCIjReObRYgs6yyyfx
XBvU3dt4h+hRlvN7Xa94X2+t4r4lQaQJ/z+nSTKwYdEPEpeB7TrlGByfjvAI4cq6AIDPofhqY765
FMNwh+3tTxD4gVQi7hu1PTu05khnHMSYa+Osm7Wz013MX+5t7aDuNX8VcsT/hg8umyuN26e7ubZF
QM3Y3hiynWWFIaVh8Ujzt7OCy71r0Y9OcjqKj6MafIJzC2FeLemnccgOsjDwl+Fc8X9MDE61ltQj
WaXe9ArOb/oKIwPAqZiWR/U3fZQ96uZxtNjT6jkUM63QIZdAoIIhv9fItQklh3Px18tnLovXtZ4+
zA7hNCeePDERhcje1LB9U7BrXdHM1d9OgEerJRij+tQam8AmmUhQZ6Fec5W1xlBg6ubs6FstSNVF
qp8yjKXWy2e5ZsA3OHqs6tOO3jlCqcMp0XPPSPUrmTnTWmSjLV3ejVAdH34Y7k9UuAnB4r/E8e0P
hBzeMOH/w3a+2z2PC3rn3eJK5JOqkzSNsU1QfdHBZV1s7kfyYmpKXAz1FVRwnETKLFUGjbJTyS3I
NyB7ImnQ4BGu1o5Kld8p620EdVXeAHCBw3ngpWsn31yFWxCPbmVQe/hIr8GTLm89q2JUmA5csgXW
kj9pvOP1FX99bbabxQn7r3wrUxhM1yVrnQjqJCTjuqLBRQiXJ0OdYZvr3BqrVRhn7ZKFkquze+Pf
FAUn+yAL4/PyHUkY4tkAHiAtCRiNTRCCbOb0jUlNMHoVc0YXiu2m4XKMfc5aQE4rrrvfCHE7jsRd
PXA1m4EO5owPZqGXpfpTRA1R8YqFypjcZuj24c9MNlwMXH1k4p2jCekklM4wdJbAnYH2jHwFFb76
kbhFUKtgMF2ohWNp6fPVcz4OVb/pPWlpLlOgM9+wgAJxG4WSOhjAt5IIHD75N7lJT4AYzXCqHTtE
rvxTPgW0YC2RS+tNgGd/7/mphQNKHevVRlNWKgl2cDGe2Tnj73sD+0xhbY6XQts5ufe9OCQolb2g
V1giX0GL3KKpiu4GyKZeRNoV7hxjDZ413oUJsCsR5F5eGRcFdzw/4ZEAeJNKOaWf7D5TpIWNRH8L
VDWeDWDnltiG+AROoEjq+sBIk0+zxSAW/EqOfEYoIBgq14AE5aNW9rOccqTI8GJr0l2dEmfTtt5u
8sQO+lv4ksq2YxTxBuzCLBLh+u+H/Z5hla1DgT7Dtg2C93WGzarOBoPH7oMsqlBzr6Sux9MTUuT+
KxUq4inqW7y/V0sKYEyh393Jcd0xmf739MOteatkZmfTkxQQ24n5JKxQ31IRZZyX+OACr8RAPiVv
HSa9df8ntkkXqW5RRpclr+vzVgNLU4dVYLJs/QtpBXNS7U0wkmZdQlFBmou0lNJIn33hgqlju5O0
Q4y6PvrE6eS/ElOfy/ECYpzE4UPaNbVuwUTDJp1D/MarVT9XMe+XBNL0K1Gg008xEnEHetzwrZn5
LU5jnlqhA+QtuqTWxzDI6S337feOickXpBV71pbzC/zeGfXtoXZ9NMxU/SGaw+LBp7brq+n0D86y
ANA1z2aAss1dIu7KwxIVyflVEWqDBQyCFkuP7MSYuxU4ODTD6oVik9hx4oy9ATb7FLp3NKClAxBQ
inIfEf/fiHjR6mI80eS882nCbujeq5wRtDY82fYKsfRKyunzCPCEI7wH88SRtOo4rD5OtreLLHEK
Sxyd9cZgF1Iugjybw2p5VNtE6nZyPOJlILzgrC5nqU7bRXyrnzhP2bwM45VrwoFIbg9ipw2iV+6z
kocg+KV7auay2eCk5NC1anWWB4/qTq0ZBmEPz+G8jpDDd5WP5XuQzRToWMko8AAOT5TpvRmZwYbh
R86CvgqSVp6n+vV/i8OBP5RbCvzVcsCeo2sXsGFrF8s4V2t6MO0Ke36m2Zxb9thlUMVxvkRw7awI
1A2eiXwkIUjQSlrGMBlnESkLClaHBun5pN5QDAVfa6SJokgmQrEYWSI92nKlbbMuDL8g7FiQjQ5s
WVf7HuyyGVh6q6QamMLGR4rAJljCTjjRQ0ltFkNtv2NwBtf0EJio0ZGagfDWf/uON0Jzup7Kwj/p
0+ruQiErBSvjNM+JYs5QGYcU1sGQ8MRCXMgQky7QnlLlxdmgatGyoGz86LOnvbUoauHIHg3+wpf6
0nA5f+z4sKfQUfOkbEMcBRlvaNH23U14/d07RKu+bnnFP75hTLekhUAnpFylMMQfxhzhkY+f9c2m
xyv17mCfHZGF/LmCJ2GIXpFd2v6Iq1PltPrq/GRb+YkFwyT3cpZ55+jOnP2AE8UC6L01xhV/Xci0
bFK/SMcIfAUiINBNj5G8gjX4tKEW/dKelaBvUOXZg3dRjgfS9F31ajSRM5rWFBoA0e7i0Xrn+7RU
9mwlxmNpSI4ghVUrbH6/1PJAqHLmGEGyx41/nOiuwPoZ7/nctNofh4mIY6jToEur8shV6N/5Q7fQ
BpqQ4g1z5mS5Bryv6Wmp3sBNlwMD04bWYdFiLeQITkMdj2yCocH9YHTnt/mXbhTN37nclFueC2BQ
DCa45ONihFlXO1XWFsKpliHR+HgK8iwU/Aq/ADWO0KO/tlRTje5g0KvYY37ULS70vshSZVvOOO3H
hFb207gwVFa4gmGr6TKkRuVAVrK3c2Uh8/rwol5sioFpsHKwgI/Rs5Yqihne+UB+/a/n0+MhB5hO
Z+Mfx2heOUUoXKKvd1LZpApIycLP345Dsfcvpb+gPhO0sPwvZsm16/YwyxLcSAe8qPM9jnDYTIZT
P1pGPb0NtFe6vsLN2Ank9RS9EVCiVNUjhExgVbWCTPJCxUyXpZ8qmBwlyC0usQnREbCcj7D+p8PE
qhGc18Og8m2v5ukGceo2J7UaT5wZaLz9+1FXJuopq3glsFah5BKP+dgcWzdfIHbmmc25nS7G76d4
uRW+IquYmESkk+uUakeWjbi7m9VY4j+kEmLkbQ14NwpmnTN0er0NioR6yaWWTbzLa/VcvU4QB1p6
AqB9/xE50NeZYXhV6K42B0IaOCz1sUG3iCsXPZGtO+BHNi1EiV9QN/nILFOieVAleaEUVUnRhSHu
j0jGDYRh6GWxhj+FkrJLCfiQgsjx5+A4qCZp1jvbgE6xAZiylIrTkgfoAPrd/mggHHII0N2xvoLi
dLzwYOJL6rmx0V8TehvTf3hsfLyut09dc2E7SxxlfBA3lQO+lwQWtLAHo8iJA+D8Gl2D3Tb7DtOQ
lZM73TtBYqs9YPENmqcKbzAj80YBHlvtiVOvI9gptT08beflEWfys9uc6rfMFQ6FDJcMeH6Dl1qX
Kimr/TJdZtCZFuZ9re8bgPOB1kFMl86RXTmLfIwAblEQzKcH8bARGgS8CGEpQdCRDqrOezoFsYbO
LJdC9eWMZMBsd4CUwTCQb1D9N2MrBYh3yOCufK8nq5HPxMyctmMHdU8gI2gL4cM8cQazb4qGbNS1
WkqrzUOk8m9qnWj++4PDT+ce9Ti0aUP39uJ7LZ/gKBjYKclth8zEEghfLl+bYc0GbZdd/bNA7am/
C6VObt9jaXm3KLnl1p3moTo0szzZioaEyi52uruH5I7mBjKiU6p4UBTieSig0qO149Rm0MypZqpO
wiPVjAHPs/wIw+3LTskogfpTvLySwVKwSoNIgIJBHz7ng2ipzodCDlnvkjavJoTuP5TJzfmp0ai0
y4cVxAchS9+09QwRu8sbG7p5gAqyGdASnHFJsossvKNm8t30XfYQMZP1PWqU/1YXu7Smu3YPQ/wU
l2KLCZpuEZyLO3Oqve/IeOPRhANCtZDPTPqZJ0fV9B2M7t7ZrBwSwhbfYTlBtqyynLgC9INDioOr
vdni8GVuKi+SZNqlXqKxZ7kqvfhfq0fVKRVT74KuXk9CiPJpxnqauAf03xJ0r/SRB0y50R98gkCx
r38VEiqK8WWa3IKQ3IosjJoE8ugC2mtSIqCP8ibh4dW5o6tXucYI1fr7HajJAXVJZkPsimH2ktbN
VuJKDSvtmko6RF+HR0ySnsELKKETx3sk461Kl33CNFWAk0qd9OyslA/FxegNduuroCJFWNDtEfIt
Mj/1A6JYF7c3SMxETO7RzXzXzJ5axK3/E/GS2PbaAwDr7LFrmNU7kHglBXe56MSVE4AHJwKpgC37
URINnNjnawxq7v89f8GC+XHXIkjGR2C43AUOCzpsYO9Di6FZ1ruu3YCptL/9c4DtPlHb/tSTuqGh
wRw5DtTYUoKSFPe2LSTS9c7Ud0G7bch/g1AGnpKxVK/qKPU6bJSHRYnMlkYfb/8hK+2zXynLm/gv
km2FRg9c3pt25xjFSxIPQwgx0Td0yMR/G8s04QZ0qcxfLRJFMFww6HQ58TsufCSv9+2XFeZM2STE
V6IdSCUwS0XdyYeu9qoXz8UFQcrcpajLfmoWCbZRY4kaH8rJA8C8qE0/d4f2MCuSxRW7gdlZ7qYq
AoId+NXubnc9I3OQK0wdZTANgmM8nXPOBX0fgmT8ceqi92qqrVh/FHvlD81udvuysJG9eT0ArYAs
tiHYfBioRghsi8osjPSkyE416odipQBfgh6UIKWs3fOtz/ieg6BjHlWZZde9tCKlTDHYQZIRfXtv
JIUXKs7/LfFml1IT/vrqA9zeu5xWheSO6n+oJKg2huM2kKS8/TWk140yZUoqG0xSISW0Bjx6MzWx
RSowglWKr8d8Trg1BLqQ/58QkI0Ot6clli7XF3DBGh8UMNtoZ7KXsVdIkmCtRTZ/4dvAx2DxfSZo
SoTR2buFk2CqRtYU5AmdvSBHBnj3HCi0PUFoTXv+7Zk4tJcKp4yEr+xP8dmGsMUDjiHB80BKfW/7
eDkbt340H3StIGzcsvMvxXwyUCysJ4xRieGUJ5iVrWqTMp0DiMSPDLpXvSeMDX+eD0W9VvG9mA0z
TX5SKAWhGvSFwgEHlZx2SGgYF8nCxNVtlpCZbuUnDdjc28DT3psCbmPo993/VTR/qztRcikowiqi
+ylIFOXd8mm0kMVFI0NxaPtG8sQ1y/zCjDp/wL4XbjAaNlFlngzFsvefhrVpcDptyRcRl7tEenzZ
qcmMe9ANl2Ksj6VvvPo5mxQDBEXQa0WF9T+2Vsns7AkN6b2sq3pyt2tTZT3Y8rFKHWYd44ivKj7x
A1EKYCptC+e/fiCLTK3VLc5pk/sl9xGmCaExtLJZ8QbYqXJtzH3jeC/PrL8Sr2tN6eMeQJnbz1sR
rMq4qen6SdJUWwumktlJnIT6Kc03h9TVirZQ9WAT6M65KmtgFiGyYp4Jqti+F1D3D8XIVFR8puY2
pYMvYBaTutnWmmDnrzRNemYgCFpnIQsPr3LLfMzhnwqtVgAeA/ajcBwU9lOTF1J95+zgobSMtWh+
DBMtEujbMKNaLxw4/pZ4u8xDXzqAg6edb+SrOxMucSKmY5/3m/yv7np1x8QJXWNY09rwjUjS/KZg
Zw2u5IRum0ROn/RB3pBfkrxr72+EzpM2pH60rEuYyf1Ea7Prg9xfzt0KuIq7Pj4oQpP/mezKb0R5
qc0MIJ7r1hIVQcQpNKyLHOuVo+IHNL8ql8YVF0ZHGUfKx7homYhDzW+kWk/xQoShi5jO407XmCDE
Bf1nwIOU6JZ4llgukdtlHJUcuUp/FUNzh/AQAA41KtRSOAcvJ/KTjtW+LVTJvKE5MweqK1Woa/LT
dqZ6D3LgNziJwJjIO2JDVOewiAKlWNNqA7Ad1+dKt6m6lU/b0IH9cn31piygEmebLfdxZ7epAHTe
6W347nHrMXFZG929Dpx3KMieGEyLWdFkMauNJe3OjJzuxAjIxHyUMLj96Blmj21Ew+vRASDOjAMF
txc3TwqTn5eIW+XzSAgykYmoH4wVWDuqqVmAv6Ck7TjuXJWpSDhiQxe47LKa3VqkZxAqFmThGJus
KI86Wieki6+Ih/VorlQBva0usa/8gk/LGZaTPfFayDMu9rMOK+L5QGjrloW+SvEFSUNDoMcgDAcZ
RLegQld3WQLqLmNsH6gjDDgdVk+fti1YrQMO4TzBnHk/MnEedEXd/9OB9zSLyeSOUeKT6ziDJZO2
2wKBvkYekp4+cmgvH5dZxBWg5BXP9xOe9CLtlQaES7h84/4egNg/kOPzpZpG4vCFxWaq7DXf/Oxh
0XP0k44GLGtVx+ZDdXdftRB4xqK2AP1CXD9Sx9JITnyRx0N35UQY378dmhg915YFvdfutuzoCmzb
HwKtGpmxT1F6xtpgyqwXfOCTgX6tcSS1jDDrJJco9YBaLIsxG0Vp7xolsd/74uSqMn+BTjDMQIWP
2YlGm8LW4hJIojwr6ZxGpcfHwlwP7QLfOjrjMy9tttsHVV9nxDnlw0Rld5h9P2P605YVv1Nepu4V
kB1TJXSYOWpX6iOkkflauLB1rsUGte1ld6FFElSkPOBIwlxXEKGt/PeglfVwVT/beDjfFCR7wMxQ
d55plTo8qPVoEvM7gqK0CMZd++/Xy7FFgP/MFSWs1OtlQBcCNC7//SPZMZHYSO44HHONtpSFzyTk
UGePJcQqdJx0I/jOYyeQeficbe05E232DGwc7GTSGJJcVjOuQUCidnlND3MTmh2qGkvB2TBo3ncu
aqJhkRH2ow4+1Z6t0KbRwcusSwpJn1lJYy1N2fvXYe75OtuzAxyvQgL8BSFh/kX+YtTVtq/J2jTA
YSCTlmS6LlCJRMplnpDjQabrSA1t1OQPBjT+KBDL+4PI9sW5Bq68ohIpt9Dv7X0L8b/gOHnH5rIV
tu7QptsylBp73oxa0qn0VXdYDtEMrsdyHTh5SEeQJam40FpJs+sdWX3d5BKpFKLeox9Oo9/EcYW0
9ccOPQecvFHYddqZINt18141nc4jaUk5S0pzePd8CP9XhtLlk+LvtPhDvv54abu9oFhGRLiDjUq5
ce2Q0+RdjPRP1VHTbazaI9TAoG+7B0mqH0aevm1xy6RMztLVglzGBrvfrVPx02Meqbrllb5a3g9Y
6/zTi4ky4mMqecopHEw8zy3q+1v4QrdaCVbHdXyLT0ZLqatwue+hCegF94HgAm+vuOW2NEZCkHyw
mi/tRI95FEz/pJp2NUGZzb0YMnlM4wcQfaUjJWj5MU3p0o5JlLnZWYJbKHiTyftR4vM0cHXBB7/h
8Qdri/FDCLdA/tIHci7uT6ZizRmfpiKBDbxVzx7195IIwZM3iowcQ8TDQo3fQKsPpy5LLE8yvW1D
grTqwKCoWzb77CAG5SWKjY0WGhFcERdnb5HOUI8atjwN11Z26ZTNGsv7d+hE35eZx2RtH4e3EqKY
bhc4oYcVGuDXjQmrSLn0tiZBgMbG/uGVASchEuViJH0z6w9sRgPAA8nPuYByB93joFmSNn2q0wVC
gcPhUv0FewpzJTO7DCvk3FR7mCJhy+EKPhkBe8659lDuDNWCz8FhtTUBu5wj7t60QAeh9Nn/aYiY
J42WZGXcjzjfF+/H595Cj1e0PfXM90cFidqMnX6hBFFWq+PwXJmm/vugxU/f7Gq7DWQDlkMMDNmF
trctsbYY4iaOrTtPLpluVCdRGwoVGTnIcYO3czpoW/uPVDmdZliVKDxvfLwicDlGV420GkuLov4J
kcvKm3hxdJnkpKBlwsMvCXPWzJsA+Q/ECBXR86wHrS1g4+0p02BwESeO0g+nstO2hGnEJLWDTZk6
HHucZhEDUJUdmcony2ywQ85w7e6ikPGIBA9JTTyUMw8DUE0kMZIhimXXwOIfkjal6khJwpPMZPFQ
2JwRIflDqnLTyPPdqkh7AC//vT+R/9wWzrRdIFtov++shPlc13eB/t6C15fLehtEdFjOySyYSkWn
bSUkHhYOXNeSQibGBS+dSWtedDVJZNPGH3ZeGyNHLjIAoiviOrVszEXTK4ZNYDFN1zVIb4jSKy+o
tfQ8L6s1PEnf6fMcU3Hn37GbjMBW9NrVsWvo8OK6ZDJFBnagw6uFGiZ+BGaXUvhATTBdemsi6UJ3
ZJlFTXnA59Rx8E96gPxK1eQdQMTYj9VVU7dcLWMamgeVsaEWzxpv8WkthA8wM7lJfnXI8sWNv9Gz
jLoyv5PXcolEmoZuioiWUFv8RXlAiijl87i48uwiSlztgiyAinPLs+egJQjA1eiKllkF3t/RQw2S
BgvXyqBQ71UY9tACspVPajN0BmipGeXLYqfCt73jbtd56B5BgPmu4Yscdmo3Z71R4vDzycGwgvuE
GDYuTs2A2sUR0T+QQ4rQ1RM1KPtgVVQknSrDDGyLiWkFugvTbFgZqCd8Hzqjwl+bjFVLPMWepW02
a0Ip9uY/FggR9yZgIHQ2/308rcxn2Os16x7kBlxfu05Ksgzpg5C9eMIZklj4+HZ01GKmYjLZHWxq
pslo5aehFYt9oy0ITJDm42J8zEEhclhga5qGCVqfCjW/Gv9DnWxzaYT5JZxuPzwDWXDTRqaQv1of
zDdesyBABhjtu4xzB5trMKXDnlKffc5/otNE3k0p1XyPUv7GjtXFJnNuWc9QgkWHijSFRDDTweaD
ykplBRJUfIIFwm3jb8rAw84Yi00Br16vcr6tCKxPMi3r+b5tVs2j73tlcDOVOkATs0JIxWfxCnEG
D89s1QE6FLpK7OfrrlCvncWXU4cX3hsLzPQ4Q2G9TWCXU4StceWtlXGXzszjqPyTHpY80RXuRVxu
axp60gnKWilvUg1tEymjP3hrRaPT2FvCp3c8UZZkz6KED82SGea+CPxmycparr+SIi1U4JgQQs/o
HOhlQIehredmPsr931jwDVZoVlfvotVm2j10sUBOZbbk8MPLM+EfEtKcEjlB24wXjfsqIBcBfjVi
ceF2oVFQBndUGySAysqoTCHONVy9vCE/mSQPvZcUhxvHk7LaZ3JCnMsIBwsN0oDh9bx1NQARXes5
de+Pl976PoyazAEhcVPitq+3GJW6UOYjBJQdnXjkjXzdEywg20ymV+JWwuOhTI5gTbOpRbUt+8IA
xjIMO+OEPnhoI+hQKERcnn8yttDHdLQu4/uIYCsEhWLKKV0aDm1y8y0U1djgCyWlTtsq/5Qk4rjo
joPGFZjB9YsZHVfPwJ/TjwbXoRTpLxLMZlXgJvNyhIQkAbO4wcVFjTgYmF9l+Dvm5xZM3cngTbrD
Gxp/n2G6pxLWn4QRugipjZCD/bGDIqBdPl1g5mq3d/FWzftay++OHUb2O7oBB4AnqQK9Xcoq35W4
wylWWEv8QjYTS8bjRmG/W3MqyEHFTcsW60/ha1N4E4W4v/YnDPAEVrYLby+jS5QBtyBn2gAAoeVk
Y0fIERGig6++PpzmRaErpG4AkYLxVGg5y3Spac7zJF1ODW5G/2lJBZzB1YBN2IhAwAPTnOR/z4Nf
9jF7hreamzy/ekMRzoFg+AEHBVc19hSjliEGxnh5nQNP9rYxzOJdy7c/vjSITrxfYdPRpzhompnZ
FfK36wMu1oyI+ZV/a5/vk3vM+W5JP66o/iA4ySSipZ8KC1LoWgX3tKQ3K7rjtnJGBaJS2mS7M8C2
kiTFrJCC0Z41zSuXDAG/5UiGFh5rBelFmK/D3dLuPesWqMEAkPUwpyp7G47uA5dLkkfPuo0TLKOm
8IMEfcbGhtCmtP+vEkX3x/iSVP6IgDEUm0UVJkoOaSdX3LmxcfEq2GGYvavADDBTUsYhfTA/ViId
QYFtiZbtY2oL5n7N6z0BxunvhPF1LqgQmpynd4PVY435/rsDydiaFsF9h+BAOmunMjb6kWqxBTui
1C3R6l+TtVnC8y3Dq0lpwmEfSnKdqv3W0kFBO8xb28KcokliKqR7rNXXmwlHlDyuZ54E/UOLBWWX
0jkXtwOtmdRdj+Y2+RgHR4UO7ssmpMDfzlnjDno6jHwAh7yazB/BqMZlev7G2L7uS0+cG5efk4Pq
xCzom4c1Zigjyom7iMFxlbgECw85qQcCVv27DGW1xc6qscisfQTL47rfnqS7XS4ZvwX25ckvVfw9
PRDiOT6FdiYVotknUsaZRbmYUEq0Dzrr87C6VL1MVTgO4ZQjqdzg08qbSZ6DswY8TWeOas+flloH
l9CvgN8mCKhnuFf9K0UAk55gRWgHYyU31CK5q5QRtqk7qy5Rq/rV0/d3lDFyAf0kQqbLixqV/B5Z
Pz3XBttyfXTkkMnb9ASD4ZqOxSDwAvzueFUUv3qp39AilhAQjBUazHXrqINaHVa/o32mK+wpjZ89
EhGXHlKNcJcKJuxtQGcXdTeRhNyXhDHWAE/d0znfpJoDIz48AogNpCBBC3EmVGCfXj/5R2HPGX68
K7zRLVxqIzxFIG9H6c6chzkKFaSvk/2cKWZXa7UOU9yilojEszjgjW7UU3zmbhkLOXSRBqMPUe7d
8aRMBxGdKnrloz1MzKte8H8owcjES+YK2JVy4zRVTI449wzHXVHysEEqhlNtuZ2fIs5lTKAgFvLc
JxOIt9KjVrqKxlK1l1Z39ngcRdjZJxvON2Pgf+fZY76IsRZ3QAPVRvaONAU8YTaojIXy/dEApQXi
t9PWQ1wzmCBsfoRPoaUI5oMRfe1tK0u0H7dufyPCLyEEKDwXbZMi0Q4FAj0MhW8lglBQ4ivO2sMK
fPjY1FnO1vtOWk0C0vsPbj7LKwDMZ8hpv3QdzFoC8cSsI6KvmgaJqUWHB6UZhvTeQyau0Q03ZUTT
52jGwTPMh6NrZYhaieTybOPPSorQAB/GYeJ5I7Vi/63jukCbpXUzmLKP1csziLZHjsJEJRcscKp+
co+EXA+gLxuGFtsYfNNB0eLQgmmMY6uLRJ7y+TdLFBKFzGxzBmyL7ljidLKrDGIsCr4kdSqmKQmk
27CxM0a/Qi3+5oiBrcOVnLGIe58Q7LSSPNrVzHPHq4TH7T4FE7b++CR2c38/P+ufwRTKfA0r8DmN
3CXfrhraUnNLR4ePzWV5YcdlrS+7t09Sf0uPkfcQyGgbt3cDZaMPnEPcOrxuSW7Gmy47vd4aPd/P
tRmsS3doNte9CceBTek/Qp/at9erBz4YpF2DoUyR3l33RLYKr1L6wsaD8mE6Sx3UxvRELfyGLUGq
wEMKQN/6V/sJGY+fKQsZycjuPemrKm+0J8SWWwa6Z9S/7CJTlSg831TUKxjEiPJqFc+sF6rrJ74O
ZB462ebKHLdSvfFnVCuyuagq3zuC8TnL0gqfwKClMjgZsMyVcxHHeUm0ev34DaM8orkcx1Kkuqrs
uGl8Vjw2Z1UAjvsIlrA17qyePv8sKHECR9CuATaXQGC1R1hvLyFAidxr+DqtNJXoO7c6gGBqmyYm
4PDEueEQ80sEVB2amF5MVOn+8W8cgoh2iYNmgZeP82cNAMnlG7Rrsmj3yoCUTVF44RqT8a+jrn/M
UiqdeKCuTezOjrJO677+Z8/soOeJdGXqMvAHhyl9/DwF2yOrZmXLEq4Z2E9BsDLxQbCYoHOe78tC
aK5ruaGMhgkoPSQzaQA0UqR8PTQRfJrp0pIyPxkwBuvTK0/Ik4sgJw2F1kZj6NCKLSArVOXYOLKO
KlbWPJvoMmwOkJWHuHowz5wkudyESzweo5q3TKzA2GnHAzKq/75L/sdkt+AYzM9fmxwJP77XEes7
lHIp6p8ANoBvzC+X2Lp00CmdSzdsvZJD0/5xzGFQ/lwFxLWdRGs0+p9ynCUbBM5/w/9yULT6n4hb
qa8RegdqeVmgvDVtVuXSobkrq65eee5nWuee3oIahW9TBLXiA4Mc7XbenzDyCpQnlWSdUrO06CJM
nDrPEi14drgbqPuHLesq2xjugcGCRGkdL35H1lo6B/YDPTF2PSHi6j7oEWyXzbiEr0WB0+Gm7ZRP
Gyd5pUC2zEWDFCJTZdQ+zy+fOqLPqET295U+wftNzDXjoTqeYThVSUmcNuby0aqtP428EON6KfRO
Gtf35jOSNO4qvYqAUkpl95lotyuPdoOc3AE9pP++zIS3kTYsf2hgBiwkJIo/jHPdQrSoOmYC5zWI
LWWpxU/N0TyHLvnWO8AyRAe/UQqlBqqR2AK5GPWhctWpO4+XHK8VUjAGxItaIJ6KRVji7uZrcrQE
WJAPVKFBT52sxLzr61/rQY5wCbmkyZiZnGkLtWLb5AlA/X5T/2ZEhwn1z+Z1Ok3IZxso6tIRLtOt
TcX5DGyxWaHdTOnvUA/GY9BSucK+eNFbjRugP6BNwXDuAHtr+NMPYyUvjzfuev1pEpG/yNygUQ9F
HW23oxrFAZXLBQsntADKZN0D820Fjmo/r/nIvZTQQK6dMIhGNEHmoIKIeurPbu7zIdDrtl9R17PY
DPVL2QpJ7Aaod4PwmcUnPB9PUocnjy7dByuETRzWOzdw59BaSAzJUzkDRnDxh0AByLHHbAYUABx7
Esqm2H+OuuKFpeD+LQ55TbgoedtB8CmYC90xf01VBV7tnWWzsd4dw7vto/Wsoxp/izoPcQ7xgefl
JuZ4e8oEJGnVp54Fi6OZiGHme1RY2F1+RDeMCzVv4xKC9/w1NJbLHHI1HpS/66HD1XnwP8oN/yUB
gjfO7LgpZXi8uGyw5UR/GGvxqf8P7V1TxtpqUg+GugQZBDmFW7R4YPINQedg9HVsPjnlL5eVM0bW
yZyQGMzvDY3sux5oSzx5omqVGkIPdgqIRz0qqBYiotoZ3fIpf5ZZB6zVMrPYWGEtrK0qc+L9g5hy
uXJXXMJlQYnT9f0glG/CLuqd+UsY9nESUERE/ATvLmMdEaPmz9HRR8T9/v0XINIPwQim1YZpwaka
EUnVhGY+m3Wxvhtws479SkvTRLc9ARkT/Bzj6TpCErMbO3mwWah4fd0niMSAFmVoLHbtbxkYIUx1
LgyzTrRBF9qN7QX11nqT0OVS0k7D1gZ1kQ5aY2+rWf9fs2ZTbP899KaYRMwbhndys6eYT1oVYNAT
yjBjEwT0H8b8MT6IDuDzFFvz5gNiv2v6zyvL30iqiHbNSOxGFfS4FcQ50zEid9OVMZiHu4Dh240U
rqC+Dh7dl8thl22pEIgpTbI9M3eN7wLjYJcKSE8F3VX8HrETOfWf3sE/vJycNJ0htfQ9hrucgU35
c/CzcALcHTFfYFOoWZ5z9LGG7WIrd1r8vid1pgP++Sob2BCaTe3P5hHnRSmquQZ9q5itQXUVyhhH
usFWuu6Q1Z/AOa94X4z4FlLz+dLFZICdZl1NDFKFloVA6HA+DCUhl3CclDDl9bSNAAX2gVOVDHx4
0lRB2Ba90lnclhIV8X5qNy/C/JJCuEQ3C+d/+kVjVpvtpDF+Np2/RdtbAIgXHLn1O4qOJzLENu6C
MmxtWvHz6TtEXF7sYfscM5mlYGdI8sv3XQAqOaUPKmS8SOT4fOkJcLd8Q9pJUWRlBAD9WGMd2+wu
qOCfjo3Ji/rjTA6UspILJIRG6FY+cCPRrJme8fZ8iP+3M2MHiuNm0p1V7VliS9983MAqQf/3WxTA
cIDv/ebC2wWHsb+7iHlBAW6rKTY90AKb3vdwzw5x/LdiXdWPKVOtwVgpV/r7YtC2laDRy4Dhgi3O
ksQIBJN4IPUEs9xzI8TEP0Evo4MS8BJc77S0CIfwGlNUreYyDLi8Yk3uMzQA52eVpMZd6qCXUgH1
eyo2x0be35Wbbub05/IBJZO/J8jiFljAxwVYbaMOT9Nc4sna9v8CoCoKXWBHQouzmcOJZqDPjj7m
JGLPOnHPLPzUChpxP7028ZjohlOgG0gz42Z3r/pnR6pL/r4EY8mwnHBDhpCFL56o4anML1nP0j+M
XWlztggvLaA7eq+ElOC84wHqazdy5k/TGE03RTtvYRL3JwRjjsu10mtXKoaVPLMXnvTjSKi1Nja8
QpovowyapZSTQ5fXpSZQtJKkWhJ2MzNapTKyW09EhzH2tzxPVCGDFcz3BjfpCFpQSh9NYKeidBcs
VUCvrA/qpEy6jcNAiZ19E/rn+TgBp1xCfbnpKE1P+33oek4dmcjZurI2avpyLj7IME313gfzasKc
vEwQ/K8iJg1ZA5I1tENif/n34xrCT2WVZ/64Z45swQJTjOWdO4er3f1zl+axDeh4qEHp+QUFKUW/
+kOsfokJE+tYtAlTIAENsD0NgsvR+CePcp7L6Vq4XFNcIVbWL6t1CmyYxOlr56Cj7biVLsaSOEuD
C/BEG0yNBnTZKMXauBiqurnuu6TTmN9E8hzQ+CssSQG71rZ4vzYJsDJQTsTmfHPk8HADdBrkQLrL
UOzsdjccwLZv264nAX/pTbMG/zRfy+Ht3E4cy9gwnvb383dJ8127Yrq1ELWL7OU8AUi8a2zdK4KS
SztyJ4B6mbLQaLX/WvT9Knoedp4ePlSidPKFvJh5k0Wan13gN1Ey2x6thLnkCG0tBuN6kms2vwyh
QNRK5OCZTOfwLVdVEjHitmI9/bJok6HryEgBdA6fUwDl1vCPv6CNlLyuMyRgnDGBQShr4gv35S+Y
/wmtMjFaKXR7TM8RpsFYJ12jTDoPBpR14Ji9CmJ7ANY9MIecxo/Jn9BPanrgrvEjbRGDQZw/wr66
xWxL/kba26VNQYx1FOHKL7VzYMTBfK69e4WnsfiCad4BDAAlghQ0FqwnjoxSnAwj0nxphXpeHdk2
JhE0QWkU/jOdcJm9dYLJkU6+h4HiP2n74efP67LDnzBs30tAqPvwclCLv1Pra1LeZ85sWtzTJWFO
C3N0DGlI7neNVn5L0seuaixa4rP7HRQteOKrN4rkP7iZPFYkr6ZY0q0O7f6WFRrhRC7vGm6bNQkx
7HvwQ2b105FFOw1FPY1Zgd5ZNIpPJFKrW8MQDTJlJn87Ys0XwzUrS5lt+RHAajtX3Dld51h7wlD3
J1/m7DqjWV35TLFrQkn6diIDOy7tiOPFK8y6UGCISqo6rz0zfYz4g1nn7iGpbDRVxcTpV7NyAgge
GdPicoYEVxxtX1CCYY+yq6Wx2MghEQ03pBe/NQoYtfWAENbAb9jmlTpmqBFT+jF5Wm0ZKWWtEW/R
+PxFO6YweLE6LAO2t6IW2xNmdlNorV1+c98qYIuLW83GJIVqndb87nANsoC1PutTiXO+S/8/Bnhr
Fvu9b/EJdY5AuzFaZ2dO7qrSABUvTBMaEEeSHmf95CKRVxF+4RZmkv9CjrICIgM+xRGV0wNNRXug
cSuWgG+wfWYGohNb2+/p3M/vCbDUpZxtpVA90oaV0HCX5tqXDv+HlxAy4UsQnaDOdvLZQUHMO+AX
J3enhsdnVqJRz3S+0avuMKRRGie1drVftLOnD6VNTi2o3v3DcKjPCSWG6EdXtTlqKpuG5dZFUykb
XpQ/z31StcOa351N/jv0C/mEoEzx96A6cVulxxDMJIUHKEMTlQLW17L+y4lH9Df67kxRG3OXIv4C
epHez1J++j5EUlxzOVmQtp8lVBYrXfK7EXZJdy2YFpEWsN/QhzEMhs9eGS8jqvmfKbbHgG0V1sE0
AGhf0t0xd1efdc0tC+yLMUahGWJCZydEI2euNznCJ6miSadKEchykD0R9e0fMm7tHQX1iCx/wPE8
zptDZysWhmnfhfCTpeSMSF6j9dFu6FEUFtXiil8FFbU5nI519By+p+5DJ5VxGtJ1IBDjxXWijX9F
DdGXEB8s/wkq4jNPpQG6oD0snD1XfGND6KXDcf/n2mVsNZ8SdVdLTv1vOXL8DJlgjhozToT8SwAn
GVFTEDJIR23/CbJzC3rhYaJTpuSvKiQKVo13YJxpQpYlMLUqcYNGSdjshJVJ6uPTl0GitFOFWgHz
FCGhLUHnZSzc6V3BW8P0wQncBSs68ia2VAUHdfelR8Re1Lbbs6DXWmJFbp+oiTOhvkJGoAuk49Tf
NWw+xUnXKnM20fkmDlkVLXlBo4Q8V6CfuI5d/LwqcN0pnl1oAMzG/48PVhIIbVxByebeXliNQSGj
vN1JxwL1kA31371sQUBOQs8FYZ5Y6OheL2Fg/Ee1FLm/NDO9wnpabFXy1XdtC37B0+s35UaGrQ0t
q+x67gY7GDEoRO5llmYv2/+yUH1EAZl0ALiP65uTm/hv7AnSqjIVfRaY5yLm1IONxRUvLMiPHtHM
BGGbL1OTAR9lgauqAn4+qgLX0ZDvsWaHVjC84Hl69b6rWj5E+/Elgb9MZboT/4crEaOFCXUgqNC5
apZsq9YhSLgsfky1rlZ6f7iwBNgnNu2KSoEOsqA7UdRCpYSJtsmaN4vu1MfGIayntdaeL5atgo8j
p/DUKcdeWZNpKNHyZzqWNZt0RwDbDXUwFadl1LhLm+vIU+aomCG3YDZkjJgrKC6Cpe+oWSAPCWt7
r/J3vIWlyHaj35235g4/bXiY+A3CtjWbvJ+KRzW9F2qLOU/VDnLYG+sLgO+rtCZ2X1EQCCJOP3gx
EDgxbbfxcZekKgB19ehZt3pLoQbejTner6nA6Yw5J1Ie3yfZUkU6X5KLoMDfMWTrxLSWWp9pANPB
s31RPBfzpm7bYyXppXkN5M/uw2Zay2bwNc1pv332aLpIJRn0AieQCz5JjRe8meg6F4Vui/5uGPJW
aLMgp3lcL1VKEo21/dRJim9K0M0E1YiT0H4hgs9LgcHzBHN9TBpvs0kghiVzROKz2kVa5+EPaseQ
1toCkkIvoS+4T8B0PfSKIyyZ10oMULzp0AZOU3LsWdKWU9hiDZTuKRjCq/VDX0cDc3/Udiv2i/Dw
lvYjLL3H0Pp4u9vewTe+jWaBSxg7CohLAuWER4PQlKSLkc7PDpjSjXhIc1WmMBspXVZ2UYCUC4qS
nX+qzxwXwN7+Ay92e28hp4sYi3ryQ5uWI2EwBLpdowVLbo/CKjN3ej8s6Vwkk6mmFtCyePYKFyBh
kabyKj6RxdE0g0KkZ+YJ2dr5gyBdv4YNBZRvW8vKR9R38Hjsy9WZcQKbn1/EXOBQ39Q850u//AU4
YowXG/k/p0Nx+Ney/xv2XLA/iaPHY5+40h1hiPy2fcADxEBvd5pPcC7kcZto9AfrDONQdqFe9iZB
Rco1ZkK1UIRnD9NbL7fMZrtGf6wn6MccVx5XX8UQ/BpMWkNmfqaTgv7Sr7kodZfNT0ka1d9eXRQR
VIR4K67uylK+M+qdF3Ar7eiyEsMjrd/p+7yuepMeaNl1HOKlERKqdf0Rv7t1X7lC5KyTM2JMRhNC
AlBtx0dMR38P+5lZPIIFRETJksbOlnTWwGa78htCEwsi0vQepoctlKkul/OzwWt9ido02kYPgxYk
IfGKx6YKGtE1C4VFvkHE0FGXxUWOk3/WSahlA6CStN8hSDxibpgonvd4p2vp5Jzxvy11o3OreoFV
vvi/FZxM8Lxzp0Q5hPAhMmELmOjQtnw2ekmd821Qp5JXDG2BVBt+ap0lJDe1vuut9l32dPZIxZ4U
Nfj6wMNljRE2kOWa9NDXMq5IEf0nFOVNwANc9rSy3cpbomT0mKsERPLIHbKPIo0e66MagEPOwnJf
ndIrf6ZIvYhJgvyPgsS3agBwhXSsN5s1joDROEnNckNF5mNFlEuhYli+jzZnn+PrpBnX++gGMG1M
Yhw69nDYv3usIoKTwWpCzHnuLsEP/nsJaYjICTerjfqybMsrov1zQNXWUCmVC4LPAcaBuIN8bOOW
NKDcnLFeXX76R1goD9E3gJ8NJX8sSWJReDOPzzKCTxWUhfT6A9RtPQSMaDp/4S4RX+IZWYKmCEkA
pdRPjDtoe2Q6DQqxkT8u7mwfIT4LlaofiJ+JR1Uc3M7c4UYCtFGpMk6/3gftMBVebzBzlNf/hGsl
CYZ9kZk7396THZwwpCSBRXv7lIXZdv9xAxxU4iRRlwbD0zD2OjFTyC70Xgm1AildCKCkUbfQP6xd
zQjVf3ZtDz8l79dQjMz+6EAgcFOT0w0fiETI4pqegLIv//EKEvfJz+SuKx3MP5Ml+x8ai0JPQ7j6
cWujFZgdU8olNw0sRImTt48bruIysZgGaNIr9K4fLNZL4RSS71A+fXqQkvQsL43chrEtpv0qjAcL
TvepU2NLaRgVGuxjAJ+fjU/HXQQWSaDvbUVZ/nZsf3JaTGEWhWZjLBscDik+XNOQbUSjZp3O12/3
VCKGzEYFU4EOpwrVxSq3kcMbAuPoJgzAkhuALbY1YhesLbPpDNGTgh8i8ft7K+XCnyVpfPX+rdST
ac5VR0YZpdCk9q/6A2WtRaY735OBEDiY8vNX/GX3zzXv1vXta4Auzkufl6ZF0GgsiQUaholvPKAF
e4DpvDPSV3yS9zSdiHCGRs3nKHoGX2FKxut8clZwuRwZlm02Ixd1SLA96NVXfQyu4v2jOnDYaxvF
OLeUjizl4BxbXe/LGCrdD10wzyi1vtB6u31D9o+AOISt930RN6b2n3fCfePA2IH2zMThapqgSTqC
t8rhGzJYrwr2mE7qDqMYpRacQVvLWJDy7pRpYA/RpWrgeBM0RM9zS+RyPRbB6D0gAyl1qAWGQU/H
DooZ6+5OJRExEd1JxY49Aeu3wZKXOYwlnnYgJ6+wVsvDjJbdknxZkiXcbmCzmDcXpqjeHzI8XsDa
tEuESWgtbBU0vOxgjSXdOzre6DolRy6TfT7Ex1rcuRqTW6ypZyd6FNAaqpc7PiGPFxMhKo+SlIjo
paGSQGziiCUeEo+f4Gx4tucBOjwkvxqKReBlJIFMGlQ++6CkeHUJ5lIm+skznO/NAdwRtJ/vjxrG
J8X/NTqrqeSDRKgOKhrmfvM0xlFySCsyyce8xeXh+QBcxBrVn+a7wx0rOnL5wE+fnn/slhp8Ve1K
IkykEfbq258jcugu+/9XdzKRQg+FIcLB11G+yOCNtCMNdAHcvbBHVHH1fMs+rKVwyhfkHAxpF52M
gw3/7FJDSO36zncDFXS3so+KxddtU4kGWvZd9MLEe4DUUjpVWgMsJJhP36YcM2ai7xqkpcrsXyRn
TBp0/PtkcqtsT2O3Rn92uePF4/eDxGcBTlnxk45dSbIRV8GtZB8Rc7IHeMPFnTkK2aGyGFwM/Ckl
LZSD+x0SHzO3NpmavWbSUti5XD69NJgD/FnCFw1xg7+BHKt6ZC6WEYmL2FKbtTq+M+rhW05e1DET
b2kP85Wt2UWREjcKH/z51pW7XFvlnIHT88KFP9Uolp3ZpKRP9C1Z5aV0qElJ4NWsSE5tCRrVvZHX
t7YB9BXF3nt+JUfJz9j2ovfV+ltF4m8WvanO2MXne8CK3iSu+mx3Y3tnjdnVuaiHXjm69XlIpr1a
O1BvFSv1NynFoBlOlvV0jajPWiQERnj9CsmGxkCeniP8Tzo6C554P/151Vij48ADPeKsqQUH/CQa
PL++mW/P5GeX1anxFSxIxnmDPcji/HreiJA7kTs1K+C2Oz8LV3Itt0iIFEMtJpHN64VHJiXMfmoO
4BN52q+Biigr1OUi2YxPMneaymNmK526QFWrJ4cmmZ9+nNJ8z2UXb/txHS6gJ50dEMM76Y6hSopJ
BUGhyUsWj/5Le5wItFQvTlE8ConnoW9awsfYo+Fu8JdXZw7tOUC2aLjrhQ2MTqFDQLcVd7y2MfhR
V1a6O11p8MXumFNXo7ejJ42xv/vnlxm29UIZCxOoPVNaSKBtMBTLdK0w8badFYVFGn/FtRtpXYeh
Xt/DjQeOmUllNkN1/hxv3LuWMOUwO8v+5x9dsGE4+ZIhPptq3pL7u0TgOKLlc+RTk33MUiXRhMcN
/kmQNjYDPM0rDDpgYcE7ufNq/C5L4jLMBrB8VotEczocl9sqFcQkw4ChxMQrzXUoUyEnm1QLpgFy
F28R2tSfKKklVVL0hE+DlRAottt9ZmVfJfSscdm2IFOnGZcxbDcjnBP81qGSuKNZFULcXNsf11v0
aAIu0TRciKvDtKTnRDGPOE1UaWUh8P/YmuPZwcfUMEZgupHnNoov2Sf9wm9JdVYq/+NaYteOmzf+
fcJXdyeAB8yOfUlY8CbvncF5S0CpOs7vRqDyLuvaKg/trSfC9yCXYX/cK4dm0+0e6u9QZGyb6vhc
k6gGyDIwycoHiDliPhrlScL6HRxqGoD1ynv8PHaAzChkRHDsltCEIIvvOZrJpqK/+KfXIXozKWBk
kFfdFuLEDKwfBx4HmhWwIltCmKNUSW4lHN2wiO0JbhF4QD7OlfhOgfmfFN+dKjcz/uAZcPF6AEhE
mknmpXmSOZBFduX8N+ngD5ufjBaaTK6tdqIUWzQ2FamiYcR2/60FM6vLWvN0n9YhQ0cQY8wq3Ywu
xAznhHo9YRh2n/x/i7iuUNbmbBwzvv+WcWI6DCpiGbbTEclhLNfTH4StRtekzoAxDZz+d5odvsWs
aVh/rLih8M0p99Ub/WhYtsnHhyAlMYw53zXk4ZvcIcOMohT1fR8i04ZTL6ta2k3hP22U44lxbR43
5TJt/SAXoOHhdIzwUsh0fPxYBEMVNDN3IK39mi5jJ316Je6H9iImbqBSGxduKKOGelf39O7sFKJ8
n/nmRyBGIXvUDY0kS5J00oYQJdz+Ol2wweVFlpwHjQ7fWpw9LSgGNgLBq3Dh2rw0HEkgg4sFqHpo
CHLm2iDq7eeU1eHl6u8pIP2HSfdBTrHuLDMRjlynRH0Scb1b6FSeg3/56HssR0vxSq8TWXUGj59o
uq5lTBNd9v7fgK4epRf7edsHGHmkjui+NUUA2EoBcZiy6RHYb/KTItXRBMmVLx0P/MQayKWZnZdb
h8H9qod5A0YzY2IBKd9OOwRZ+Lm3YbaGR1GsH01gzIvGE1oU39bA40SqJS84wo6PpT6DsgwWepu8
NtfLKcfMFrWtWJN6Eo6tJMB4yX5u5KE9/8NmFqKrfhzpSj4kZKt/WEv8QBXTBbNHJcv9Dl/dw/kL
367PZXUHZt1EGsWNFmTiiIq4v6WeppYsQbyU1MSwS93cVfbcqs4L8pDyvwE5JjCIEhuVlkwHmr1Y
msT9Tg6zcwBhqZyUprrfCoYnrMyMlcLotY74qS2ttreXm5bIGjqYwetqvhBtv4ZIgfWfSIqc5PRy
BphXtDyKYuQ62o5NsF5iuXZ30TeNTdx6eHWRQc7zqVSY7BfBMHPoxwuPLOV4+bAY3HyEvdDl3sNB
OXeevFTmyxmNyXYCzBv3rs+PoYCNsC2sGj70pp6vsw3BGjqm7fG0y+U4q7tOn/wOHJwAMzSG38Zd
HZkYBfeUi3n/bNcD6kdGgtRj+p5zRcDIVgUO7+WnCpZkz5VbNA45soXWA8KQ6pyu3mU/7hu/NKxr
R6IiwTgFh0kb1KRcgxfM8QHKcp1zkblq2RX36+6WUyX+NG6S87O7tkJTWWRntWlU/+naN0fWwiTf
sWpMR/7X5NePGsxFwMcjcmr/krxfUzozUyo9njbDOIh3LKVGJsZp5DcYhTxND7ARyaJNYG9FofET
TFh24/dHCFdY3b47DGOGhIbvzwvmgHo8vJACvfEADTjDa/UNhaW8wchaSGfVVHPtlPL1ORjpwqg+
ndzZWz7nWTu7KxTjDWaTJBhOK3AJMrTOtIoesIonv4JeD6h1c4wB1SMgnDGUyp2/CPbMfy3yYj8m
CLV0aNW+c5SnGI6TDP3h8bgy6mDVz/Jb71C5mEbiQK4InDHIXMst9cnwT587HQEhqhzmfA3qi2Iz
ArUNlE5DM7nPd7gdefVetyRBlPfnz+ZSVhGnI9Zab1ywYyAKIJJL1MDAIXnKKyTkyzS3xXM97QCw
lPsE0glqCySz3BPBuIswgWV3U0EaKyLFXafv2hlrk0IJJ6yk11gp1zyrI1lc9cql592FTS3kKRYO
2vt3sEKjAVFUzDdo2t7ZlFszkcAkPRwCScr6SW633dI2/g21UCWHPBPci3tnrCzsJX9HnJiTccoq
83W0Lw2468TDdl74cW6W/XYk/DmG5iKWkUdaK6YNDpz5qFQtfuQ1IyYTb38m/F/PNqiSoRprKKbN
j94a/tHFOiZjHBAJyE7XH9pWfzOuDngszgt8IfAmRRHnEY6clNRU39A/TWiQbL5p5xrxuobV0wyn
I9jhw87bdxTaPclMPCKr+rSAay4N8p073IkX0MNMwwqRHNZzQmMgaLS8+Bps6YYYOa9sLCs1fpqa
HC9yfLnP94XUzyv1vczmRnF7x22Bv1w2Ri60n3R0FdBkEJBLfNMqjtMuWhFdPG5myNIOFXB+anak
YzREiV8wVH2x2w0t/gVl+E2p5kBBu0oNlP8Nv9qT8QIZyGNwKGJsUxww2t4uejM8crPSVdfK5J9L
5eOAy2NU2foCVN4LevFj0ZQdkR96Pip4hrJIHOR4Rj4o4unz2t6vVlVwhSe88Svb4fCm2NZ+pRvi
rN7sKYkxP1g1SvFIqakvmAnGXvDS8BTr1m6PWY1t1pA52ds5Tm1oEqyf6VEpMyqALHhg4E+inhJz
UaHMpAuwwBMue3dpFJs8ddAO4m3OzQnwhH7gguaWf9nbl8dyySRPGemUxjiOlFO1NMzO4Jm0SnJV
1NzGywv2AfPDpwvh7r3VuAXEBHEO+pjdKY+sLgX/z4GPiSfOddKrvm3cdfxnibanQeK7BMo5v9in
UvxjhFA9Ox2Ulw0BLQlH77J76Qg05EgvEkhTmcsnjROHIVY4cP5z2Vs2rL1EgkcyvqC2fFzhGSdr
LkCzHo8Cci5hYiwEEuXra/lVUPzquKUOegZ8cR3XsdBpkrk8tS4OL2VY2+933FGekWq3h16PzeWn
jo2auGl4XKkl75JwTzi7h9MUSsM7BYOfH9ENmmKaPCfpJQxePlXnyVPayWzJaus8NpV6SrKAUJhO
+dojdnf4ZDrTuhDn6fGN5U4a3wm3y25eiunZfqjRSSPDIVJnqKm2oHBRq4x1DfzMtrqiszQLN+yE
X7xLpveXrHtKyZw8PHiP+iP+d7OGGp1fvZyguJJf32YeNOwE+sVCi5sMG3AKSZqEEgGJF1kW+7rb
2MWS278ZOv4LEmHj1kd6FiobzKkbqjMtfaswuF9IFx0MaAu3h3U3xcraBYg0w+TBG8v3wgMSLVZ/
VGv2dSm4NjPJwhCtwXQ9Inb9QQwEOjZ4VCd0uAZDWBaryUdrpkTE+vWRwwFptvGS1kvldQ/2Zbxg
k0HBbtx/t2m/Eln6gb0MOh+3HFCe/9lIMPsJdieXN9/IDvkXGilKZEvz4REh6ZLJXModWxkiJ90E
NbJxABGHs2bg/qoYwMHJayLmOday9WiU8W+4rIEMCkucDqhH6kAZBZfke3XXBEcmulBujW1ChIr/
TuNZIfS2UPdG/Edchzl4WxhqNzm6CMnJ1Xc9znLGtDvzlaYPpIsgu3IrVRQ6MiSz/Y0dF1UC3mDu
DDc1iFAnbmP3bOExZGSrwoELnGn/wn32M1alb++WuiZxJQFm/SyneLoS0Ilce/THBlvXdFOZ7JVT
eGYfepALap+h00DBwkk2jlw8d6HE0BVuS9ajvhcAoMwhV3TSev+XWtbQFUx2eujrwqTOYuqXeWnJ
CQCzvpVp9ytGuR4znzOWUWnX5ynyuC9XJr/Ud/dc+BUgmK4ZVt3kGk8C+pjx9KiPlZ0eOzDhnHTX
IxafSP4Fx9xA7Z9GxhpPaOa+KPDjnin8Q+NZg1yv/jKYwdn+qneQlybDeyidOu4yOMXuQdO9jAM2
QcwyPeKri59m/4UbdW8j/toPTwBrvZ2Zn+mdcMr7jfiWbwfW6vPRQWyP95/H8ZfbOfSlViGkpmhX
5Ts7ulnk0kS/VFEUSZCMQk9/3ugfgAaM1ZY1hom0/fSJTCgdsJCHHSv9MajV9ZTqCce/e8NzJQEw
B/vnZRr6WRolBz//YwC17AMr21kGKy8vvsWC7K9waXfchFBIUn9QYCHfp8xzZvlW6CBum4waLK51
Wsud4PDx0/6d1t6ZrU+ym3VJLi9Xhk58aAzOB8XPdHo769XQf+JN1pNxOhdljnOj2pa8iSz2mb5+
1SJxcQnodV2mytlTD28dyoQ3fTskA3qoAxUhIFTeelOwBbHK0IGrmL5twn+KnRUA/1hRFka+Dv8R
N0KjKp0t1IgCav6UqbjqMYKrXUiiPDkdI2DHHO3XXlrsHbgYG7eCM1wW0A0R+Mhh47PJA1uR5Tjk
DYkcvZ3qVGTPhsrWfH8i0dSj03NpoRdKmX7/XQYiDBFyi0DMAM70SP8OtkM5o3mndP5fgRVvk8KK
TnfGwsmy2w0ToWncRyIWIpb4mbnarka7IyilceqcC6efkLtt0Xt1j1qVkSipRyFa3udRzl0/VZPq
wVnDZhDBqaYm+GOoth4Yodre4iBPe760EyooxoDqgs0d9nH0rzLs7dw9f5MG8ejtAltBwNT/b9l8
iC9M9WKgArP+f4MlWhRQXc8oQIw3d9P7deouxDQAf9fqXC5ttWhrrCl8+baWGOQ5RO0CczcM8dlw
DB3FYUfQusKDrpzad/RTvk7DP8/lfF188tPNbruk22US6BYmILokItBwCC66eaR1+V6eoIDkmYVL
h80ao/q/0i+oKtIactMC9J6+sY9K31orEgYclFdGrLMzvuV5PsUjhZXP4RGMW1aUkmfKlxPAxhdP
9SYYK1F5mUBYrAwC4YCpImlOT6bmSmv1Ry8BA5pyj3k6uRnR+NNV2+tgDL6wKxIfqoDb1E4WgCxE
rFVE4nES9sKnRKz0vEGxQjJYbD5y4v4mOPtUVWBBfLGIoXjpKyaj7qCWEcP6kW2//FBxtSrgAUs4
qiQaSHS1SF+b37hKPnXkcjWF74XXJWNXXgUpfXSObWv//BlQWPg9Zxapxaq2HpBE+CwV0Tbu1tw3
xZPT/JQIoxoGzP9vZVkbgixOsG6B8yK54iQCFj1Hg9+9cHMiNzCdqii120ZuokC9EOvJrhQTIfhf
mPXTPmRlq+kcYS7tvek8aogCtOYygDjbLq3VvP9NE+zJ366uJW3UOskoiCiM7A00EwdcXakQdi+W
26GXSdkbwSPSRLWC1FXokTG1tmRSD9OnT6nz+r2e13YYgc8ArmKCQ5zojsn5E7zIIRKKYV/HoaCv
eoXtchbbFFsV5k/9M2vZGiyaQlzlxGgmv8DOMjinhGauUii//tx5v9F9QHqbDB2mSrUj217sQCY2
+5Nd6/JUxMim1ni7jXPL3a3jo8fLT2HsJU/69tL6d94PbBXzqu2IjLtWGcRpnsmAbYj6EXLWSRV3
9Bg/BIxZqx/65BahEy1WkixOZ/xwseOfvx1rxu6tgvVHYIbG9g8kncKxNPaKKC/RHF8n7n+2urCg
24x+dgCW17/WoXJMKHWbYjs8GIzW7KZS+Hw3QFRdA7bto9NgMAr0ji7toV+EeiZcbCxZOw+6BMGb
rtUg859lnmiYY1aQ6b3w1L0jF+lnWYnBoyyj+b9EPmbIwKMrj41JL26KGoQr4aY823pPlnh0HQuY
JmZpfQwGSR8Yrpw0aRGpLPHVGDs161nvMRf6tcygjEmwHZ9Gq4DEHGzcC56xY8LbAvxMZHp9Htp+
oZBC6pxi7slzZ989Uir3zZ3D0vh4GrbVqh9W5RRnVNY7qkEkgqY+N8s+J7oeQhTfwEPxeRsESjVx
6d5H8oUpmvQbKaUvayLoVlcfiIofPgwZ6C3PPGc+DkWh3BHmcz4ORA5MF1mGPC37uETnzmbzoObx
MCNry+saHHud3mmKCTErkbo6/u7+iPz8woGazos04sRUasJ76YgMH8/pGk69jlCEUmKfu6Brsn+a
KdXjuXRDh6LOXQuFD6cegpCd8/89soZStH9oD/FckO1BRem29gm3V+sa6qdVBbkxR8tGMjmE8oH9
xq0EVZKn/LfaKpkeO2r1VSJSubyJbkjmurKeHz06HV2u8LPadkYzh2ZEQKaL39+jqKoasE4s1cFK
W3KuGTiMVekjic3n4KbE3Zm/vElTfYxWwNsVkd1QnfTM17Wsb3NSDINNOJwgPLmgGZEGw02scui6
PtzXip1TlmxOeEbVkve19XmSo7FJccS/gS4c83yOtW+NniROf0tp8VLG4CmA+yYSNwNZy3fBVvsQ
aqfr3XnbmuXA7fy9cpJ1kaA6Z2wbBjSPCd/XQrlr2jlhST3TZzwQKfepwFbJKuo1WDXPZPAw1IE9
ptTtIPKybSr9fFfcMr3P7QZxoTyx9DvbwIWTK+HEjSNBJ+ZjPh/6zJJSUGH5c388Fp9LDEJOaC/r
/RJkg5IJOtZz2TmgbtFwlo8+EJWcBXWoCS4SnER7HM/hEEmZxlZiayuiek/NQnrPZ8my+sB/0nRO
Gt4MflNu74Pmo2x7AHXhnEnvPc4EHyHCxQwi/tsvxvRisi6mGEvZ8BQ0OhwbaoDJ/wMCTpz94yIG
nfdDAXRo/7A/0Adxk7t2dyWuhoCtRUbyLr8oAyksHngRTTxD+mC2otzG3B/lmX6Sg03g2Z/VydHi
WGytoePb5y5yqyb/CZSGvTHAJuOhGOyk5joDsWB5wHCAmsAT01e5BGBiGu0r0VbU1nQXvlfpcs6y
J9iUMp+0aPOtVxbVXpQ1miOH9+WEgUrr5MmurlolXk+qgxaqG1PQjfJJbo/eROYxfBe0gKZQcHap
lT8DTal67IRZCJsYfQMcO1DFp55l87KuCmtyUeuXoyw0CrfL4rkC8vzKETICPvCbZllQ8SrZ/Y77
+byH75iTvvIECN5SeZa0jUTeTaI7pQj36gW0kSnVyTrzM48cqQYgGftSgH7SO/xiRu1cwQbSoOn0
/MNUGObdv6ZTZkRdamoj/PRWa2Tk+eU5+sst0BoejhfdecT/axnnNC+ANS0Xd80SZTpKIrF9445+
VcF1gs/Awt2jwIU2sbCsXanFrilkoIkO/v1BIvUipZE06Da2RGzInKeKuKzXG191CPJzyDPTe6Q0
SfafzO/WaKxcdGtzF4I+v19aEPubra6aKrzk/ge6C9W5orWY72BS4bQ2NP9UsbtzXQ/Ti0kuea+v
eYPMtt0WW3NBAZ4z0XO9whZnACiXoZf+0Xnj7FdNu767YjjAuhrpAcKRiBmchI+zvrZlaVIL5I/U
WfIZbq8K2UfkBozFWiHzku63KNfwDrf+iwF0oHKHnIAayXQl994TdCUsRv5mKwiGoOgVjLhd+zjD
tNLriDSnGz3zcDz9Eo0xhBqQuQA2vtYNB5KzgEvGj+YG6cpS6/Rh4YnUjwgok/gGWDUocoNsaNIL
MNLgOsvk4eMcRemP+brE/ZuV5hqD6rpntBbvSmCrr2pUKs+PZs8BVw0F7w7t5hojBVr+YoFlv6gP
Txmm1tFsBdzNB4awWUD/oiMKLV7Mu687a9BuRW6HIbiLyDBLbkblJ0A+n2m0CNVrX1GeCLLaNsO1
QrpjH14DUmOcqWhmYKg+e3tP8wgcsWgsDy3g9HqezTFOu1LxuKPawxxctEiJm+S7mK/kMcTPgd5G
jb023A8mFTHqXRPIC03iG190+VmWm097rbv2o0NKL1Py/jS5WCKmYhumMB1XcGfY0bg/QC/eMLls
rV5LuB0rsjS7IOh/RTbtyImHUeQli+AKaG0cPkUFlrn4nFMhThQMxTfk/Sh3PH94uqLCyQmzLFNM
zk2we7Ql7ckl5aPtvr+9DQY8b3rCqPtn6fp30TY8Dkbrm6tfW4g3YxpkE8/kfD3sRPji3KwlvnjH
b3L9HIG6GOofnABnk4LWJxwfbPicZ7rngXbLM6lI7vEEF2AsSOlkUXgAgoN+xEhs9u/MRjELjY7S
DrfvXX3Rhgt42AukxKa7pNaQtN+2JSxurSmbpreXaNxnyck0IGy62Ppwh37XLqKKRYWjB2WaAd4W
4boUQyKRRM27P4+yzITKgBh7FXYDOsQ3YlIpb0ESSLUASRMDzuso5mWtbAEsIt3+UY29zIDsvbBl
UAJt8qrPlMG/ua6ECPE6WajuO2haYDe0SuKC4g1BQGwtCa3jdSyJuC/PKoFRKxfny9nX4gxuJWTs
JWytLn8fZWx7MF/DcCUcPmYV25krGZNVcP+lY+rRhG4XmKkrF3TaZpV8J0X2Bl46ZrI0C4tgyca5
/loVdYWwWmfO4iDasKCbRba83rDOZ5b3BBZ3ga5FdaJeULrl0gWRK/9HFHgHUYfZp4sHvCzAc67m
gGI7MPSpjvKnQ7UUHTUyGQx7JnirJbMArz8wgYOQmjN9bWAZdUtrN+XlAHc0FE12NfG6tz/ETk1i
jMYQXnM7m53LE9uCeERD1UA5VDJ0v96Ea2NbPXfJkGmxiOmF3SJM/mKVagcRmBsu4TndyBpa7CRy
SB2TKLazCoNwyTjWQYdb7HqFus173hRm2tUIuHacJZS2Hf+6y8B/cB63uTJXbXHK4KFRsV8GEDKj
Nc3LoJbt+HsxCD2nHfhPYerGp9m2Cf1onqaNGUKn0qVc+TbAbQ2FptewMkdO52tyjcXmbJJlMWCx
TAGyNaQVnLkQBVK8iTzJZnTvVB93+IG7NelV0SiweKKak0ySSjxQpsbjlqGlvzCCOtZWwG+Qcmsj
gx6Jgu8TSfCeIBxoI7nNuvqWlLEimG5l+zlsdrke1bb390w9hvebmgwfKQSXwnQqe5sP+e4PsS7M
k3yKBBKgmhvoOO+FhNFBcNHob7jTuM3iUY5Ps6A5gVuMsah73yPLXOBN7Z3cT7dPMskGL+IyQdEA
Lujfi1OMJrY3qeEnGIII322Jzn/TgEjMzD9vQQQaYGlN/gWXQcT/3JbnjXUR1KslGlccQosQ4t45
NxCiutNF0+bAugEcHyYmjLqukwHipa91KXay4CexBC6lhi1tRVCndSPYUB3G7FvNVdVEaBYYws5u
w5Skqj5Ak+AFTzsoUkYzfIormsu66o3UVgkb+j4mCq+TvsjwZWtTI6sO05a28BMol91pEJLhawnI
fHKOSQRfPLzOR8oaRqJeD6Xsbfp9yzJGssqiSn7oZvtZXBPi79969N+Rk+sdZF27Tu1IKusIVzDd
vc2miPzeQpmLLckN+irqY2dDR4qmbr8e4I2JRXreo/ZNNsMFWhWYnV83ySC5HfxiUL8UkIh6Skln
R1oyq7S66VZYp8cCskn+jJRqje1hxsMMv1lYRarb7++kVy6LwSkZo83Lsnh3UZqRerW3VdOH6KFx
RjaIoAqdiBpP2BE9m2AmzTFA79tODR/9fQY1xHjr6BdnpaPK4LcoBtOZdUi/vMn3b1uUBdsOm716
k17YYUUalYH7VWkeCKrDpffMvg+5SE/zGQQ1XCWkntdcHmU5GQDFck8TkMQk0qnUagvKC1jNeEvp
yfPx2xgBcFArpIPUWbuMPfdX8YEwtOytvKzwARbnhj6reu8SwNndI7kD1hyTILqqtT7mH8b6bkT9
QjV8emQcNXuwkhtqLN40pdi2iydYeyrXe4BlM1lnO6nydqHvEOvY0KgFTC2fp8ijiSVJB78GwpGx
bDxe8jiSpZJStrd1qgwY12XdpEO/d7oEobNV64aOe1OJ7E2J2hagOgkR+TZ8ap0ku508hF/YaqhN
1uiMOTClCvJ1PZYKPvBmS4TMspVZ5aV723oN+aFFxDfgqiNU7c9melooZY4/ExGNluA6krCcSjRg
O7+ZfogiDylkoYYUf9T+xR8bbeiAoMZQH+NqfpUIgFpLTflzfYREt2C8fbsev5E499H+qg3FLYEm
4N5KHtCg5/pzmKnXHwuaYY916D41K/kh7EUzC3RAqOqkn7lx5Yro/qBOm24ieHmV/ZQxfBr9D6SR
6mAW7CDwymURaF3hKL9Vk24m9cPwXg/JN2qJ5zfDGAA5+6T7zPJkPEKwYP3ea9aaQzX+5DPAVirp
oyKF1egAuvBSgWbXjqg41/dOx7AQ2jkXKIh0nXOlN+w/XW0ZpeOI0gFcIEN2mUR9cCkBM6HX1AxN
EmtUwHjJiLcIBlXYTxoTe2rIRtXPjTEqjiIgk0dd94dfIhTa8fJuwlnWEHL+/WtZbR2zmHrSexE/
MreNlLktvOcduEq/YCCr6SvP4mDBrVvEtP21XzD1IUr25ob4BZjUwZbe7j86i/P2gJFAy4hs5gFT
rU8u6LT7dMSxEdDUtTMuEamPYoxTI+tN1r+ER2uozLpnC34ssTHcJxu+V5G3O/y4EpUt8JzG9g8U
RSNs+RlA2ZT8OuLs7G0wga6zgnGLKOZ/qDKIV6/gIsumB0KY4MQmG+A4W92BaPiQkm1j/vOCCuD9
I5JbdyXjgzrBj9OcGB+cp9TCa66Mi8cRIfl3emHTlK9BifZS0BM9EyiZOQ5ZgAmprkdRlDcbEElm
R8xfvkZ4j6ugfa1OGZSei1RM0sBo4Vd229X/pNOfZkR65NseoSNzZfOYvxOl4206LwPqSc3IQICJ
eRT1eryGh31IFfyLFNP5qswlpNavkT7IgVB5QxnETIRvgbrJu/RkOXgrz53QQS2OPmIlxv7xVr47
WDXYrQxN3OycJU7ndncW61zsFZHu+x6HNu3kxDjnMqpxp5HR91x5dVzWcKiAQUZpsQPQuFZ02gMe
FbuqYx7YrcqfWhgyQAaFdTnnPsN+eYXAZnhc7sKce8o9TsxWQbOmxL4QbtOMhDUfIxa4klrAbf5N
/0pyQ8K/2zwUgqGq1YxFS+QO57PoO3UBZja2oo743pZrfv6Vx+RhKAmgUVyZIoDCTfdydvhkzk8V
bWP5M0pt1YN4ecvrocTI2z+RYhJVwcguqFlY9DQ/kcTSkinfvpdPcIkXstc+doAXGOZBE7tQ06bj
410zUFbVzYExPN1IwNjGFtd06l2sHulK0Il8MK+8JaqCRnzRNiFUVHn+cTDfuF0S859a9KLeycym
XLQO5EQB01SCPNpXDuTGZqvXePQJ9yBC00k8PXYtsjdgEQlqyWEPLG9+P/y0ZF0vezeO5ztOOUDh
m+/UbedM+/fecMrSxfjcf7/IKbdkcX0qKFf59jOdgDg8wZT3SFt8DGU+TBaBdkxZcB08dx6xa08N
JrMZCBCn2KPeAyqWjAjWfjzN8L1NE9YgrzLKEiY+YRBZSDm0j9InEpizqy33HblGNG7/PlgUK2RL
gcArl0htu8JH/8x594jYlXTyYbV13zibMUX5dIyYQj4ED+TcZMTAZVAIqUXUmjL1RfGLAfG6Q/l9
c8hzzHZOzTQmMMYmdAd986E+W34KHa9++MWQMw7SmZVDw+TEZjwpQoyGWORsYpU9oo0p2iZUEcZT
n7zZ/E1M5wS9kqpPWZ5mxOem6FwLsMR1jd2uX/ItULD0mVLlIV9zmGd7g+l+TbOaPS8CO2RKXEzh
tP/78DacObvL9XNbdyehQJageRk0TNtVcTbQXmlNpQLToLE+j/B43m5kqErfeElyOWWxX4A1DuQM
TpLW5HsTEDnwG/B8DxuGgj/PxCiTVkCPczabVkRVCdz5stqfFThC67GaLwGPukOidyYgtvi8+nTc
BrtxKNMIyDEY7Xk2SaLChmafwI7BuMbVqnKIde5Q2Apx6kD7N1yFCVSORm2dWOpBQLK49OnjErx5
Qs/bA+DP0o6SZL5A9WHb27ZFpzYSqJeoI5Ww66CX4wKXhXEZy/4RyPLZ8qnF5/MGtxZHaf/kEuRI
ouqem50hZhxVhahbJuQDBvMpWmXJcY0+HJrkLvcwHB5wfnEOYHAxZfYdje1F4xve9AyJf5eJ1D0y
m1aMmHSGpR7Ml9FkyR0hHEECPuw95j+Stmg9XKCI8o321O60Sy6/thPnlx1FNElpsOeACJFI8NtG
TyAZCtf/AEnWE+Jfkch481MTG09jjHUle1vBtRkIBZh6Ug0GXv2D2cbRI2mop7oQbNCGQDnx4FbB
4y/Gc8Gb+wIsTXwSQvru/k7lil1T40t58SQBk/AwtNF5ykuDfRSKBPnOwN5IwzzFQlKnh1XP8sKQ
1LpJuy+5uBMJlxX1ag9bATCMDPSjPzzOZP282gLBAVpSqZ7vcPikMDwYSDk2E6J3ks9Z+UMlnxzY
hUhtU4gHk1sOt1pS3K8HPnJ8FBDTPgiTmONlxvBh8S5+ay5F8uIcJE9F1LdSB7Q8f746qRIKolwd
n5tEiQfq3W4YiIfrbl4zIyTmOFFQxdT6clWml16uBR6v8fE9gKLzNDOXaZPpzx6A7PwjZFnmtSx+
TsTGV1G0/mynkG7IBSTWaGcuIBJV01/4wVE61VxhrBMNJE6ABnClATv0LuSfVDm3CKak5KPo+uyk
lEnXsf62vBlXjGxG/iQI/skQXVp0vj0xJKUKoIbobJnV1O/eyYphzGREzZClXc91NPnV/qoqYaU5
5DLXAS13BLAVnUlZFAuMmuVOyK09u3fTJYMzQW06vF7M/Of/d4obIINhYhvuoVJacEDbskN+g1Ex
m+nh2FawzmVdvLt0Tt3UC0pxFWqxClAurQsRbiyJWJ6rUMGXgb1m1uODPpXWmk+ttDDxzcO5py37
QDFd6YXMCfM65X6sDBwDGbNZh+7es6B3YFr4jN5KpL9/xZaXOtGWVEu2pzk5qTO9leirjLKJG/Ws
KFy9C7YG0tN//lwUt4CF2MQGt4TKYSw9YfTGquNCHB29S9F5fn0ccgGGM8h8XYSxy1rkXEKaqpdq
H23qlgrds7/kG6ejn/c/SNGINd7GsZrKhiIe12Hh7suZz66WRhkE5XVLnQsyonexgz/is65EW6rz
4n6BZ5mKPwFLB9ovLgATQFRfen1gzmuKirYyA05MhleE0MqO1qU/k+KJaTibxCscXXnKaTV68wR2
JeJ94Ma0TBPbC4eaBXm5von1hCPQ9BHnP8VT3eYDcP9jkekJn+hPY0eIP0Uv7SWBRr9ltQJmUCTn
FCoc6kIojrrklv4AE8sVmt1Ts0YYtqo2L2BAv3busCTGiwr2P1bKCpPQxZIRlMObPhxcIfpbiPCc
lP9L+t3icJiUi3DQGSiFSnwkLbevSMV4u1dyiJiIGrSlpPYksu5mKSwNZeLs51Yx5D64wgHccrN3
vqQyIqjdJC2A3KXTPfdBTcviSEBZwZZs+D5MV/dfProuA1fDbVQfRa5tDheQ5fDds0HS8Xkpn5lT
YONJ0UfkvuAtsi/7jzmnDNSCghf1NyFzxTvMIA2iZMs2GNcNf5IJW0UxXCd8Pm9oFXB26AF7yoQk
G2TpYmPzudv06VXrXqA6zJjyQi7yg+sxw7JcFvl9DRSRngfjdFlNN9qrFE9PmR11yjFH7sF5n8Ru
WMffOw4AhUHvapn+osy2LWhLVArCs9mVnM61dsLiizofhpVjaTf+EC2FRyc6lQ3qwaQzaCh55BC7
MXLeQbQX5LfmUBja9UopVN1DX+ETXgXnCWxUMXLDlUWVkUq/mbD+eTKe/0ewmSDXHyXy9rO6SbSR
nmkcwth35vTg7EcwuNjWb5HGFJ9yE+5/HD/or4RJv8jv+9G5yyufte4n15x0K9SL5OUlCpslCeQR
sBdyOqS7RW0ws8zKYScrjuqmXVZCK/ujZZtk+TUDBk1dnrJoR5fcGEcDF3msA1pwf/5XfKSrJsRE
meDa/14y9v67pzChQqmDC0GuqI21La49gPh6YR0+YTTD3Fpz5XSwBZIgcMonS/VXKD3ue4Hp0cTO
qM9GiAVlO5JuRev+z+il0ff/wHx0kNj6XQCjLOW6bTM2xcPfQv3Ded1TlpBdlSc+nxGXlwx8JqLB
NK1Y5cuRch2eW6ydysttqsbtrekTpv2OI1jqWKHN60dY8O/4wMbawI9jYo6jSdfztg9HU70QRJgu
epChgzOCZJdWg+4mesc7MrsRfXHIObFPYP6NZ9ftsReSy3iaFyXXwP2S7Y933pj5/CM8sk3Xc3EM
vV9iHsXeiqMPMekzetUsFtXwTVimvV/nLQAmmfaug+KzG6Be9VkOeboP00/YKBBycEjsrCETZgYk
niS9OrxNDB1hFLxoF7irJ3MEaxjs3kkpHJSKU5VEA2xSY0a1fXjp9D6rhs8iL6rlPftMzZZuFBtI
JtG/Ov/GyR6BqYj9BYWrv8/2EE2GiaFbIAeMi1nUxGiOcHj3mvvGBtmWMgUchO6vu87v3BtMvxsL
/T0jOGqY/fISWIObtEKGgAE3AvjG3hSom2/9khb1VsO1h0FGrSMZc2FaiQDtXDnwaoiFGb+8vCeU
R8k7RQ16cboeQbPLqceQ5evrHBbDpGUC0XwoSXbF0GTBtwSe+PKDx0JXz0M896ORljp8Z7zYEPQJ
NyAUcs4gwlwZK+TxSVeLnUWlYiCWQ7wLtmH1wyySnpOlX/hZ7puxRn1fkzdnx7gDg0yJ3jjTxgS2
9sp43N2IjpPV1rn3RNbvPbNZzWEgoTXTGplKTHoEzdDPlcsX3hHVtQCJue/ip4eaojLc4ufomx0U
x9NGXT5DypUd4Ei66h0J518E8JlRsTe+DchglMKpQEFSPvL13PQl6JJQh8PcfMUAG7epJSoUekgs
gFLD7ZkhFQi38rF3CE08g25RFn6a2K/BV2fo6Ns6QQuA8R7TOiaD1yKu2G2+AbeWaXy6IZWFlbPN
HV0tls/cqAAX0uVlwctvYbr02UjJ+vNbOQOnCJ1fHna4HYMPFECdxch55WfXC9bGYBPVfxTAd/Rt
yPsC7kJSV0Sywx6rnc76MkrEpru+ieBprVL7SvpTOdKZjqz2/3EqwKfqhmDWtZIzBBQ24dxi3cGR
Of9B7jCZjdjyzppKp1RRXTU7qBvKl2xXTtc2FFQHpw6Jtdby1bRwLgebrILcJO/Darp+fbEGtREp
YMAJT1qgPVX8CvypaLmiXvDa66cq7nbX83YSUc0TleKPDOGwxKYwOCh4vXpkiEquAhkDikPNWFqf
rGlU6U9N86yfkrPY4d6iXrwp7P+DlseScwewP8K+GdDFm8nx1nRsVhatoZ+NPFnS3gGfAMVHB2X3
IIURsFjU2BEpcjCK3rszJigdMO7e92d5MmqbIjI/K1Zlqo8/qQG18Jx0QI03J0MBctE6Fc8YNVty
wQ4CMEpWolGr2HraPT5tWegLV2e7xvH/1lH8UHZ9jM1/J/fzEs0CCgWYDjYCe5npHnbV3l9+jiAH
8Le4vpOFaCVZjpECIQioqyIIcsEFinxTq8yYHtOOCIUx7s1faXHAzOCCDXy0/bNu3SRtqgvz8jrY
3BNGkQ2FI7WdbiHoLPy6jbnfetqDDj5wMNDhBzYGIK0p1yvf/5LRwiqO3Wtdnvm5PCmeDn8x2re3
1rr5oFfB+i7aG+/belvcrQn2n86LoUPjv990YhG/pJdccj7MkVOuyGQlwU6R+LyYHWCj4OpMG7ar
ZjGqkT9GF8VW1iffjemNeNROceUlyQikiPjb7AQ+uIe7mmMt1WynPp8BkxS0iu1J7Mlhao0Q/1kO
IZjOec633MlfnyhhzvZ8QKS8rg+jQEbNJ3e/33CXdvdGoDWtpQaEWksV70tFUVMTWb/dO7aVb8cf
e299HYCl9imysLuHjR2YOWIqrHo/7GmtsJGCIQZl0lTkfKPIl4jKhjlbkfDoRwfh4aItj7j3BVRX
FMfpBq3sCP+c3l0Rc5Oq6WTQEl2pOr6fjXjZYJUD3LdWgg2s1REjc8SFbAbzajdpXhP0Cp1WSqxd
Q8xUHXeLn7TKYD0G9S/Zp7H6sFa8tKtF0rVuKx2b6vnUYIt1r/JNUSVacRg5/akRQVjmKD91Nr0w
/8u+pKlp7/0Bec3B5HjDaFUjBrkDA39zZKIPIcw6li4CHRkFgwzdunOS4Sx7+qoY73xN4X8HtfDH
siSjt92jwG8K45VdprMr8KlDCd5v5Vl/60l1YQuaunh3nNmNnQOUvnkbRC+Mx1HSp+WdPcMGJIYv
25RTPAqcCoJONET8Xwlnhbz122y8H33MGM2XiYZTrH1EEDdirDH6rUzblpeDaCT2UDg0DkXQkHqT
/26zQyMkfr4RrectnnOWqWwFpLYPtjzXGjEc3CgaBJ/SFtz+A071jWw2DVhTZMbtl3z2cvJGVNB5
EAMQ161aqW3ES/IyREaULNEWgVuxnGu2VnRjAgscDqeiBiAOIcbyw6KfGAsYY8QkcAdG1LSl26GV
bl8c+TdJU+pk1Y16tgByi8/Yr3M/MBXt/FSi7q+dpnG4P4SaXrxbwZAKb7KJBO7d3nhjKNNXxj17
LHjQ8yJt6sGXRcvWVvYNdmsKS6T8Ardfnog0d6s+DS8I6xFQqEr27WXJkAKFF9QpSmBjhzOltqI9
oZefzNsVusA3TDPnkLsGgs+eLZToC6GOAx1r4XbXB452kB3nUaaaxozl+ssA+x4fS5ETS+3P+xNZ
ds4cWCVQPUzbpgLfqZQuC9tpintOBM9cYSJTE7ZUqegZddJg8hx4w62y1oVz4eVAImR8HYr4A/hj
jOaz90qsQNA2iPq79ZK0mTrzuvBKLuvZR695OjT8CvTZZYpznBFLODQGMuX57C5Wg5Q0bYhZsDSS
CZZnUfNVqk7F4lKyyMoa0FXintl8VVzVp+BWSEGqsdxamGi0lGascuTcX926jKtRJjy8Btn+YAVb
qzXn/aqVaNbc2lAsvnYRtHOekhGpWyLO7G2z7XLQQ3ne7v9DMUJX3ovSEh8tf/0JwLi6Vk17mOkk
jpOubrTsey97Ei9U5scHo+Wdt7tdtE4aL2Fc0JSgTzThZdU7taMZNToVNGyIX7+VKKjou0ll8o8Y
GPdkfrcHwzImxSpzasyxx910IpvUtxsO834NaA26VnEdoUitAj6l4/maGUaqMmnD/zgS7QZ8ra0u
f6tgIHETT9DXCrVf7if/W/sUXV70mGpSoBch9fCuW1O8tyf/j5jD8SO3a/hd8WK+8sRyLUusMMoo
f+GyLoG7zds/XgSOoa4QUBtuwVEZfCjIbkHfAKybntS28Y2cADpeUPxnofBkQFYitnJYgmVQFf6c
uyYhi4WbJbK+SO6x9wIIUkdB3b2VX/JzDvkcPCfYELzgXG8Kk/+AHcijTi0iNEyFYPOCkX875iO4
pxVaWw741FbX1PVqOXFdQcOWImunHnTPGjHS8zD8eEamFb2Vlkph3AQcQ5lMbvgNKe1AKdgnO3sS
FN6gbR6Tti19sRxZfLGm/1UA3mW9jNLkr1sRXhM/f01EBnsfwUW+Lj8yMCEu8c8cVUExzOsfi7xx
/BUJ+T9zHvPs0rcyZXi2qsp821FAJ/zxdl0sFrFihRxHtR/f92rNExbjtzPnj6684Cjz1zhzrRXs
7XvLl/40CodZnqcFClMzc9tsVhe1R3zlRKnl2/2GuN3pfKNvv4cu+xpLaig7lmIxs1r176QGw0vY
ToPSFG/PXEzlpe5wwC0gGZRW+pKrQZiPF9J1xya8QbOk2s07CgV+0WB4BSDUnk2TxTPQSrGVNcnM
Aw6PQqhgV9Tzo1Vi2uRoHAR1lpJ2QQzmq8lCkY9LBSj9oGhOPHXhiZE2g3HZkbIiFU4PXa2N55dZ
JlMC/kDNqaFlwC/TYPcEp4huySqLq+dD8KdDj5DW+puAeNhDRMB5LrayPNmRCT6HlKTR4hn4KIke
W8wQicKSwjzRXOtto4KOpLLP9r+IgNZ0Sa/+b0jxyhTQFApBwhvb2YzcVOnKA7zCQkAaRk+z+7E6
BOccSKy64hDJ4utkCrvmu5MLLQqf4jxKjb4vwSt6HkkK+5teok9SM7xWdKfstPy3YnF6ZiZ5oZGs
pPmg/a5koN0DfAf2wLjc6zhHhY72r+ha8QCwuRL5pYfxEYqUlriULiYaVKESYntpa3sBmXYtBfhz
E5WchX8Lsk279ST6raI+3lZ3Sb+QudfB3fH0ooUsjUVAl/FAFIA/Y4G6W2du3Q4wPEFu6/1V1WPD
zYUMgJHKLgq/buMbH3vWzEH7WRp+WCqRYzH8g22sQCnM0rsADrm9qyDLJNa8Xoyt47l7t8sNHYS2
ltEyut4rYueVfFi7CfbyoDPAjZ21gkaFjpdJanlN/RXQqCEMXQz+mcGHrD5NQkEMYc0ua2dszRj3
NJfFtOMeIkbaNhXPz478VbhtM5Nmjbz6+IO95NnPOUq1+/8UW72ZSuM+qqA1W6WkO+cyXTcy2PzK
EFGqeJPO9IFjUW52xW66mrYUEgtHX5DgoIIJLa9if2apLfw9aNnA//H0JMvq9tcL6tVXsJf5KsEx
Xjz+3nbF2Vb2afUZkve+/gVSlpmIzQ+LntYyzsoLcwqTw/LagBBYMikUd4jNscmH1waSOBTgZrkY
lAB1GaqVW3eF/v4yItfB40zeWO7iuSVOHBg9MOcYSXiDRrUjb8r0M/ECuWK14sKAl7FJSSjFCxyK
LJFhJ6CRThZqNRoAZVFdB+6FEgYONMCxYfSgAQFSQUG2Ig0pkMoepF/zHs86M87DzyvKeqezL21H
ODU6RmrLPduuzwr10iaywQW3jkZGJDLQyWEbwNlEwzKFqJogPcJTluZeHoWMnl15iUWBsUOsn45A
+45zmRdE6wcFfW9p3oYcz8l2ZFlt3mHrpY2XKfW7gPbkFX08pSWnJxRJWa8FDotxdd34hbC6vBQV
3kNDyVttdYuc66e/2OEBwoNQ+LWrcCNl4S4sARcM/S8qA1i7qub5G42XFfV2shw5BObj2nEcK4n5
SpkZsAa+WNaEVMPzdOtUzegbyTG5NjjoDWGsNUN3E2FSlVqEzqyP8hw+FrLft4es4lw0s5b+5N2A
rfgrgPDPn6r8zibj0YaA7hmEujn0Kku+jckiD1fer2Y1r5nwT0Pvenv9ZDZ9etKnSM/8UwfoAefk
Q1Kd900b4T1+oeOjNLqXiCIU0ZsLL2KxMiKYGSto3yqdo9O/evpBev7qBmXWbGclYe7GXGreihYX
h3YhDcijjyWJ7z7IV0jST/VGE2qYN9STs5TmP0oNO2VbRcrZ++0MQ15OWwWf8yC11gcAfgmaaK5K
kk+rnTUlhH0M8tKpZXVj4bjctS8IAp/0vktRWy7Nzf7URGA15voQ8d2m7WpkEEEjPyFGiNJc3XHQ
gzl73OfQDn/sD8mSH2mKPKdAYmNqcQ/3haOSPPr5lgK165/K95LJYsSK90jWsQ50YgFFtj5/zuSN
/ObBni5uUCkkRZ5DB1RAXsgXsZCQ6Y+henQ2Blec3WWpF7aQVd2i0i4b5YwAfDVn5JZdawqXe3cJ
5DOd3z1Unw5LP/9EoQf+etOIvNdMlnt1KpXXIyHkfwHWN5gwPjddp5V86pr2kwNPYwaAvR2O01Qs
bS/NdFZoIMqgrRI25VFp0aLRoaNS7e+ifjhov2gQ8J9ebz3gs0yDRVZxET8tfbSnIwOU1giFhzhG
6DL0Ojbk06IkxUNgcLxJ37oqwQol/+YTxR4jFnJaUzQB+TP88Ppcdrv4XrGrMyT7nBJ8rB2SOcAg
OdvT8FbTnD+Red7mxK5ilt0Riq/DBv2jdBiFCK5L3mHoJKtdDL9XG1Srv+l7n3EAPHuTZCUruVJS
B3gKlYhbkY+qSw0QdpZB6ComXiRmpx12zEzRT7STBbr+wIkZKdXTzFe3lDwj/gqXbvX1V8bAjtcv
W/xPbbHNBMQFDa82int24I3kqidzrZt8349wxx/3d+kD6gVdZ8sPMBpQJ1WP7iBXQskFS0IfoQYN
Wyf+5S7cnTVEMjlHjMtegJoGMpr2hGczoNBRteEK9i/GszhYml9hrmEPa7Skh7eQK98MMgCaLiSa
i/c7Rt8or4MKdVBnvAFngdT2qvN8RkKyNa8t0EKK8X6xVJ7xlrTlz9ILlSqWL/c8FZ8ABoXdVYyw
XNx2upt1XhZ8dpEGjNuij0tFZT2we7XZh/FZLcVLgZrBcEi2k45VLQz79ZFcimE67+P144Z/DOA7
ZAYT5YuuaH/t2UzSj1RbKhK8sP+++pEd54iHj6Q/1Qf0O7lk6huLA8rbO78vWxOXwlt3szmHlyZT
/8gnM+F70tRcBzWNeUa9N06j55mBfpow4Blv/Jm0i6iMiXNNIlYIKqTJdCHIQgU3Ix3BIut86raD
2/HxshodX2MPQ+ZirZ+8kn/mUABs+YJradvjGpZAeBqvvp2EkpPnTB1UliC6gXhfj8xAShsyeYqz
9FFzalbCi3gSFoY+1NrakyMjgAqqgIKd09PtKuOXQ7kFQQwyOuhiaSFt+em20kiccRXNQh8MPqVL
eky6RkPRI71lbx8O7Gtqps+MnFHGC+YbqoezOkSwVWQ94fe6Y9nzwV/IKhtzjfWFj/ZFCNqdpbQD
4abVgOK9EQBLJ2VomgXvUX/UEoJUkavCAv/9Q+8qD3IEit8SBlsktWYB0A47yRCrpGj1NGzmb1Yn
xiYYBpvnjTt8+fjk9zUu8Q6tQoFKpwSvvJSikMPiG+aFAPkmPNh33zxaKJWCKuAaj2QkZsrcvq3p
3/B2tnPOcUhtVrSp115N7eybshUeNCM+BrO4d5xi1zyF3BtnGuMFo46OVYrawDNX5QB/VswKjNQM
mZcwWN1SwwcmkXSNzI+5r8K+JQ4PRuRmfK7mdKgmNIdY1oXX9763t+6wnhEYwr3IP0fJx66u/tkG
6DR2P03sOCcUYQVNr8QCwCB1kisUUcZB33hdkOHS4fYfykZE29pXj33GakmZZnkXKHdaeJG8jbO7
6Q4X/hwsTx3kenFHs912SXD1cqhaA0tewmG76phTpkMsdn31In3M/MD3uU1vT52RU0qBCHi2fRhL
Q+TrIf2h9TlSDzbFNs26f7T2HLGtfHXUZgTi4XnwN79MG3LpzY0sECebI0Q83vhXvUCr6UW5tpEJ
BLHxvgppMFLe+bKEOn/SXtI6yo0t/95rZ6UYsIUXQ7G0tsQzBG7u0Y3HyBAZZNAmoNU+oAO+W6s2
Gs2IMnX7sXtCeEH2jzfwLt/rLS2MZRQcEzO78RRdVhioUabIEOuoo/39Ji03nmpSO67XJxDfXhaL
duwBaNqSvvrPxCCugpXTUMSBlbzNApYCj2njoNlYSije/xZo/Am3OFs+7nr+3CFlD82Et1ZfMRGj
R/oEnPtib/YYjo9qubNWJTXZC1mmlMM/CyIomhGDqxJiu/6An5UrSC9LFB8+VYqakY6R0zYOlqv7
wnWPjLNdqS4FR2D+G/Nt4EN4ExKq5Zq5ixrMZjbHMktzi8feVjRaZiRcB3AtfkSEfAOusR+ScgkF
ZGk+CFhboM7X3TpRAvF9nOrR9YIJji9BBB57ci7p/xa/0zBa3kRbnn4wiMH1WUkstgjBKSzGYJxv
WrNcb/vPWW9vlUxvoVEly+9pGpMJ/8N06OmCdWTzGzmbdjWtBQ9PIDM91LMFEL54W5hGbbFeQxWb
Z+xeL2ITv0SHZixLDQsTKQPY6F8Dn3Owic2SLjhwRN9qDJzpikz8lggcbFem6m13OKVphtrvSuvv
kWpzrOEBbBfWbh6pBXgTTbp7ULHim3YTRHE0TXqgzYnUZICnGKvDjwgxF0tplo6eLuuwR8+KjbrA
jCKwH8FuWDFa+fp+GxRpj+bd/ixxZgRlCQHz+a3foitUP8CiVymDVIkiMi2o9pRc5aoCAI7AsF2M
Ln9lTx8UnFDWVXM4D/UZdma5LvHKS/XQwY5ty6ygwI8NG/pLJwyRRpgVnsAwvpTMZq3gCz0MEEVy
nY8nTCvFcyCoXAo66r22Tgj3na5I3hkOWFLAfilHWQ9PTWRi99jUyJqirjdF30I3qDG+p7rSWnK1
0lsBpJAzU4eWmA5ipj5Xek5UEkOCbsJQVmPLnOIYi94VPdJv+1kksRJAtSF6XqFdOTFAeucHdMdo
24/IaphVDiorR0BK7Zc5Luds6tR0+xHSiA+KvpI8ZonrG0p+TkiuwaThrGQqSz5iCFCEO4lSZINH
tez2xRblIyvjHeat7XhfGitQOp+STeutSnUBjtInDEH2vJhvvtOkgzF+J7FW2pYQsXUCy7DXKZTO
NEhD45dQead/fF4flGfX0qAEkORNzmgjR6ZKZ1Mc2D9V6+DjtlKB4niRcFG9PYjMaggTVQ+tztrU
ZZxEcD/acV+08SFaC7Ja4M+VfNbjm5XD+8Ip4dxBUIDz42MZI2+4jW6thoi/WTlIXrKY/8LMWivE
Dnp7waAHmpu8K4sdKyf6fkBF0d/fN4eLEVICgVXFEx0P1nChNPaVecInafigdJUwvulf/zp6CdC9
mgvzyLNq91OoOc5YOMGTJaGEl/r9nfYcZCedPCWI8P1aXdiX1AwuQCDsHeH+yzHw2sEdiJ7hSLG7
su1uqYJvvv217bVQeOoItq0fDa3spD2MDhR4KOj78WwFXiUi1rdTfxgEXJmzfwSwv5uyd0Pnx4U6
14DhBL2TiAprLJY/x85uFbc6nT+Q5sFg0do7UMkkw/t0080bBWUSAxB1HnODyX/R3+IZAcnUE4xx
cHDRp4j4Jv3ZzoaL0i7ztdNXoXqX3DDdoXEdJ195WAxNOnRaFWDDYFE0eqZnBK2pefe+QWMeHq/7
GkLRDA1MvBTR+hjc9kfwrJRvTDTqZfYxbTJI7hGto0jBT04tsAEtoFtx0VfSo0LIL09FDdLjkuBI
I+BuKv8x6WLgBPHaBXLfIVHL8ODI5mi2RGXumqKdtyV4dsIWat34OkQ0Wn7wnpGgGPewbwiT8SFw
bTIV9O5tiJZZeLiOU193/SBt+p6DwqvrEMcixC4uBgqNdAUt+Ai3UXcdoFqGPa+hRbFiJ4bpYK+J
v0I/St3oOENvw5AhQMwmYpXQyuBGH2Ig48AZJhYxL9Y9gUDkO+EK+NxNthioU8soKIq0AUUVXfPt
0TLRKVM7Dg5OomD1eUdcpwI8cx7zcierDcuALr6uZ0irWhmm1gO+uwODJsiQ+A7udl+LZhH6oEwb
v87sn4plU9OgPGKQ8w8Idj3lFR9b27pYAHARNEV78USRqUnwKzRYrwplNBvsrfKRqyGpuqn99SgA
cJkh4XzNXvH+cZhkPNw3+TAMNc4v/wedsqtQQpCJJJRTw8M8RbiXoDdY/C6YETYwyh19TeTd6hTa
XpGM0ws5JcneG+l/2uoxY64IGaXGuwcZxJAtCJ7d2Ynh2cRLDkXayHKDeTO1szPqn1FUw1oAFYsI
/lWsQtSw8ua5ZoCwpnsXemFCfdKvO5gb1T/G/KTCDzymRtauUkNhn4gdOhaPcgd5jhT8Jz8xVeBw
miX0gqjAOokzLrZ546YzZbaCJtA2ld8S5XG+P8Y81PE4E0FN+zvmoceflkebbouIFzgjLcco4qDX
+PCCPRvPZHUsiF4FqI70qW/QhLVsHLixiZPDlPZSVYRvMkDu89D99NM35n1jUlGi5Zv6XNHVKizy
9GYjCeWnMy3Zz+icnW2engdlsX/nnTt7LZfy+QAmbiqU6CumXq0tDhcBhPctyJSCTHtjJmMsrlUK
wJ5n/jtMkoenfSEc7QqzhGi8mDiTUpQXZZN/gOrR75HtnKo8bpsGMcnzXUWQV0Z8oB1BRs+80v32
s/5ymA/Wb565PtbCbJdbsnuX0TfHYerjy+d9vE3Klt0GixdsE/ciw3dO3zEMaC/5so5OVlaHt0aQ
JTT/YtVjOOb6Im0Lnn7+H60SRsaTculkHOLkPNyyD1QaAdtuNwbyBxaAzwIDqaHeSYY9/O+CF+f5
RcY98lyMbTRUvozaIGTctc5TDfz3IEy91iGI7ITbDigOBCdGKNsdWHbU0fWqkk66kQ1aefFaqzu5
sjRqR2cCRwMYnHPtX4nsgZEFU3G2V21G8KsdcmcjKpY6rwvpyXoXUgTXG0WaripDOiwTmulYVZcp
P3I8BGEjmElB40eMpRFFn2lSKKJhd9rhVYjvTbi7WeHPm7OKU+Z+TS7AqBGGCSvpWbJLPNqoznHE
BJMBsWV1P/Lc4LEitbNQyU2Xmem9u1/YPidReTEGCkliySagEvZpjF+3Tnk7rRnkcN9WKWIBtp4g
pwL1N22kiki327/zodLuJSdRynTu5kbYkm1GNjD0WyZCbezrzEitKD9p6dqT9tm6+hlmdTSSStRK
YNieTqHQmAGANDBb39bg2bSHfS9JC+2Rqn3CXCwqaPHRwv0VMJXFnO8qJbX90P+lQneviqexRdQA
Xk4TDD3dmX16lz5mFwncZ3Ix6BJo0vqOeCizb2PI7kp1NTsWCerVzV9zXXYBeaHvPuYXEM90YrOw
H7YBHej1YGuG+PBc8EiVj/tPAIC0XS8ADVODD1OiVVFFz7IGO1guPFj8TQhX3Utz5h7niL28I7Z7
MU4NzeNWeOyBOMRjTWTU0KOPSYx7vHV/hfbIURn/O4fW0YFzxvJUoG2oo6sd+9VKqzCevnDuCIgs
svsD6yIqE/jfTa0ih8Y+JIlOF/tHx1hCN/zu6y9XIUr+cPiAGLOyb7ABT1CpWhRGNhK1wRPZfNIw
Myhng4Z7lNqgGEBRKHYkwtqv+5ugctCtZIT7YNUnZVC0Dnswqpwii7HSYpHWu6jJ1yQKdqCOwwwt
I6pTgMZTC0q5mk9L5C2bzVUfOSxT3UIYkDWjnvoOvDclNNTXxG93GTdJ+/l/XzpXW4hK0/F5CvCw
TyUc8JliujjO2zmUxBhTGPbE33ZNcN4SILUfY+b7eH3D8bdmdGauxnFTnUcaGl9eEnbz7Jd7U8Di
DZfoWsBeitUdavwoPLBZJObThjRG4y1MP/zH6gd8IunCR1T8Jl9p1nHX0ujU/y4+O0uIWjZSztIY
2HOjtrMO9IZO7g88TL/ybhxpjNlJyhpNjb0xG/NTytCfj/PONTl+q0thVpjZ70iwRmZfvem19Jqs
YpEEbRFXSo9FrMxZHzZ8vUQsHsakhseAiezfXFFEKd0eXQ0R0E8efWYZ9pVM/TNeZL2YdRzChOR0
PE+sj3J8a0AXpfhrcTrcaj1lJuiiu/pEPBFG3cIfp43ryZhOakNYnqCS3U1z3O+NJ96s51vj5noL
iI2fyCKO8Z7fvZiBgrfDVfPVL9wkSSq+WJQPZMFXafXj3Q+iEb/PXZPn8HCFJCzXkt2CPw9aMCAf
iLUo5tsvE67HgRMbjjAKkGrFRynHVNd9x0EtZbCTPbr9VBGrzPZM9CTnvnwBaRDcxK0Cmmx7ZkPp
plelX+JZhB7j8cuaM1YNTteO15169736cnZ+eWNRuD3cA+S9AAPlSqK1xNnzOF0oJNNgPSFgbp/D
vh43DhcICuebQ5lCrE021OjUogVqNzzvZ3eVR95JMK48Mpggr/fKAbRLrwFmU8tZFxtoFLNjU0ar
bQHF2gmSM+3RQhKKdb4C9LwVE2uTUckZogncOjnqSYYVzb6gNCChbYiWa5MLtTNu4JrKqsIG5PVE
5qR3XY2dX/nw+G1kBZzkCgSOzp2S+oA+CWlOSLssqEmdf6NARnndMSMmA8Co7uvYmPRYens3Fr49
8JFD/pr+8eb3qB+BBNovaioRA8Asu7HxVEsg3GwYPOynR+PE6RU9/6XamqFGTo3t+DxSKzwA+aiO
30qVLdI+NfCJ27FHGA4TBiAox2gBilrtvFzTKmkwv7uJIM/VAstA69j7QBFsY8Ko/JNSKSeiYDzy
HXKpvuNeakqzv8wFlhq5efUsspGN3ky1jy1PUw+KTjDarmh8u0qcCVwT0YyzOhFfDz04s3U0Or7Y
ciTp1hFoNZZRRwmsAvssrt8v6ZE0JQWu1qT8CpRKT5KUllCOB/hoBKkOTVS1VDOQj73gPtgf4VE3
KyTH8vsRV7OQI+jsHUp5B3LSB9skHHnZdIa3nIsKNtAzQTtkedtL1WmvxaHH/cDW4N5fh9atsiqO
Gq9x4TBDcLh4382JHGY7p2abKBvE3sW2AMQVDj10gv3JpRl5M64Y9Ev2I89ensWr2fQi4jrBH8Qa
L+2VADoFIqQ+M8f2JGQXeYrSHuCo2g9PSrt69x/cjGRC2mi+OE1vmW1/qnDW63GNvMloQvSAuk0k
o63VoJr80YH5GKwQyYW5ACRf+z+BoC3Rv5k+udxkXgqnnRWQ2aLlJPWJ5x11RugqmCwPaiUjP4e0
MN1ifUwLUxCmlzANzgo+91nzmz1RPNpVe/XuB+CViyPCYHmjIJbzYaMup5Uydb9TALVGyiq6ssUK
lrJZC1gWMY73bdQd/t/a1c0BEmfT7aiVnpViq+7Yb/ZxEQHl0llr0DPLJCj1Syk6YISIHfIb+2ks
Gn/0KN/H/i7a0n4D9SFYNPO2PG3ryVmzaqARK8po/4fzhMMRlHg1ZSPOry8gXAbsq+ONozoGNbj2
OaFIKb64nfn3307TF6rztaL6Q1WFDKOHVn1niF3mU9lpLC9lsKuJ205XXppov1MgK9upwggIJlkq
DYsTYV8hBt9Tli++oBoATEpbvvpnElO4G00Ys37sUSgZaZz4r2SGjLBAjOiEO4tj4GUGzt3XGRp5
ddybihUPvng7bncMu4Z8oxxHFT1FEcrlIi6JDl3m4rvB9VVmZHI+V/pK8xMBHNn76Qb84IIMYQW3
AjxShHYl2BkQ0i99O6fT+HcWy6fQGR3AxAn1/0D3jd6TBWpX8/GU3PzIbDhBmA5HuCg+VOvU2Src
Rsf9kFnQaKTK3p8IlWyFz6A4G8c8TxJSNJZ0UV7ptDYnThRTv1IcPdq5XX++WipRPVTTjj8dm7nB
36xzUwGdE+ZiDpU+/x2DCcDQDc4n7ZlebcCVQHptRzqCc52QXHE7gth5foiGUD8nDIaFy+0kZpX0
euZqGxGAcrnPQ1dxPzfSlK+QUcvgU+EVkRfUkbFs1ENL4uMdwc0DCBOvlp+RW+PsSeAHyIChR+rE
1geJQi7FMhZASCjPhxsT7m+G+LCe2fZsT7WO0VpcydagqS5IjBPySIb+AJt1XMUWukzbYgL85PJs
BSdr8yzLx2GSP22VDY31UrFfhI0KPHaWDghIWj4AoQCSMKNMC+0k9VBIVc1B1E3chuLbwDQz6k7P
868PLtWXeNU7/ieXyv6LFJch1ga2FseNXWu5RSXHDbkZvLs5VwrUxkVYqUCHeCV2qUujeMHq6MbP
dJsu9r2zrvwwnKCt3VHa5fzfOs3B51PW6aBSJ2q48/Ry4ZfxUSK9FpPr7IIqi1kprPa91H66l0uI
UgMZdTZ6X9iIuE+tc9uKoK9wi8R2Temis2xkSs541z/8+PgsxmBmnTcWk6GoJeY5/1ri4BbM1Gjr
xcv/Fxjj8d0kSMdpkqgpLGmmCOnyveDahLNIgkhab6DQFqj7HlEskw8u1+oZgxRPC2ICF90pMYiD
Fe8u2i6pjX1NdfSjQjJnpnZUrmF4v09IlaYG4/filmPz8x7GAsSbUxYmlQ0qrCItJeIL+fTcXb6I
pY+rfILi2M0sJrZSvfefphEi7hZcuYosCqFF/+RkOQ1tGNohSWURNen7ukuJrFqbiJPxBkEhbjQT
rhNoGgi3jQaJnEFIn+8NWJEOIiUXXwRI36YG9GIGhzggth9CcN8hHSU4NQ1chL2KAHqY9jAuq8Eb
44DMYXQUGeHdPFE3v6T2yiRd/qxcWQCb8DCj00I+rYScoxfvvQ+yRUZ67X6LlgTevXF/ZHgIH9Ko
D1apdK9AHcQou6EJ3pgeB3e++lFM3JfKYi4qyT8zdCZgtjKD1rfadjy/i4Y+JgavrRddab/sVE5z
d/LFFyXRnkFxKrXqcL1o9ZLlDES5yVVY+9gueSsYHfrJgMr7wncqfgptewbhQhqWtVjMLz5q4w3C
KDUyfrICBkvIwBIt/255R7f8jJb63IsXDj4qgUlgu8Q5fN/9Jpfbal7dKldfZWoBR+TDE9Oewvft
i3zOJYG3iC8MKvxkEhyN5QAWrWdUk3Wq8Y2SAGKde+jjNMSgzU8yvFd4Ovot0blDYeXRkWcwCNI2
XVR6pgxoYuflA4VvxY7IyWhtVzqkMCOcN0xuXv8fRF5Zdd68WXmKFdNdfipS0c7v7OFFZJjabo09
QRjDSHpsDC9h9KqkzYlbrmRrdgKjND6825yR9RyTjLGkx8nP7RhazU0jJ3YR/eKh6rAY/YPkzJYj
LjYv71EfplwJwlsDWFsq5c3k2OJprzQY/1iGOrRSsnYDOyXqRUxCva7yH1Ws91cvZCUESzeXJM/H
CMdph82BbKHhsN0UFIT4cwHynW4z7LQQxXQOdm7BW7HW1Td9fEdIgui7hI2QnDNwgTHQekCcyOYI
nIPTdNujcreOtzsBljY2B7EEll405Kv/aT+2ZA8tGisdKGyFQJmXwAFvhyhxoE3wwG0VaiTqZSH7
17CQc4ZpyvTjs1zPUKNjetfGFe7pMNCv7rwq5nz72LHrjDoRNMGUvUegVuE7Iy5O4KzTlcWhWAMR
cmOxdx+Vhi9cy+dI1bk0zxUjGMGka2rLQGqHRsN/+k4sRWJn9EFFVzCQOWHTNh1jn4IhjMd4QCmp
AV0XvNCGqsIO+v4W06b//XgYaRN22PioF1V4HOYF24C1qGfl4zgA3gh/zauNFEpZQ73/vb83KTyr
auxOiUruyXHbnDjrE51NQZ1LxeY6qSdx0Zlro5VbKol+Ijzol/s6L0Gv74NK8hoZuzz5CTMhv6rC
bWrF6ngAuN+XzHkI07fbdmve1mcpmqtUvyTv/QHlqevTtzzDAi+LyaGGSKtxYlIRJnLQj0pLCxZy
tMHZ+UOIPQ0PxnBvIxcQ6leqRG0025EHJqcsLfgAX7SDw4ekOMv5zQmiNiGtMd9EhJ3AmmifP+dY
NW49mpXQjeNVVjYKvYhFfb46DSzs5PIZF/OdzoNimduMMacNTn0dym+veCJ33CSaPAb6jROvIYlE
xcrMlXoRNbgBIc7l13HfBy8ujOdLKIMorUq6eDgQuKCZPArAQr+jN/T51Vk4DWU06sUNtngDrF6E
QEMbD1mI0OyuIzJttvFBjrHfDwOR8fXTdHHAJVrHvEUYU99Gw2mFEsaDKjYxGpHYatRAI25sSVNP
go2F1HwVIqm3N71KF673zkx545RwGOPPXmj+/VxaZm++3A/QbwFUuBy/AnX20/NW7OisT/mvaJP4
UdtjleH75AHCo2sPRgEO+O/N8EakDXoMUcuOQ8BQ3BOkRwQIBFgNLLB3O1X2CP8VBB/Cx+sCZAZT
r6Cm9CcaZDEQ8kVY08xdHq9iuXiM9vPuMZ/SmAbpKeNTyHxua9x8oYCMcdxmFmayQjaZMagvBDpr
V5MBteocs5BPA5u7fndkoHdqEvQH2malG2y68hRbpY4R/8SdwdyC9nZuO1RIGvqcVvUySdAuPly6
MBkhUkKDnVZHdIScCi8DDJDKNTXyLLZyou8rspitadiFli7rFuGh6HP/PGspsCMwmL/7TA2hOAW1
p8lw+m8vLO+MMZNBL8z4NjGONH9v6UTzMMIapQVG49c558ZYndUkedkKjBhh/JYIuGRh/kDae7Ar
liTkEuMtr1crvV64BnIskEXlz2ARYjrWQfT3NaV9rTuATzKy64Hg3lemt1jcIZWPpxZKNbriHTVB
owisCBZAtmVS2/6/l1MrWCBFUwTd+P7vJvWhx3e+CDQww1+GBUT1eL9rztUy0oaU9yfUh+exV5AN
nWfHT/V6iqmTEJoKPF85TvCSpGEMgE1C3Gm4cB9LeMYbpKexbNtaeMzOJJECRNqiSO1YJ+glux9F
RLMaGZq2GNm3nXpg3bQNqLQ13zlLVBJiyug16hmpK9CMFrd+iD2aODvN7JV6T9UxQLFM2OdrcC4E
MXIntzKBShk3kqOR6f55wj036kM0RFby05TpTe4MbpVuPmUK5tKt1MLnrQ5YkmXTt4Ga0cqSZ6Tc
jc2vF37Rf4hMioy9B3zhRalIP3bLJfkWqogEX07OqyGJWKk10gttGqGw4c/q9JClA+K/viWLXUCd
asVB++uW8/iaQ8lfQD8wKVAEItXjDeJd9v2Mcs+RUDVFXHxUrQ/7Xj26HHziyOdBnEkoY2772P4f
P2VcP/8X0r+caccTTqbCxfKDhJNSDDmeXjS7x/iFqqeK8hOH0kHL6A77mqgLfcOUHkHrDJhRHiyc
Q1Zyz3d1HVX3Te+kG8nLQnevhx9VwYpJjRly/0FsF0ulY/MCC5r9KdKE9cXq1Y1qmkAuR40VAr1Q
srVun4MlVk0YkieAzUDu6yIbnSzWoX3b6dKiLRrdQgnuzjcXOuRW0wTt9T7pJd0h3bIdSDMMB0Sq
2qlY4TkPvqzq8+0IRROW5qzT7IEeMWT7pYBSW226ZeHqytOoqr2FVKoLLvhcSfpLUU9FauxkMP1N
cD87bXMSoy2Wwceu8DuwAiahIkpVLi3mvx4lfwKNQe48zAMPmUBoKDI5+mSRn8bjxYQTZYZgrnnA
Q17lFjgF2RZUoF3lPIiPjmAHcutAPnkmC5nv/0HWUbMNgMUbMSDP2xsPf45ru0zYjmftl/UQB+4x
q0GPqF3T0od/68anClj3EpY8WggrrB6KHspxg5e827fI8XzughXfA81kjS+fwulkAYK11bBnhs39
mE+M2czgaChjvVlakdrET0TJk2RMn5ZxFaTICRjrpcV7DnZWunNN5dB2iS/gJ6Hv4zQT7MD26juL
1nVCYD9UPmE+nGd7HcPB6mMeF5XKVpx0TFjreVKhQb1ohBqj0fC/xC932LfKmdl3c4s40j+esnUX
spe36QyY/ukdohNqEKmpeQ0z8QJu/yrJ5u2YRc8oE7jYnG7w9PHEpAELC/tIHuY8GezE1F52N2v7
ibNdLo3o/mencfhXJkGrp22m2pfcIN/eTxNsg5BeKrGdtLUVWUYE0cZj5XzJq/hnXFcYbXcAs71K
VTc962HNWiW7qpVvPfW6JvRtYPrqAwo8JAivMOGgBQsz/ifB4bWnAXQI4xcLjFc9HtnHQYuTadbg
1k4JDI7XPp37AYsYfJ33OEMNuxH/Cw2WnVH5MtN/blxpzicd0ha1+BzBRKvNjcmlj23HcVeHxdtI
157fY4J705SGhly4o/2FVRrkyQOvY8jwVr9e7IngYXSqGaMKtRvsau6ua9tYFov6uaht+Wfdadhk
b3P9RHJVWaiKJNfLcmIqygYquQ1zt2yw4Aruau8MlyvEDlQdiZJNFhF31mHT81az7Elm1+MQkmKq
2IPY+PO3hP/LUwMr5SLMXyrlHGPTmkfLwZdVltaMZDiO7qeP7Q8s+lGiMkrE4xa4bs7CBDBLqDvj
rElIMU9EUhn/BLNVLWNfQILJOVXOOQiWXDGBzagOPpQQmGU4ScxjYy3ywyFAbZp4Hpx0bBiHerN6
6Ha7wS+/WrMyk1W5xHA3GEIuJftJd+Z8HHNXOlSUOXs6zlNPfTKU1sXzPnR/6d/qPdQovClWyqdE
jmGvcAXW08Uyhp4o25Lh+h/+dEw/qDyfPCJo5wIS4elHfTlsBW+D9hRe2kLSlPQn3a6gnGibWZD5
E2I5I9WNOVX1wjpm8TsLe+SWk9AoJJFsELNaTMOghfa0XN/7U37OpmWGh9cZfvWHODyElrclGp3G
SzxV42fNcxphbfI6XdAJsL7cCRUUJqyqiZETC/DDKC/iBwhwwZ6TwksfGK4KU4Q11T3QUsUrHvL5
zJzfHcPXTBh0tGPxuL/RTtieOcCBbsCuFQzjbSBMUKZwie/zzPPZTsRuybrXp11yVMt8CCRihzao
ZJGTj27WraNdQpgouaK+wVpWxMXGDj4qBAO4ALKpjWy3BRWgeZ/VsWYDDHizQ3mpiwmROOspXaG2
XD5JNAbf5OSuWw8lnL3NPtB5ObvLgY8UQBlY1/Ug1YOmCVdjZJDKWI04Dv1MV0vN5uhrvDev2yt/
BzPRGXlhat/ncfF03WSRgoKoD8IAqz7g4MojxvuKTZt1L5sTpm91YEPLyV4tLfGI59S1+QW5oTqh
MBnS4+fguqrJsGHOwcoMlUi7Y5Tqm6lVzT60oUqMuRObzEKbAjzOv4x/tuXMLAahEMb41EU8Fwxo
62SIUHcYH4VEwr4lRwvfag3Y0DfSYj+bBtA4YHygPIZ/RlaFUKqgKMhlyhwy2S9qu0d1iLBMo7Rz
kySI6Hqwcqextv1gY9qr4queYyxvg8yePs34EsSmt/JT9u2zpScgDrZqt334YwioENxjA50yGsKW
dUewtwV+E+03pUKWwH9XxqeNS3OxskA3QlGPfkBchDpkZQ7AKEN4xF41fSw9Q/kLyDBqN2FLqiaz
H/1k2pyIpsGIzl1hKEhevH1Bb8anESwA7+O68isO0iBdiaSCgrW3ErM4REL2m3LSrE2xLFT1xNjk
OiKQbwOx/35eUvMYCFpiTVUvBXqHKBsak9mvhVDCD7dhJbjo2xvf3LRmiKOdEyDoBupeNG2+UjEr
xpJKHczYS1etLb0erZXgBRZadfptNHb1kVPX3iLzcCdQ2O4BC+VMDqJEVgNgoC8KonwnTMtsmUyp
VHXbwOmV5r+POgmnycTaiX/D1a4stD8aVzmeaABZf6kpv4t07ZVMWhmE0FCAhx5qGcbMty64810V
TyVjOaa9ETsRB7oRS/Go7ABXYMV+acdQu6/nFwKAa92X56/pqs8mqjAPB4V+QooalrVzM66lmiSF
Cdzjxrhi+75Au/YOTm0vSegQegKyJuNRadbPo9CfYRR+qjTx2gWFwJVQpx4t8fpetoJNkHEbmL+j
H2ZCwkXBUwkA6iPlQ6ZIeXlqEyqS54oIyqu0uqKLZmQ3+4fLmu9VEXBSC/rsCXXXPgsUkoVgZNV+
oRDF3qG6bhETaHVCx+UOP6g08aJWC86wqLiMS6Q4OHFQafijv1d0rR8iWvHAvxaRU1g/FHhhKgsO
Ia89yi2Nt1U8jssdHkSlP4HdupCSSgSFjyu+xZmaxClVOsp4wAzxscOtPr2lWSSuv1LkouzPQevS
kPfEvCIUjlVdE+Qnn3f8O8iQy0j/dXu0pkzIFrs8N9Ark3xl/Ef1ByccQoUqi5/x2qzR+sd5fMk5
UILzK4bLEQgwPs3L6DMUERlpBLcuHbfnv4Tsstbx/sTV6Ahp79BYMWiQ2RHzQBlpgIGfH5pDPeNf
P0nh2W+jARklsFnBIkWKNU1vNSUepPPiOMMJ/nWa4vXQoh0LIGzO7mFo97MReb0UnpQL5jdOOK7V
tks707muOY8KQOcE85SUTEGqoTph0SPiohERIcOK3dkC5IZNVXnvniRCfyE0I4+BPTGQKVtW94v3
DxSpFr4muKS1n0TPP2cRoj+vx4Z5XVVJDDn5uSfOFjcSxjzF7msLASoE5MaOVzbrvQI2Af2QslCh
DqVmtUSM0MBQ881tq3a3IN8tLWKbIlYBNTSshgRCaGuzpI/15fxtBIaYx598/9HaiCQVBTHns+Z/
UjJ/XJWwStS5geCc9AVyNtuLmBw3KCPGCRIvxpgMqElHcMB9MG6FU5+AQ5btuiFNaXU170zkd/Gt
8sHYrGUkokeYFzQYyVaDvUEsZg4chHSTkS/aLhdJ8oI3mqMCFoUpCk2oH6P4AtFNH3YsjD1WZcRr
IvI8bqKMwqWnfwLkwT5BX9pCi9y3nrHDeD2hPOiJO6o91P7jPBSYQMQpgqAC8jay/QQdlLZDWjd9
pLuVv3lWqK5eW3jID67GOoiwfm2E1lVKfIhqHGxFLwkk6FoDhNbkH8sKiHYpxUXOm0oLyGw2ms1V
4vVDvJRFVFWpmI3YQPYTWiZfYU2G1m+wMVprX1LrOUqtn/x/6KIpFsUM1iS1kNoKU2TntpcLHG6d
EMMNCbcMYE9VPRaOpAkC2Cy5+iwVXTXZ9I3oSZE12FZekKMAjseCG4RxXohl5omwfrh/DUpARfae
TAC/GnXEfdkATfpyUbcWLa5f8igG8uD3za8jmmC5LvHyK4rE8G+B6fuPeFaYR7lWv1uEXhVHwgqN
G0ceiOtf2yJNsZlE5bqfvYz95bvqsfFbLkzx9cSzJXo4PqtsaHeKemNXKwQIyaXuG0Ut5rst5wRb
cSPtfO6rCc+663DBcJubZYgQHpji5uUkT1gUxikqxL5ls8RK5jzR008UIVpQJrG9QprYIJJudv30
+mlPTlY4sKR2V7pNV5mnjzFdnhJGvmm+Vz+MSieDG22rOtD16ll9FCT1vgWAPxL0a7O5Y9xoWRgd
4jHET0Suyule8NcARtz5wsXZrEgRbcV7Fz2aLtEXbnFHZ4vJPmL4FT1touMjg8UviXHi4CTrfXhy
2UKjYN3kh1lQ6yKU3XZfd+TK9PSWJIJ9+Abfwofzno7VnX5Dbx376rm2uQUVmAw7+axtQFDn3pvz
3NmPmY1fJ1qelHXZQK87UeWLGOSJz6HkceXPQZ78LvO9nP2Ewmvb9KnUiTaxhuhfxqHv0WGV23Iq
rw7MorWFZr+5lf/K3zFYYZahjiazq/vfKvqcelsxdU1VJkGb+bsWsIXr2323eiyVlREeM3TGCs0a
jdIQz+kIZJ8WIaZdfpduLRsENmFx6di6fImmUvQa1TKW4ln19VVT+0ceJ6C3eiHqtkIs/vXo/DvB
yrYlkEwXJTpBJ8/SNFqaV5aHD4t/wY1jx/UTG1nTGKKN3R/NU31XTz2GEO7MTN6Www8E9pyWsfzo
hc8sC8e8dbl+B8JQtx0UaiqvHgRHhbQYkDzsD9A+1Z3XcRsW6BpxLqkUeic2qObkgAhyLLz65F8/
jAKMtt/ADindrWVCAm9ZwyWEOnxrhSf1dEG1trvXNeqQ5Hf13grHqoswaAgBE9lKgJ/7qk55Vl3p
oe8lQss3T+fCc7UHW4Kyb7650egKO4kwT4JaL5IinvvlqnUM8u8gxvWEq5qqlRniIKaD9Z3ad8L+
ez8lJHsx96YhpOK13xYWy8bbWzeoYyuHubpV4x10x7jQhqneAZjpw/n7r8cDcRW/EKdNlc25Uru9
0BZynWU/s0d+L3NS4MyLjxEh51j6V5DBW2Oluu6st955jZOb35D9CJzHsS2N/N3PFwVTBBDEtfvo
6Q3QqKka5sJayL0IjxRRvd6C/2PGHHA6eZhf9MYjnlOEQctoKcjXTDLrM1vo2qcR4GEdvxetTPzp
e/2Su6xogfI6N30AhFrh80pQrDYBMY5WdJhqRSxSg9D0/VNBbVRz08ZhbtXhtckPmD1ekb4rVCS6
a70ByNHLQ0HhdgxXn1rUPOtFWooRBYtuo6MqLCUXmE0uZopw1mqXEAY2QhnQogfEe579U/jPrkci
iBg2/j0cwK3+Ih2KNE2dUTK6v4Vz7P4Ff/veJDMEh6Xysq3jlIHAgHfjkwKhM8ahcxIeKcRaxvwK
PTWJ07ISlgEpqM/tMDBAxvVaedPA980Ai6ch41n41j+PXcyc3GIYUrhFcAS7ZSVc4LHjfRFEogFs
oJgpyiaCNLOl8OjHFD9Lwlk54F4iziYFpQbh6RBbzZV0iPGchpcO9A86Hb2KJAUyHcTS/Zqb41f2
oacb4rJiqv0nnPQcI6U2U8w8DpaKqGgvcnSh1myJ0rBZH0KQvCVfxkZif/a2W6N3oYU7lGTzpuV9
moGKteLFjltFJ2XZZk7moVxJ1yA5aivIc2DJAc2+16olVrcZ1t6+A1irE/UdTy7Hxo46hxN/ZrQ2
Iqr5TZQfDMMxfYF3JbGzI9NVxbDGh6lyL6rhU9Qt8Nog1s/KM1RdJBISd+HzJBPST4olE0OqC4jX
ZeKNKDheOHAhWMi1hg6CMx5zkjlW2l/zFMdGoEpW1NtHuV9O3G1jcYGeY0gmEGsfXcZQntUPUDll
SmOOcxXyA6FaFOMvaMddYYtmAKAufPWyw62vq9/BRY/g/df2PRUh+w4FJc15o24vN2GVsIasFAke
r6s4EO6FnBSycUrQhCVEcuukByGQSPr+OKiv946ptb8LsXh6NTQ4F7P4dqPuChArbHQCqhNFmxKh
k9yxn69ZkN8+gn2Ek8t1Y+GOfon1PZuk4rkNHa/kDpqDE2G/XxglKkXk8oSQtxt22wpzWijLnmC0
jSP6ZAY9iNl6nvKIzoYytUvTrT+TvqXZbaK35urDV8rtjzb671zYJ+kEC6GIs+5rAV4tUUU8dLqM
0+opHDSrvco9u+m7ZcPezRaUoSVNy5mzrQbmQSx4kjrAbDztAdCoLAReK0SQZU/xrXTbDUBB+GKT
mob8umz/K0348bdmhHaa+tFfWDVtvfast3+3IpAiDmhoOcYyssJ/NyfoRQS8vs6VIE4TpaxJJ61U
4Yl1dKtRn/ePfaxxbgR9Qy/QVwZ3hklCemOG2LbDYBI5PAXarPO2g792UVdMJDETPLm6WDr+ribZ
4KH7jOdxrsOhdbFfguxHIL0YIUqBhJKhLHryBx7g7ZLLqQ4F5Uw2mnQy/R5uVix64lLBHjtCsXp9
zQHiQgs0F5kYnRLUyS46anVKyaUPx65nFntmhx5s2HwaKFVvZbSmcuBA8nX0aDRLXOAZEqg6yK2f
9dCv17ju960l4fBEgJcVPBlNvS2qXNnjkScsXrZwSWorZPLJVs4jLcqgIZkRG/OR88jGF8L5UJMP
fj72LSDKiAmMds0yRt7STw30l+ZCyDllig7TwPaP/8Y7z0vUgoDzj+mg0/F5BU2eZLizYaYBCyNL
YVKRV5u4NcKtcbxcefvG/HI+BV8FvzsT3uzIg/DNsNbGRpRaMMZUtj6+oUxlbtPshO2aGHBnA6Fk
w2RyatOEbnFjwEDrYUNlWPwYlFSuinebldUdQ8Z0HKnq+hbeh+dF+0nYHfon3a606fw3tJH/yzSZ
HmVsLAUL6a8ym5MSoV8XHtrRs9g2/+7VWla9CNAMR23x0OY3v/XfM5svUScVpu767mmXUHZ5wDo2
6GqWCDvRXQGIdwo9phT9UmhYeSdDk8cuPL7x8VxsUiImD/+MBBUuy1uVJX66PXRrfhKarz6svqg9
6s37e+4PcR1saKdIYJ76Ec/HIQOoc9vwuBWimiNi2AcvrMazA0lwsdFTgeDNR8giCFz1V6aAdS5B
gEtdOD5FMElbXwduWq3NFDvsS9pKH6MZPy4WSbldf5NoRC1Hej84N9m5EMZAHHCTG2170JzlZyxv
Oj6nu1mXkxhUaqXCjfm06Y00B9DmQCVAuQYWZf86AeunSci60ENvbW7MlNdc7QXc+xggwFpWiyPL
zNaesmUncRCR/6qe9mwLh4XOdTGNPH0zcpOOINF9MyofvD9QNT44gZ0g9nHTudt4kGqUY61UxYDD
E1SmLUP4+k+1Y5XPMX3SV0KWpXmz94aKgi4aqFhLZWZdHwbUYLcbe0EMoL38EUI4cM3mhpH8qars
dP+1LFdQWtgs8CNOZHvxXVhAzW7aU9O/Q9E5HaYwDpm9Ur9wZGPousXUxiXc5ruV7HyeAjPRt2FG
RqYSTQD9wxa1f34up+72Yyyi52gnKSZEbFUJLtvWSfyZCAjVeSIGyPrgR9tepob8n1BOtYg3ohBv
dUKS3gWNrv1GRbR2bN5yN5WsGuDyhumSHgSVSEpv3uFTEpbfnmqMh7ro73v42s5xzX1jEIFbGlyB
mwmFvQtJOM2JCkyzAefKsWNsKwuDYu4iluGZ3t94XMw09FqhHa0BAmMXS90WOhHBXHxfoXLT+OXf
kFkBDQRChDowyRJD7lzzX4Z0d7iN8Cm+4UVllf67X9qpZifQ/gu6jNppjZ2ULxoSKeJLhLKEqbz2
xi786+h74BFUoEMkvcGlRGwx9p27cGq3QU+/8dr7aXDFKHb6Rdyb2ocjL6Os8ZANYdFLXLgb4dto
+RDlKbuX+wqlbIEmFr/mMjgUmoP8wzzE1C2Pm3aSb6kBgZ6KCcCR6bhxryJ/4EGDVHgfxeyIOxDM
qoZZHThv5eU25wDTjKxcwOBr1UzfaZsJ/VyNgdcq+8D2cREXVIdxVPCh6rc7xRizYs9YRmci3yeS
6cXG18GdIdyD0oECh410qwZSHocWVss/UrtckpfRtzJIDwfhDFZoYwv1x9qYm9yoR/qY9do2tL6z
hJmyeKNel8lxPMISvrEVG6pSBW4GDcD7agnhzjvK2JpSJNLeonaen93kIa69U3eshh3pQBWzOVgb
wBjzTYEIPGPnBfgGiJ7Pg+RjYeGYge1C+tJ01o7RLBHwx6a7gYsia+N1LoAR9boGNBv98XvjvnvB
uqJeM1dwNz7dDDgkc6rmeivKzGznleCdD5DdC5wJ6lREcjtD125+P2Bw4pZFzCgGopC2p6lkHyrC
XXFT4vMrja6OCMmsfCRIIKgoDAuCxsdcXPS+7bF/KT9vlMgXa+O7a3Lg4Wi56G7U3Qjbjf7F1Uu4
H0vWMYZrBDoc/OnMOv2wLyijOXzQjli06dwog4Wp2x7aXdSiLyM61g5k3wqfhln+Y+amJW5qGGtd
axpGAARMucRVXSVkyaYyw3nbLv74RDSGcpxodYAo+jHfVEtqZq2zKp+Wqyzt6BDU5LtRAchoBgdn
Gz6+jfzQuyYHLvxIECgAtH8Hq6u+DsIC7ysg1P48WFEW+pshoD7AOVnm6UFR6+MkjKlGV1pKYLCg
u02e/K0O0O0d05Bs7OaGJcvWWbU/O6w5GWWHML+2z1fID8EIfapCwwwNIrie02vWKCyZaphKSw+u
+jpbASYh+kHngO++ESz4ymPPep25yKNudq/Y9kxDT2+btEkAgjzU/2jLJ+OF1WrWY6qARSc12wQD
zkZv/WrnpU1BOeLwTa60B43YvJVZ4cmrNMPOavxLw+j130b4/if1D9QMSE0B+2WbEooN8+vaTFEw
pd2VeLA3+Nz/61IK6XL17l21deSZGQJ4D9UBnZqJsnRNiBMdIoX66nHlKxvvpofz4B1l25d46NcP
ddcAPNn3qFvHLepQW1iEnMZEoPWntt5WaviSQDcCDmaKnHMjEt+VCLgLNwyeUknOLe6xfCDTHyy9
lXU2o6EuqM4jEfEmFXUChvCaDwKVmidyLuwAhJx3+vRBY+3LwYH3JpJMioLDJZE9HZyXiBvyoni5
7Ql34AjePeRyu14l8G6KpK6rhoZMXg4gL8KPQdlHgSlPVrfKT69azLY5kCP5RRpX/FGIw8pYLPA5
jnhvNq22fu1j5UOiesq79WL4sRArbYstPxxtS4wmv4tLa9gARvE91lppA6/Ul2PLFKJbDBAtZkQk
bPTYEmhoI1YGo8ORLPNe4D1UFScRliWj3Lw/hxSRkk6RgzPAuiCibf1oJ5vnY0xPmHeUgPLrMhNG
2M08mXvWT+f3Y+VJKquIRFBJtLYfnV/FAdzMi83A4jnpaSR0Xds8e+w5u5IqqS3+SKLI6HtVM/oe
dE38mq5j++84n/riTMoBxKS7oUMt/gPhoIYLUKWWkxbZdxMLuwD6/K05zJOobdG80lGKzc8gbyG7
8i+e2juoIcMwcqTGy0swYk5+mMNTCPm8TgLh45pnLeNQXQnzghfrWzai32I9rjYVywW8k4pcugQw
OD4UrzyMp3MaU4QNGU+VqZsas1FKQSilPwl+LMjyPUuRLP6nXpD0MiNEw8A8qSkZbt9NpYYfOXHU
JJCqxf3z4FYVSww/NV8VqU4vNgF2NKJlSGnQ/O2/IaBSBVj5J6S3dMXFtxwDND1Ajdo9/9Ci/y2t
dLyCw31TbQlyHcJq3HC53fU1HH3l0Y2M4yaagr09UBaL/qpo68RQzN0p/VcRYf9/bhNd/gswCgrf
ud2Z1DVqWNThgSaUtLx6fyialsWPwx+VNglzL200yeEEtwij07G0XuWvZ0go7q1MGcAeqaKUJDa2
SgBY2Ph5m7H3QLSky71kChp7maZRpHHhQAyoita1klPMn2P103tJeAMef0QHmdq1ICUHy0Ad3M2o
aZ5GgTRu6gvOU/Xs+l1aur5OOCuP5YJ91HFJPwQNMyUllbRqJPK4mshkjfP5lO2nT6yLTedq8HhW
IQyi70i6z7evG9Mz3G7XAMDDRFnsrWPID8XjlAbEIX6jcoaEJPWcqdUFSrhPuLs5d2nDjaXPp7bG
0QyXON473QTk3xUbY4qhrCs2D2pnz/XvKHfjFBD6YoP1TJhtg6lagnQvAGQsc0FNQDJI3+bi2zs1
xXfwMnwvoqxDBU97C7qLrDabR680oZsz8Y5jkFnrdsJqqeb6SCnLcQYJBNQmzQDRRKSQF2yPfs1z
rB56pJU2bGaQMzeAKHFg5Trm1dA5mFBfYcf/HgLe3ALWrSKh3G613ewvBkkAYSg0xdytsNkYqiru
i4kcFA7PnWPdxucWseSkkUkM5ipQ8JVAp0i8u9lwrBNQlhyxX9B164NUO/p6QOmgezOOPZKnA4ON
kYLpwyEFbRJQqdeXlgvL19tOyToIOm0CBCCH5Rm5F+oOC9exGQ+T0/aMNNOibwk62cG7Q9Pe/ci9
fxe/RSqk0t0L0ln3CkL/Iy0Q9o1z2NbLyoZISiswYd64P0vP8PXaGqzFo8qiLPtKyBEBXTRK+tIs
173XCG7CIDKvORhjGaKWLfwEGIvGJR3xGcqplmoXShRuHet4P/JbKO9y5AgHRJUpAng+Tco3XJ9l
vT22n+Q7V4otWTM6Kwtbs/A90HOyZCmasoBr34hxICFChpqiXZpDvAWFAuYjc/0IjwGBdjm9/O3V
b3bAoGIdi7lDxOKWE+r4CrnXjObRCu3v7NbBV9jFat6dFxPVnw6I2RGtVUXfYBrJatBUPC5bKZGY
eNbecNW4AS6oSitc3LILbfSlUCSCprCsoIhLT6BvcLoCHnM2tDakypjzZu3zBTN822hsnBBkKdNE
jQaoCOe96X1UIGEEvcXeAEdgN3MplmFgHhUwgEgqoP4Z/HIvkee1Bqrs00TUSJ+tLefv7X6seSTH
kd6t2czbuxR5MSNkohPHmWDNDOR4Y+mSdfOCeXAMjgTsk6tklaiFbsFkXM4jkJVj48sp2Nb3YOwh
T2C9Ni7YOGtyNHw6iWmKQVSs7gq/9XzbbvWy5A6sRrwDDqxh/a6bUc9qR8kA3VAX8vwKViG+r9bd
9iBWTn2Y2NsVg+kpTvpyyXjrVj5AYdCMKdmZPz7dz6fHrCcYqzAWInhTWHAKssTyFRRLx1sWrWQO
IMG8tMKdBUZLKXFlE/28ujk/EgO10wviT1gXy9soFG5zxCXW0P+khSt8Cwn3HbwPy3TECIrsn7OJ
qWlDaIHEp8CwvcrdisbC4YLOTnRB9Rkv8CtaGYR/mUer8qdZinS+ZSXPVPcSlZbMQk70CEx/Tsq/
UkaxP8V1NG5NVSUWw3icPkM+RRHcB0hzJRSNPjLY3F6UZp1UTeSILJ8l+qx750BNU85CA8Inq228
ypt7ZO3Db+ruQGjgrMvT15MHdhkSQU+qWGWcAEqCKrfMZDMKfWYnmkMRfwXEmUwyJFo4nMr3xKeP
ZHi3FlsgOa3w0nfVFSH0nx5Y5cDzKItrX3KbHwYO3/Q+tUqahN8bCHDNpUbjlsYxJo6V4NgYxkpN
8WH7QQyw+ZBr1u+/HrPp84HkZWjtPhlAc+zgRjZsHaXySVCywdZLh7rm2Wy6HXTNpZAS4g1Sgka/
5upU7RIWLAJ0//DZmPk8TePGQhV9JjsHAElbXC4T9m8G8z9n5LSafR31qjXLqWarwCxQImq4U0xY
nuTxdeYSR3yMjB7pwp3m5xgjjkMGTdv23HR/NPD4hzRjDP07fCwxZIdbxiiS88JeJ5yVyByC0rxB
P12Hm6sbBe7z6Crp+TTOjgLudNswgerfZF93q0osiDDAsmvMSaf15/u+4LUWczv8XKpQp3Cq+t+H
B7s5XfgWCsev4hQYULYwLl7sy1kmfCsYStpcHdn1cbZMKiVyIodfUinGpEYOT1sftjYIP1e+A0qZ
zJsT/lBRQIOmH0z9luVKDNioNg5pxHV+mNLF4ZbTOSfWqzXNfhM5oJwKl5q575ejL+9kqvjpAJ4X
WnmyOYnHZkZ7EOk38Sxdk202fgObY/NyJgZZ0wVo1vsSkSsgpnbsYQcs8x12B9FlRidoWKulNDkJ
MmIxHvp4urRUnG1aFhSVagilyNQ2R0sNQU4DR1iwC1at5nC16nVn5RoTehKY4WZ37a+i3bwXnRWX
2d38ITWxD3fFcgWhgMmPDqhif86Lt03azKEBjk8Ffxus+GuEoyScAzUK3cxirOY4QhEySlwMIAlJ
014hB4R1Qw7t7CfalZ0tP3DgCnYbzX6zZuL7iUXrsEcXAKVpqJRZ9Du/mnISJU6PIabQbarUGQKb
zyLKftzTRX8sghpWK6ubjz6sYqLL7S4D9UW8fKXKsslefwDqAdZKbSMopxEikvghT5UUkm/lhHj3
s3xzNEwD4hzNHgjO4OdMbCnIdStc9ZP3CtlrTpVWMRnQk+IqYBjRyooqHAFZqgZzRuODKIjSAtWJ
3W/1l+j++nBQap1bDlwKZnJBP/bHR6teDZahLAxrBhiQxnjXfO3owIE5I4f+r9d0i5p5R4Z1ytV4
Mtc1x7AiSXAyHruGlo2htmjVtRbdbD9hAAlqqZ84S3xNTxYPA37It8ZTFJPfSspxergAevm7MKTG
lWnwk1JygtvBO8uOHWPlNwGv6zxbou/uf0n0/dMsMsUY1QenrLLC0wbSfNGBxbz0vwrLeDgZDSk1
nwWMuIZXLg/3fiCNbA9wctEi4FzyU5YEE5MSokmGFMcf4pmsC0+WcVnLI+eQ8VejlcJoFR/rE5tA
YAxEBXZ66tQ+iIgFiYRGdTQQp6DhOVZwdH1eQfS1l47sWRTbhj8dhKFTg+oRCvrS4PnBlXb8jMn4
5OhuTDmT3F91Xd+4AMSlyE5TIm/55v63zH1VZI5N5qaiMbhz9s8nFhaJIKpe6C6mZ3tkNtKj2/CU
Xh8t4m9Jl7AWgibZhwe8QsG8/aZwTT940KdWfgxd3fX2kY6L90AZ00Dfffpn6T/hAuY1FGWllokZ
Qc04uPfek7LUF8mmOXWT2dnyPW4EXKPz1sWj72LCz0E2TotEZT4GVp5Nda6HAs4/HuljIeC0W7f6
GR8uJubD34KkgkIb457VwzUMRS+JO0BuUtL6JWIVjdCsxNT7Evj9XoICUi0bcDeYO3AYWOAYzd34
EE/MHkVn02HtPuz15lIZvDD36zA0rJs1pbWYNuRfjFft/LnTcOYPqJEoD6YMPDPwHUKFmkBqkqzA
mfUAuXVqxI7fUSMbUieY9zlF6C3i2ZEO7Z0b4tiR1S/90xFXPJ7KcNSTunfWvMzwGFqFg+GCAIQH
zV0Q/nSxT0MPP35s361KkpsFoX/t6ZGJZhFfG1+3MeqwNyZefMFMdJ4NmgON2Gc2B6gpKwb6i6N/
ieuy/i+e3Kf3yAJhyhtERk67i7w3H3AHSLt2BXCTrtcM9F4p3nhVJMB5XGxImcOETLyBQf4W4k2R
pnhUA2F/T5QQaPDkFnJTwOCjYvqMrCZbdxRs6KbaoIqzuREKlQSfAr9FFZjFAejf/HJ5Vne3DY0K
w0jqEWeZ5SCO3Z+hYJXLKFLbtWC/nik/kSqJhSDxjtkFgPFdBToEgUpWBRimCgfu+YaSHLLnj6bG
Rh/TrDRs3e+KlcZkufqQzaxmdI8ydilmpLoEy3S7lranXRkJZM3T0E4ZiWaCO+M5vIIDTVrXFgel
RmDiH9WVfMFZePwP3ZBcHkE0m3ZHS7BadcJr/FzvGE4sJHoK3vr8mCFRaQ012uiwpkhKr69nAoY7
tdApX4xGSyFPXtDYLqyJvlNro+dWAOacrhvW9G9K4MEWil4xH03gfM26hI4e6RfoEJEGKUUFlovw
Ose9G9jtitOPBetmpLVYpHzIFCYdJHnWVQOwDNvt9x+sztfDQwELXT9U0rMLlZ6ZQxc0OU3sBGmQ
ZayYoQ1CUchARjzAkoe7aQgTQPUmSIRhOxyZyme7vCKBe6oVtbqnkq6VVFEsTn4kUduvtqlc141v
P5CW1rVcrhromu0MRDzgf1m+vG2vru6W0MlKwNaAI74EbI7Jp06HiTv+Gq59Yeo/jyrqyubQhA/1
bglzfQU+JWN8N8V6g5JYf8kgMSE/k+0IaNMxu6F1Ib8OOpAEUwlffAik6ELJp3eZy0NWZZhdhQJu
dioJL5saZ8Bc7PwebOUHg+QXttKWKFdjDfYpCgnVKltcsppWlgS7YydxHt/jY0SU2q3J5NMBnzAn
uDnXGERieeGG1uMiy/6SGChPraZ1CSYhb3ugRVN5AYgrNP0qYpNjyLXp35jOEi3+FfZStTRq5Y/x
dxvAryVqVdbXOTaQO6X6fewOGetjOwU1htAKT+rvBxkWtBrSP+SHkT3LpSzIYPVrwklT+ggBasiC
2TT/paskgOrKoLAW7KqSbiV2AfMc0lLDFOLIBKgZDws6GHiAt0cjlxOY+X7LCSlYNi6D0MuATRv3
1nvbBNdlOITAD/AI9Y82OwpA5vyeIxfYsLLN4/reSpp+YIeAwnjpUIra2IIfMVCC0RbBrZtwkKWO
lOUVaeYSdm24S4C5vUzGFVGVJktEZW0eSH2M2cfZpcn+l7PxMIYpXAYHF5PYgP6I0LsmkanmtgNz
VIeQPZonBVBAMKRKZ9F8IIDY/rc9KOuucPV6AbGJbI3oBEsp/+d18w05PcCCEaVwkNRTSwChKzBj
EbCjNImL/9Hpi3VNMSDN3ckjAe6XoTwzIvaLYyeiumzGSh6nmiZKph9fSsCh3sAOj9w8uGlzBCo6
f11x+7KMjpyfNlHi1mVG0yuWAVtSj5QaV0ZgFFeGRGTLBBj2t8ukx8T/TL6OGALaszibGAngX/1T
rBtpQI52JLU1P/6hsrDlSKcVWPrgAxi+5VhTUbr8yg7sVeuOKZNczqOcWFDkFcYlEOb5bl6cnw4u
h6FlACtkirb9VtBdrU4u9AZoHe0iaT8HSABZGsErmbZJHYefSOHi2ImDwwROaxxyhklkvCrpL2BW
o+Fr5SeXAUDzV0otTdXOT0J3Fa60+Lmkp5zlsXC/i5T2qN/vKAJq5QLd+/T8slQk1Ug+A05Mq7wR
X6fFtvrrzxqUpN/Wqi1XpQFYad6RGS4Zk9Dz69OiclE7H4CuXXIlEqZUHYyrVaIXTXYLfhbR9e+w
D20ZvNeexO1sF5UT8kOfm7vKxTfWCJtRO6gTz5BiYs6beMeyc0cyCpSWo2dZtDiBtAs4ASEWauZ1
8ZJ4XOe18bJVQVAuLqWuQT+v6FjRTH2SZRhm9Y3Rk7DmMVOwUHlG0u1mfdddYu1ImNtJ4iktUOO+
CHAzbwDdPdftS/MdRquhIEnHdUi6iIrRgTbZov5pbRsG+HgV2qmU2aXDCNlQLHMXF1OkYF3DNEir
ommIrLOsQJd6SEQMym9DDbaw6zEQ3/uhXm4VlqWUnPM26XdkzwBJyfVnktr2FiBxSU4PjMvPsBHE
XkXUempezq/7xb3XLoocpXmVAMxt8xbihTbknO7oAQOJhe5jfs6s9KhkqyOw9Zhcth8Qv1EPLHYp
yCHRJ7uOdAeLXjNme+SYbhOVmeIyBVSpFzrlPOwjZn5bu2KMbh47L/cEQ+Q9hJF+aFE04XCC1Dkh
eblO4rBcsaClCI0wTtAe/sOtUQ62BQlqzMjVSB8ARNLD1BmM762SMPJjzCdXkqjG0EMaZg7tLnlJ
YirdVVtaBBoPSE2wXv98e0B0gjBYvd6cWo3nePHmLz2UFxeLjG4UsgAfZhE3OyKEvZ/5HsLUNUQ3
kQyjB75KNXU3+jlgJ0TUDdqiB5FR1qahNRIxAwGcciNyHC3xRqfxboS+XLAK+V21PshCZEkA0jJp
+MPi7Xgx9/kS5v0j2hhH+OQUt1VaDjiSVo97E+zolYKky/U026CpJG3bTC/QB6KR11liTNtGA9Rb
6BzwCrsIzxKSFuQVWpLg1+kIisbIuJxMTWSNDvTDsmGsEfb1M8YqzSadCV2OWqYtgF+ckAk5vp9d
H5Wpqh+3ElWNf7HsMgKZv5fXQ6K/LYDekLd4AZjWzgR4KLmd/JsPv8xMzg/H/4+YTl/r354Y+T4H
Zt/vub09/E/hWlZj8lv1v8EF7Cn2nQFwOA7imv/uRYJKUaXrACmO1DTnLdXCAu8xSJokFow/jtOf
pFNSRe8jSWPSVsCbbZOfi6Tvg8EC5c9KzCD4PUXMU/fKa7IJZ37TBg8PsFFhSf64dmvX0b8hzihi
UiLV1L3nzeFPWgRZfWVEYbKHJzCIXPaaDCOkNaCPQkZ6u7kqeaG8ED4Dq8+CapC/6gp0x4nNHpTm
/agTcM3PmoXSpV24psfjkc+78pQYbGNy6LVuejIK7a7COaEu57Do/hdYCqgvr4Uk3TIMvn2SA47N
cGZWJctTL9Z45lDjHRD1M8018wu/TR3pmz2doELNRHdRsbefCWmz0OZHhP53lGG/MAOMDutPjKuD
d71bJmAt+EwPpMD9Ag+tEMej+Bv67yOJJVjb8dgRIziDdEe8RpVDioTMGTUWiWcrXpHpthCJj+47
uPh158I1kKA4rUJWoVAaJ/CJaykNkIiI3iYeWf9h2ZaxahJUVOwV5lRaQMzxZrS5/domSdDw5eRR
Rc6czCkdISF/mTQNa4LImYkOG/8P/PxqRam+ajuEuxsOr24+rSINYnr4DwO9M7AbKFJu5I95/q/a
bGSk6Q5KD34BrgbphJSwFRQT91xEXFkXKWN7T1Pb5T21wCcjtiTMIotgrQq/vm0uHpodkQUvsf8D
IPstbBdGDaeNoh6kGJ71xTe26A+vTRRuLgOj+jinVa03xIIqbNkDisFiNwgtkb9LVlDXQdULXg3K
A2pUZ3nLDiogVc9ri/5/vLIZfrrs8J9rQIFW1hKRgrILA5mTIbuuFGZ2MiAB+EFnYC0HXbfUScsS
t4a8Qr6Nv1KJx4SIKaN0vIF57TL3XgeVCN1a5K5blpuLYADC8/+NkSScq4o7+2yWx2+XT8CXYbJi
jopSPRljzpenX+35TbeYwWbgLhyrie2y6CyrbHFZ5vSdL2yhCCnVvxyVLq4HhIf1ODMIfimZ4+SW
FJaROogx5VdPRIaBsNxKgCYbDdfWYszHXciGwzkAZ4zlNpbI6+9YDxq3ZQJt3h7LaTNi8y0fWTrQ
Y7zyHlwfDe/p8UsrQ8HOk02YGFicffmfkpWW83vC5xMzgirKw7bypUsb00STmsU20Kaau9b/6oVr
/tGJqM6tP+VHhVuYHbVjOWACTY+mMOrEtjbw93uMOddr3gGUAcEkXI/ofzPgHzipyVQTyIbc7QSp
vQIAzeCGy2x6seWa10GQ0TulKAQV3VUEkmSwAQy/WkWMSMV9+VMT0WvaJreVSnzgrhoUuWqsbCxJ
zphsCRSurdCo86Mxzg2I8k7/upem/nbAsug03Z8qVbOsgNvVxbwD+BMq435ULaN/MD1NR1+csu/Y
NZhrnNyEFl6oh5YtgGvR7WuHZrWD36Q99uKUMCCKZnnj3XsMuh+Q9WjepfNMNJUZU0F83uDZdV5n
BbLo+CZ9oDG4L1e0tip78MQ5lZAQVUH3Q7FHawmrevMYpmzDQnTQIKyVkKLW5HltEeM3C4V5wlsL
2egB3MX738OqrkEorgG13lo4bVtdlx6WSeIzuofZGqPD4u2lWgyQrnEwL7quvzHcw/3VhJR5z+MP
bfmmCxc03vcGxDeo/H95dDgiDa6jiKs4HyxEzBo76bC6n9+nmovDMvw6C37e1jwPtHdF0zVI7BYI
U96fCok4C0e2UOsZeF0KDPuj/uH1b5q4oFUnCXDHykMnnuCFIl36TqSJlVVz1GPC9VxDHlagzkDY
20poAYL8cdATmbzgPYXU0SEP6rKY0lsJMAdnbVNjs95zc8IO/Z6sBpnDetBh1qMiP4y9HImgZolv
i5vIq2TIvPuxy0v5bzzTjuYpSwQWD0r7ZYLtfT6o3782HFbShigkOxKg+2zZViUSqaqp9Pf/fCYA
uYLsHhLvFZbQMyP4gyJlXqHiPTH2E0gZKLhmOTapZ7qumhDAYm+eoMnjA+hgEp5j5YSkIW8dlPHz
+VkWiQ4dK4A/KK4ErcMxxBRRU8OXyfu9ZFU3JkFs6STxORAW6YqxcVnHiqLQdlJaDGN2COz8i/jZ
BOvoYgwnPjzj4+QdKapdNobYSVavob368J1AUlAm1/YvsQQSJR755Z7SIfyx1iF49RvHY0GuXNm+
baIblRNY+EARCUVoDJzNLfgr7cr7lxoDHAxzPCLNzeQ+RQuyHoy6VqOhPwbFYpH9Uqw1sUyTCkvi
H+5QGecoFR6P3zecIBSHt8q9wmjtB8AkAa++9T3DWFQLkkznhXzOgUknZCzsXrYxIJviT6kFpyyd
/dMXtjYDoWj6F2+CIc0D5uBC7Jy3qtESGwZMPZn9/Z7yp+Pdw1beEht2kvzmEuYPqfvNFoE3skMu
Jb28p00NRNEE17mUPe6YD0B4osPPrwh7cC43qMaZSpXb8nB30RW+PhA6RKvic/Te9Mx2flKNsHmQ
dqTeW/jlVTmeFjLsBOB3kRX35Jl8N6IuBIiLAC1mCJaDO3/YrzZ+jwV/fl3SOfhgnjLR9Z4DB/Yw
kapqH3vMwDK8UZXYPzy0JSRFhYYMQLhg5t3GJU5kVpzoa/h9E26w2jYLahkKbiaotHLemcPuTU6d
AXeg4NFcVna0zitrAGs7uCjEM43uPRSr8RG93O9qRxYu6iia4aQAXMm8gYNgXQG77AeNJIxMQ16e
3zH2UKF93EgLKOAc75v7Z7wBgEku5jZjaXnIzXhFI7y71iXIGs5uB6tWKHGLLHvKF/HdDakjRaw6
F+kGrdlHrCVe1CKCN4jH1Jz/ggoHRsokW2RAvhMJB1ohi5o25stMQ2wtUgsQse4s2J7zkaAYlBUb
3tvq88vXDwZ+Cj/mTG9evsAHLrapTHb9/ySz6vcJUrTIQPmuK0e70iIdwITRaRq9B3ZRwSuMk0k8
85TjT977LdEappkzArLuu1h2LwUm0iAWS8qGWN4SjqNaXeme6hlaq7tMmccdRYh8iyO7S+zyg6bF
MF2PUnxHG5+J3la+6VPjmKSsWbvEkYOcuBEIS366Pq/8LvwPtk33sRzW6z2sqO2nTIpuNE6IGuRm
JrhIvx8RZ7Td2UWve4raXgiqc8yRw+gB4BkE21sd8SauQuzgaPu4BQRkcLVK/ZyLZZIKauCIsd1Q
AN5TOsVfGR5eCJisdOXjqRykkKLyLnLY5wk4unhL2J8wHM7n26MaAUZxIMP6cEfKcWsPStnW1L00
6d9XC4L7ikgNfqib2bZUZrssDuo4orxkzbiYw12x1i7xnTCNmcBImSm2Mq9lrvgf67nfNkLGkiVu
/qN3pVeL3nEZ8DaDnwJSuLezok9SSLORILZM62ncxlM4uLhpxPV0kV3QOnxjUhKUZ2hgz+U4TC36
oDtma0bEbchoVPIYFiOubyJakuHTFbrBUegDzfn21TZcEaLXTAuD0qp9WeeHOkVxcLuuA7xrT0cB
zjELs53/GB4CYit9CTFFtO3GTODTPzyoWdE2vpAl7xfFD7Vf1/ZHq8qncPPeserHSX06sEc/VJCF
oBdfpmGafOyAaF4nLkW2oWXqKb1hwUiienEhQriTtKTBOgRsjivgQzbzI/Tm0EPkr54MmVwdyHU9
H8gzdi4Oceiq3ZyG8KOR7ncnx+DrxF/gIuAOiKRTIcfxKPDz7d0NyJzDWs0qGLrK5StZzKvfsIxR
xBFkRG4efLGKvBPzFeKM4s9qj8qCQdvcx5ll8jleJ8Kpvm1yFTCBMGK5Bw9ABTLF4ZdHb1Y5F7/s
HQ2JhAPGaXtLoJOlPAG6860u8mpX8P8SKFrqSoL2IsRLwTYnrdvtfohiF8/AmMh8V7mL2zPkd/cS
yxJqTZ5tpz+hinw2B5ylH8zBhhm2S9SNOn8wvOfKoUqyniCceVBvycQEkHtwm/Ute21FwDHf3VBJ
nm5zA/jSXwTQQuSPX92b537XOOd9BGPe1evuRo5kKD4fwXXdUKWVds/l+L0B86/aa5Q726mllKmK
Pdb78h8EMPKc4IcoULRN8EKWm2eS1AO8qBRn7sGC8xXAYCOv4FZAekmCF8ixHoRtEyknyJfFjRFp
+KX94nvswPCpOSPC+fb8+JuTu9kmXTHow8n9+AwxhmwqpTTasy0gkCUbJaljso5GeoCMPuOP9UjG
HM69lPONB8zVRc/RitPFvFa7ZgoW9to7hSbvtG40dfZ1FHAa0nqyWNIcGyGS+TDkravWTX0/W0kd
XhosHD/rPkStDeZEGoFSTkSLNpo4gOZ7w49lS2s3OWlVt2VMmMnUSBTO3xwe+plKZyUjM2w13EkB
BXNs0wEveRZftgvTFLMoI3o/sN+6kB0M0uZ2e6TdqfWHjWp+VZvNm7L6OKJFjqooZ0AzfnHBrk4A
HW1yPWs/6nxbrkAmq87I/lUowc2/lAUZp12RpAaRRhj2WHiY7If+bp3jUOlIH5OxmL9bDPvfmVb7
gceITbX5NbbT3X5X7s52tuhZFqyg81HEhwtI5Nrdn0FIe2BJmrfklwgPnFXb1pa4u8E/RfCBp+Cl
13NYEzPdcYWLKVKMk5L+FRrBiJn5W+1cg3bOfbkJM1K+iSqKTg/qEHdqcixT1G3cREivA3ljUCsd
3d5T1hNyHHPHjusyu6DTzzVJDj6ZQ75+jgpcTlDjG38b7jvEAcIzkO1sqpXs1SiAn2rR+8WCm2JK
ZrYmdELR2pMM5CeYJ+j96aU6BjoFksCASJoVRqSEJcP2SyDUcm1F0nziOlVzgcmL3+Dqs96bg6Es
ssUIrsb2uL8Fgnj+b1JJ67ai9Xmla1mVXZHqQTMUOtXWYmmKjuodseMthowslhrCQ/dznZlegPG3
1bVDHlo/jdn+m2HErthXzA1LJ70/0DbnQTLSAIy2W20/ENO4tt5lMwx8lEbMh6zmZMLSBN354Ptz
nPXjCRcNlt1ODedQw3e+UINaEhenwfbn6vIvg/2rttlUOSVQm/kELle0qSwuli/hB9fIpG/Y7Snu
kheQMv/io9XDanbJoxUEp68E3ya3U6nlKrQMvYrktAW/0a6mZZz3qSaceaonJXl8l2wiVwdNIkaf
kVdTIwln9BwDBsO0qV7nUQKVo/1zEdn2dkgTNVoMDfr3mi+PHYYjLyYlop2qM32Z06thjtAejbxe
DzM+IhADWW1EX9Rk0m4ZJ4Neo0QKnxHzz2fFmEdw5glByAqSCUH9c8BZH91n/EzMPsxIluL+7ahW
itZQh8HonzOEcwe1kRegpx48dtO7DT9PAG+6MclGOnFIBaQJ9ecmR9/caNLWDAJ5xT5y8e8dzKDd
61tULHjzwJgjeW53FhoTZOXih9cRYlDhjLnv3ItnK0hyzzwHysGH88XUUYb5NgiBdq9JYcymufUb
w6T0gJSPMEVdqt3nPdezxVUFRk9V7Hr+gs0CQob24W1sYwZQjfLgPuR7vhxb7DknQf0Qr6ASMc0G
kvC1DSCy0kpsYAglpwyuzYU5MOdMNlbutvenOLo+4koh9OZGO+3y2G1/ULv90ZVlkt99zYg9yIY1
FF1WOISTNBDTJod4Zsl8AGJ/13xoNziPy9iOrh8qiC7fFl/KmBoZIqwmnt0pGVLvE0OFbtmOsWUu
Q69vy8PIXQ72V4Og4NHamimdZmep5Yk4ZBYdh8+c9zj7BNW/WUgHBB3AuZBgcwh2HXlnTit5ACFD
a3rC10x7z62EFWbb4VvHOuBIQlLv95lT1biuxUvT0ZuQqHTlbWZisGmePhNB/WuxdWMAJtmyUTqa
8fuHRrVrBS4YbcHHaAlPF41v4CZNutkjqVfNk0b7w7Pc8868GWd5eosJXPAUxZhAGTDiTT8tprhA
xmHUakm8+j6rC81hEynC/JSBEj3ovHAAkF/fAjhK8O15jfEbUX5u45SQF9Mg+edL1uMH9XbEf2Nd
j97FomptSMb1/Pljiu5Rf5+0euB4MIyDM8hBnKitT0F3Yu1WtG14U/0ZnIClEDI+VHLi3wxn2gs7
DRRg3Yu5IfC14SM6EJ5Y/kNzxeGRxAO5P6LBDQjqK4j5m0S194kmnjMR092aZ4ffqeJPQCwbk265
iSGm7vJ15tt5N0qUPhdmX25JWL1cfLooJ3VpefsYoIDU9ZQmwNQa/SFx+mdG+8WzceMgEAzR5mDX
YqGXIoR0oSJDFBAJcgEpCVYvghb5/C0if/H4ENmgl39WZowFowbCLFCJ9687RuIenxGYtQctoi0U
9ZcUPkDzIR+8BBruyzryO0c4n9bUMNzSjmHa2YX2gpR+qrUErdGYDFH/oHd/2R4yaX12O1WEjj24
LWoLWdUmMspnNqDM1AGK6MdcAPfqcFweojw/iTPP8mLzxQJ0RQ2QVrvf9wB5187vCiTgtcDOaHmO
iKR/gysvEGyfmBQWph1mAnf1YeyCQWFB21ypQmdhrqvY7WwBajVzTNBN54kJA2BNRnJU5zF8Yr2S
xUKG/JpaS8P39iYxTa+4+WgSccczneKRvkmdsH/A7lyqj4FT4hQ0RPAS3w4vRavWLNUzf0LvPmBb
Dwny3rMRpuFIxLUm8Odja75ked13VZC2w7PqJDl858othrL6OpKeW44PUErasQK9CkGfKr9x2tpJ
qlnhspA0gS9gJ2r4p+Ny8ZTeDeCInBZVEdn3KC02fhMo3OilS0/pjM9CzhlRddulOcbbl62YjLlq
ebi0uAJsBY9C3RrL54N3Cg00Gt0FPn3q5pJfIngvKxPl2P7V/MrWR3kgyQvTic0KZBu4+ou62pXo
0B3InrjvpZ+Psu2Xw3s5OXtApYUdBWHjep3Hy6//1ciuDXzzU/OrwTy5ZzI9hbQhnXQVm6RaoyC1
lA0qSvdIz990afW5rV1rvdwIRAR/VvswobeCLX5GHk/CjJkF6x0G/2Uo90PVglQ2YKTkaadVlkAd
JLdZPz1Ct/gVDyyyE1wJ9xbjBzN/vThmYWC+SI+610sbgEJfY+r11uW7bXr/UmQ+RUUYJl3iz0cx
toZHfdbWG50MfFw+f0FP+Xp4dS9X8K0x17iXomdMFwhwHtpL221lGbmPdycZZEicLi0yqtWulimC
Tg0BkhADYaHitMgNT6Kia+FgS9dKOJ2uZQ8rq8vCX9zazourH3tzU4CNG6l1PVTDjnOlP1ebpv+V
RowVBkwsZPcuZo/pDzHwgf28stzRKNklYaEihUuQUhW2gXV3jQpfDunIVHi1uBLalsIsJIVYJ2TC
+pLfUWzgdMjfSJ+ZY+7lx0hssjI6IsbESN7+Nkp5kWSLKIQVQKwB6rHM3tSPOqez8r4Kf6q9hhwS
g3I5RxnAhBPcKza5BMGc44xuA9gPWg7rS/Fd0viITEB6A4AuSJntyfsZ+nmT3rHBUKHC7w3Ur6P6
2XoSZDOvFqurCGVKe2Aww4nMVCSjaETUX2v/wwAYqE9ihffjLSKF+VFhqW5UHrvkJ2+SiIA6HxzH
3GnHbG+0SbWlBkYMukH8GIA4DWQfnuTdj0U0HeFtVNk3/fr+ljQlT2wumRSUG9G6pz5ye9VrsHBl
/zJh0RFoXXSmFe0+hYrp+D7dF2/6YbLJjC3FEJD3OjSKxjGDo5Tyi9DVrFRpDJQiw+yJxWO+l3FU
MeT9nH4uxv9UGuYCUk/g/bTQ3sD/W0Rant7ShnsYLEjUsqC77lUeeMyiko6tX4nB0+xc6VEl9nTK
SxymI7ImN9gw2AlIZJTJWQc08S+O/yJCaUUgPRWUVbHTzxWlmG7V0omIvwskqxYItnoSRqH9ej/B
jqR9zVPO3ZU9USWb3L/GDwceaAKfv36DnIi6kmSrIvhhl7MCyId+bYbImZ7R8ZczFHMyx9afoGBC
BsE+FZ8t8asRHIICzUYzg+CvEZmnS7heF40MWM+xgAQ3PoVYgfoWnDkQpq9pYFvkuuRKYYIk5O2B
+aIeW4oxh+vnSYDREa1R/XwYKlnQFZUq2AVFMzLCzIoSqIsGY28swEAbIQ6FvudPRBfz58Teu7jL
Gc8cRmJ49oHcW5G9kSkOdcKiFkH9lSGhBu4/GecGVWAOXojaHKSb5esv96mifhWpe36/Wgj77ppa
xFFTVoPy8t/gPI0k5DRu9toh+Y6ZkmthhyUrDZe/93c+NoPxqZLfnRLmYthQi9l0Efuj5ULliZC1
SYr9DHu0vq4LMfwPkMYUwllY95sjbF86eDXHvMw/6eRduQNPmxOYrIXmekaUp0C9smq3bsem5E5A
OCdjBbjXaN7XiyCUMTsbQCsryHvGT4aloC4Kj438s0wDyOSM7s06GXBDCUWIpARYsRo/fHJ5MHw6
hY+NlDC9cpi8PAuNpvVgpbXgGIWSymOWyNgDYGPynUbU/zjogf67WsKJCpUYSNOKZgX5/XiYbDfE
oz/VreqR1WzGg7wHAu+APRtKAhUhCHUKMS/zwyL6Dj9j7MgRTHES5UU4pOs0R4EKY9aQK1vI2MS+
NbEdIcmsWrVPItpv8idcdtaqj/g659ccV5w5rVF/YWRV3frwZgkHG1BpjzyTTa4imRk55T7pqGYW
iYoAh2EwHV3KhdSCv+fNLd7FFfrZRvvoLXrEFz/QP41gecY4dBzsR7YYi5j4AveRZ4mYmoKXEdbL
LYeGidgCXjzFlA6c27Vam7+Eo/+nWVGwYpw/87lZa8FXL+HUyakdNz/NUsSetgiOtjp7kOY3r0Tr
STMWZeVU7HyOE7kQyKzvxv6WBfkmRJnRVOgpk4CFmZosnMHrEsZcYYE+GvSeDuNAPIBBt7LCJE28
KmLZR2axbxC2g7q9Xf43+kabP+pttimJBbJMeXu8G1XtldBXvA76KSgx/nQFUICdN7JRR2sdW/IX
NMw7rDfu+1VfHN6gYwUtZDRXbICnbZTPimuYGi7q+Wh6zxPu39MnFSdcm5vEilw5+GX9J/QgU6tD
cRAcZCijq72IlhRc0u/5H9FCw/0cCYURpAEAbE03XT+D2VfiHBYLExrGZIME4rOCN4DX6MLOe+8K
MhA5DYHdIPp35o4yxf4u5oCc50BFEVS339QqQ4KKXfEoZSqLQmQN7doLaCkAnOjiL25SoGCba+VB
eNSNVwgt4iVdrtXj+qTtDmSPlMf1eLBRvbNqdo5E1/UEV2MP6c4Tq2WqXWd6SXovYure6KGpxVE5
aWofMwK7fhzN12kSmurZTHBDJWt6mTzlGt4UXinEph4Q9rZQcVweFZfCSMMWEX+T/ZrUKSTCBX7b
S8JkARqJnlsPkXsAyfEPX9DHixgEtdGiFAp61jfnYmmAcxqiAHP4zzbkBgSxPL5oaqxVU+mPzw9Z
uBGHYD0QcpqBR3Yzfyp28HidPfjgscoMWMJzzjanoxWL9S0Q4PVkuR/9HZyMnxm1EBqxfxHsa5vs
+ev8EM1lQKPb78to04aU1ruJplzf6/n9IeFa+ElfFuPVigaICCYcdxvXOqAxDtZML7wa4ekYc/Ef
BZ1I5SYLjCAG4pVaSQHBXbvFYKi54vt75FcmpgCPU9LUVBoMzTQDdRQrIV0pYG20Z591zJrGten0
GIAUvQHYQW1YwYG0Xu+JzZ5MYqTbPv7tMeOhGTO1BDpAZQN0DAlZYaNMQ8UzJahIL5JcGjEjTW1t
nTxNksOz5tFDGTDslHziZh9M5u/MuI0UKxoKrLg7fYPjxN9Hwzykk4EBBQMZ3lPc+jWTPDUIId4g
o8QrzGVXnyEjJtFKntzNa+VTQLOzH1vf2RHCsNdAhAv1Z+ySGCffBiPcufYscC95sUw9cGMf23PF
393XHt4rNPDTnU6/LRBN+UqVSlf2k2Iw/Au6kdiuWi62Z8DcASrQOfBbPQGZU/UFhMoKq3qQBcoy
VyPTmwVyrCeyOStoDbdx1kGxEpZXqViy0CvKUQVwrmiXRXSTo6T8Anf4ZeZM/WTmumbaNEel3UGO
dTsRZDqdrVVriK7LuuGamMABVaWqesln8n2ASVwo++BjsxGVbDzKLatOrXSfa4h2Ema+YxXv9yva
mcePy4j+m2dIc0/y8ueWeNUFtL8OzeqtYTpx2rJyOTbBWH+9mbddg07jeHoM6jmi90JXoJ3wCl65
71A1wTrTAyMAKp246svI6svIsokRavF28ZinAkfw1O/kcUC9hwRL5FofI6pPsS73pkt2EHRbEdEB
R25opS6cMy/65VOj408zsoy6vYMz/e8E6/4IuB1Xo2e8FzvSRh69XZiCFdtMU/X2JpJE5nYwUY8I
tgWLo7XazFInjXETWs8CYgpZHhWNNmwXPbrjOPX/v0N8JTt05lKrgUBSHM+qrxuCukmF7Oz77Lsn
PAX+p5VmmKjypNam2g8SRnFlp+yK4QizMp8jn7ifEBKlDUsjnLQwU3sPBcuv6p1GWp7hLdyVvpu0
xERFN2q3iwDDDgLbALeH8K7x8fomsHB9fogZXmL4A0M05FGNvqR813SpSM28J+BSqfkK+/FyjrOc
Fe1LFDQcoElOuugoScK0H/Re5910EWuEwaeaLk0hV4aDr3AEHGrH6fPnzXc00aKT5FgLCLs7ltxX
WVAljfCz7jMiFdLxBAkok3lm38XJBCchy9QTJ9vI2/V6RDaAGlbkvG47Fe0KxmCodNbSL+QlHqKW
rpOJozYCIHTBXWkoUkcrv9KFmgXS90A/WZ+IDvwnsi3DMydeKub2n9QlLQ1fBCh+kzvmgMyyNM6q
Rec/E1nDqjdOCLbRK+RGy6VJmH7mU/lS6HUi/ZYjQvwFtVvmO3b1wLYoMX6fIhJJ5T6CSCvhJmnr
DYoXd7CwUBrgW+rqd1mlMxqnNC1nMqP2REvfeqbdU+mOPvnKKjRHiIwAURrsQKSChRtnfrsg7gWo
9GZnMDi1MSEXykmA6zsZEXVOReOrbJU3i3QLBZxDC/lYWGkEeBUE2gLzlps8bYJgFGN+BFJH143M
tikSFv7oWfQQTNE/g+srt+CdBI9JV+OdbbAZJTQ7X9DAYgHgOP7ePLo3ccbaEXXyrcI3k2ztcTlM
wjupK4p16vAdB9cuQd2B1tWQoDZ81rnKmE1E5523yecIBruxTMk4muz8uJeDKi5EolpWtqkQr5bb
zeyplFv4rUrOh99Utx4YEGY9/ccAdUopImPRdPrf3JAv2tEkabYhLtzZMEELQCAfye1pRLdBb0S0
KtIEGVX619d3cU2+3QnNHHr/30rDa4L5ISngD9SCR64YPv0lBROHGtplU79YTeeiuaryKd0vWAYU
GcMw84qL2XdBNvV6BjaKKe+0g3nFJE6mQa6r5n4LkrKGzGaS9w5/nwUdn41ZZ0CrediVX8kZeNjI
j3rUXk3tmafMy3AXcVbq7boi/w0R3dL1Es98l9RN53y0/5lfckyFMJxLzkwdoL1woZ4/XE74DoSf
WJ8sfodbif0ZeuIeDG5Sc6qxh9P+doRHUdp7Nby4hNFfmsu7Neh57LgjJ6y8VIAqegwN/G6qViZj
GL9hPQBurehNGYnbgsk9uR9rXN8e2lGHKPA1oOjh/qbsXPvWsEd/efOBLTbKh4HtbfuLHePWsbpm
+lzIPatPwITmejrkGdf9l5dK1fSlOO61izDqDATWvsEHYdf31UBAly1gWiM8+esqY4fzRT9gkO8E
3v47Lcpq0YEwp5t8lLlDg2LorvOqTOSLafgT9WEGx1F/uabE3cyy5N1MFQgxlYcpmKx64rmki/W8
FrkLWgOp7JqxoNsMo7G3ArUnx2657l8HixNyuAdfe/GJ8a+a3wy/1u4YxeBE7k1r2Bxql6WdO+NQ
E/toKrGhzwZH4AQj7XkXkpNwkRXPo/v+LiYOtf25xJMlbX6HQ7LiEnHhfwZ7iBpJc3j+wLrLYvI8
IdlOSsckkjqHc/S2xg0dWbA6B2OFQhjgD57iTkP9D+rmJhlkIO7yibpEExf0VqDy/nW6UrleCImI
FAV77obPQLfNxtxPSVLltcVqVgJDBawcLB+xYNGgr0aBiUYK8/118ZO6SZjl/msCwIMkC3Lbtn4b
9Hr0TZtav2bS+jWtUMNeN59rPfi4Qd1/XwEZ4hbiYdFD657gn6e7QsQqTn/ozBsS46JI1mBrs+x9
bdoWJycsPckdZYay3sfb4Y5olCMRyKozwWyf2okBG2TakPP9HylUg49/hLJmi3MK0vF2OY+eRVkP
BPS2NM9RKpcIQ8sCsj2TNNksWRKPxNfkY6jNageP8GN5dH/xXA+4IjAgYRBFXD+YAk9rfKkARgji
XZ88KRJHRL22Fk+SGkGJlpf79+nZG+O9Fo+sIF3SpU8KXkdfJhnVsX1eY+Fne6AepkEnTMfNGMFD
aqteoadqTKKq+FxLrSjdQSbDQLwz9Ma8N9uVFhnKuXwZGwC0ESpihX1eR+v7E3XJGhnGWHlqafvI
0FjkLttUH7aPrRr5NKzicnpePObc0FMou602daRnCAPMbaj1d+AIpkifdFC6wY8GuYGTxpdUK8sg
GDNxpJ56pQztzkpsyoWyWA7QBdVjilU/hSIGfQ5z5pgJ6LwdmjJkeUw0eZE9rHLMb2mgBvY8+0oU
FhgYey6YKqP2341hGWI4sgIlohyZtZ1qStw33EA8vdBJOZzEvwC4KsgBiwLMuTLAm5NQkjd8eRKG
eAQPizv/jNa+j0FuBWf7iY1gs3l/uy2s3aMTetnkOMtImygtu8N4ZBjAgbTAdUy69Rr7S0cx5Bry
wmksDooPo/4F3nesDdVm4wE1LZELB4tL1yy6Gqw6G7GuFi6Td5X8NARPORWbMXklBRSd9c659IBh
KxwfC1uTLt0JfTEcAbtCDZkm31YTJrhV8m11rtyDW96FIb+AVgk9Uh2EIm818L95EmvrNTvc38pV
18ZWwjU1e4t35BkxHrRGVc4jWpRxFRNPIQhtUCNR+uKdwxrDCw4hAsB9ryXHRMQnZN28wSGTcrhO
YBQP+jAHt7bpArrmzWe+GEaiZ+ArSmGhDZI9K/clBBkpMhb1Gsmb2cCUbRg630fcYGAbqL89vOzU
YIHnsil6XRdbTZwf9t3iBSDodsP2jdWc/FyXmieuUpNeKB5yNEEtBXz8NUZIb6+6Xb7COK5SbznN
zFPAT0hJkPHwakxcog5U1220UdrqA+64r2As9noaROZaaukBLbuWbjcHFB5zPiix+AFEhr1wLyN5
OeNwKUULK16HlMJot3fvVZjPsk3+qdm4ceDg2gZlUey8lUg0dAr8aAZZ3lr352uT2+soI47qX/Tu
jpqjJdI23TZBA2xurp1dLaiEG6CXCPEdn3b5oRzkhJxijJ5l2qlXiiTF2ZWrGM7fwq1tRE2xDMIP
Yl9qhNHahuznRQWN9zVvwM0fCLJQfZ8RwAMG5I8WlZY46woyDglFzsFL6oJPBC4Xlb9N+JIC/VUR
s8IZuMZ4PJEB74B+woTzosnAiCYIje//GzLD3PV+Wv5v8xR/mIkOLszFG//QiUxBj+xPtgg80kuG
F3iDgXLpCQuutwpO/mfvD3kzUrWy7FJO1eT7nOWasTa+mJ3IYwHzLhpvej3L3BX6EthVKKIwIGcD
a0B3zyzt+W08pnQU/R7IFJO7rst8Ks1Ib5oBFiPVti0brZJuWdVB2uk1b1DHPZTuk/n+DJSXI21o
AZ50XTuliVXvE1jdHfJ2A5ZXbSVYzbAyuGdYn/nn2OiRJScPJ1XvWoh70Wf/0NMEfS8e4397oA5o
yNh4ccPwDQuGzjGs0UcYI78YkNpk2piEYSjl08SlcLyFtyPmTacZCNrsK7ZiRFXsdbabBF8EKwyd
Efvtmc3CA2a8xjapaaIRAbaTrWw6VTudhfDWUGfbs20U7v2SYR6kw/cRGIrnRylSD5SoO9Z5D4KY
IVbCceg+JkD0wRaxja/kZq7SI7eF7FY+7eB2Y1aESXPuNWYiNi7JGZNEZN/daE0NBrjTNPfk40UM
AIFLIMxRwhIDoyBxzUf1A3tfiOAhZtpOV9EWv2BgR8HkvSSVrcZvH1tyN36LRth66+N6JPVB5Ns6
MV+kjBuugyW7UtcBKaKkiH79MNFCZWxMmb3i1C9oqMGC6VIpGBZRYUHwnX8i1O/6IISqCPQO7DKd
AfO0ai74FhV19GS3rNS2BAMJEsplwlZdrjhqxQfNI0KiajMn+0xG+0oddbJrGcEO9xNBbzOQeHOJ
dFvwscbb+iSX8kxtMdfAshjC1C947yiN4TsmNTXAOi88B1PdQEALlEljK/Mkeau0pPenshIsfzNT
68KvQS3rdl2NKwKzJN+Dy2AXB7QspFrm9qeCJFHsusmWWKzHNiRICnR+rFprK/NoPB6OpSvY3gWg
xFjGMPgG/YQjwELSzFJObWy5QaGqXeqW50/If/+l2aOUIVwbwl0srBOVGxYfxIQtHCrt97/yvE5k
4B7aCms/VUx2F8iEpfo5B8gMJ5mvVROi+sjv6r2x8usgq5Gft10syXYraBks5XgiCewqemugAD08
CcmVHqo+fpi+I1DQLf8LYvBLB6lyNKGkr17AVQ1FODLkSyh9w22Rv5uGBE6BFWkpH67BG/As9NQP
r9J8a5ut/xCmM9OuRigX+X9QXhxBt0cUTDXednW/gkQJeH9Fa31mPwoyn/Un4qFWmhcDJJvk3ydS
XEEHr6/ZW0iSmTLeCTuB8pIFjGnvW3/Mi4gikf6uXAdQYQl5lAfh8T+zU7gwxj0Anl5AKPLx/zjH
r/n8kP40vyBP5Gpl1K6ow+KM24qmbmqC/hgpesdy5m4u8Wz6Mtu0zfn6bb28IPKOd0sUleAyLtwI
R/iVCNkxRALOsfWx3diCNEUDtUV6jOVZ8HDJV0MY6pYr9qXo/3TCALVI+0/A89FMzGxXVORV0oUL
aZ7BOKPrCP8OJmw2VmVRD/Qwa6JIKwHrbuAW8hg7ikNqFEIukRL037+XAipxWt9/wlDGL5hB0q3O
MCbe4zsI708OiqlTvNO2P1N6rMQMwFH9+ha4lMAtz+E7mzyQMdnHgT40MjhjGp2G4lwjVWd7PyZ8
oduRSuG7ZQVs4Mtq9oy6zwZLURg10c7vDDUJo8pG/WvgAjr79Z5lvlAeFd6cE/X45+nGMhzbS/1C
id8gEKDFdrPUTPafbkojK+tWwdLaPgDBsAKnqQcaIC70w3BVB+lclL8oOkgHhSJEZxS+pOSpfchn
v2FaI9BiMlXp+oMkYzKxRCs89z5HXMiXPCQSWwjg90/YK42qeMe5UDimQxZ/TPVTJJ5xAbST/wCL
MIuGBXbJ0nH2nXj/ChvPGYPnlmRXK+a7mLOvvYkdHMXrpAeMuZNv7BQDDGSsbaTkJiaCU5fdEe8l
Yg026IoUPXPJsUqfT9XsNXkS6BlMpWO07y5o27h+lrX5vQXtIlIRRO0DF66LSRuQJFkiRP921DwU
1J/ijQXEdDhrrIlgXXGJG50ZulBF/mjBz7XeRT2rxqZU641chVT+ceZiwC97iSk0hoFM69m9Ftre
u9GmoTYeaqdXMItXsQB63wjvpWAFRpVDJq/vbuLK0Xj0Qoh0nKFpKnmf1FMy1IUaq8ya0HUDZooV
yjlPz5xqM7jjjS4rHn94yVC8oo4MqzlsN/I+QoXm5mC3X4wYNJGWMX1Vc6+cFiGN06XUy2Y3K6nE
ljcQYKo2ITczFV02xiuMSOnaFq9LlpwIVa8zDB3L0lL2fCmpAIrAdXnsgvaQCRdp8r7w3VMwcoey
Y3uJaKbyrpTxIcQy5CnKrQ0s8fjokYhQBwTei4VWfLAXuR6os0gw2YQC3dZh3i5UzzU+UEnjvgQK
kWMnhU997Wu//YKZBGfrQEs1zYDPZy51KyotjAqaD5PzYvoQ9Zx/gzDgeAHfrsKh5IcODBhIkglZ
/U4R9PGInfNVniE/WEqef7bb7Jx9VKR4qaDF1/L1QLfsaj2b/New1X8NwQTLOS3rEuNoHiI+bmf6
Nzqjj5PYZ/h9SyE1i3eMI3/lZ8naRSHSgxi4MPfSceaHgqE9Hl6jrpGJ/VBDxhij9Bt4NGeiRQBn
Xvyi/HcGpppHm5M689Ml83+lLfyMHBzpQ0fnZyxGfFb7UPQTsh138QOdgfyK1ULm8ZchgTuaHn08
Ab1gUP5q8jSpEqi0eLIMZstmL4njqg2K/X3oXNHgHiawlGD5HUMZ8U9Egt10h949TDSHch8wq5s2
XVHqdxvCwn/aElx3F2Iio3s1NFsvrwghz94uFz5bBtzGMlLw9abvQCia2F1VZls453SQuZESZ/wC
flkaQoeGRBI2HIs+OMBw0uAoLRR03GrRgLsVYZxQF5eYwPU8BCs2RebnszVca4xiOoSWr40s2eO9
OKUbbt4UkzHJZQlSXbVYtxUJo8OGP/ErWdo+RqVRKERMFf17ymejOen3hu1CPpG0P3UWJPhmKAz/
JX/JCcTae62aT2f5f7jAV74anEfCOD5+48Na6HY5NwrqHnKyKjUhtX2nQhOyhNYOADM1mX/Tp6lk
qkVTjt61FDF6jQpnYNtOV+5iRzcyGAiVpRc7mwhgVTTYCoeaMrEG1+wFvNBShSXwPUfNVgcKkvTy
PYN2sdC3YvRQgx8IS7A+lVzh0GTtFZMez9pYbcWUK10/n0SMLmhHhRV45qobjClA0wHRcxMERFGE
f2P83khkxXyptXGUKRCcr8lVhaLRREmzMyZYFCO5GcFMFzqFCDUD/ywbSZ3+OEWmq3G4PomByUXB
sXNdS65x3jd6smuJsFXSFd1gBPQhUUpO14ezeejddeu5OjQFbYul11qpxYAJpHIU4yzuRbg8H4Qi
Dg+Lyc3kaLVMCtTSKfCRzTVpb/HNKEPaWdL43yVVpSSoA8pPbhvJVHIgV8h/yCQh8vpZVZGUvyAP
VqCmlnpIJZxAc5o4lsomy7y/ScGbL7MBgdrNxVxbNgSt6h0Jna0+kDkH0YNnNAc8P3FghL72s7nZ
x84lYAD5PX2R+/NIGxP3EzpZQUEoq4sgkuRVZ+YqpwNQKYfKzsvZXMzTQf3XUW/IDor3BcHec5TZ
MeKkMfu0sHSZdtnB7MPps3UdY6GIYmsu0EQDwOY1RijlZQjzsIff3QlM25DDrR6yaiCZx5Gbrwwr
OGY6WLdh8YKhz9RV7QhND0u1s1GZ+oKlIQqLZv3TT3fpnkqJLXUtvLZyAgfQAjK7DyOMNvNZV5k4
519HfiBNWtZgcsuN+AYFclzRAMrZplyAdqSN/lK/xIwrzGdysqqM/eWeA3MLT6H2ZmyxjwE55602
APVrfu1vbXijvN92tzhchgdvYm3B22GvsHM6z5KWEtqYzyU6RYuw+GvIEayAMhcVlRfhkQwbnQVS
zQJU58fbLLg0gNf/gcjbXmBa/ynVsTLXclIU9OTn/QinxKocG5GKOnpUokFht/RnBAG7OtsAC1Ns
HQCFJxlrI0hVrl4uiS3E4+39UM7mxC15CAKJw4myLoqxlvBmbMWkjBApuAoD8u+fJZpcVBdg4cU5
fcZnnCzAEIaaLdwQZUuMuWY96hrmD+vY4ZJ3O4NsoKmQJRLi5O//G8L1hhofzO1ori1j9qPwDn17
4j53Jon9RMlKtegkAB4GuH/ngkcjrH4GfcnEEEytkVT+M1Z3/wg69KTm8TWPbqHqfWOeRcvSD4OM
FIFJT5r1nT3mqYVvR2KMUbIp8XfN6zUXs6WeYkFa6ScZHT1nVotj9PYczd+F8WflL/8VqHiHLDXo
JerzYXo1EyOReUFErbCUR9iGTgVCHN4ckcnf7tJGNAj/KVPRr9BYVjqJkBkntt5haQktmmovTEAQ
h9Gp7/WHGqOemPoDxYpGkVGnSYYdnBJl19UzHyHlfa9YxtqYKWzm9YP+U+ZZSafMkB3CkTAqHAiN
FtpljSKGNP2/L84tkkCzgO+jGkkUAnniMwNazB1x78dfXkojTJsLdvZPtM8OEArCc55GR5sXRt8f
3E7N/nT8dAmKxbgI9YAQYwPdw7XnzdhLw+DM9i7xswsxT3tOw8KYXCghmdBYCh0Jcj5AB+cI2BjT
0gof1KEP/R0sbxlh1ArsCQ/Tm+zh2nNUcHvYti2lnks7ZPQZwOwouBO5VKynTyqIZ66s9enZgR5e
99NPdVIxOnA/SpRNBaBSwPBRLa1rqHG+RX0hmpFr36TKxKZf6Ij/HLoDm3QNUkYXTWlMaS/oTjL4
fWwLie5G4UKsOJTJnAf/B3bMoKS6/CMU7/1jfKtH/h4+WfaqB6UnMFDwpKaD7t9tS95lr9rBgU1t
+E29Nua3Ut8mIgB/d27EvpxDhidaT0BJosqOLQ8FhItZubQFbGL1KtM3cJKd5oLQP2fs8gcvtCZN
e1EUpBK+4WFl5FKx+q/K6XYC+4+y8QMJuo1Pd7MOKNIUR7XASUV5o2K+gbXlaFODT2SurSrFbnkZ
YRYI/LkuqV0yXqVvcOUbQXXP74uL6nulglL2CRJ9TtTvXwq5pIg8SInrDyl/p0E1QBdx9bs+k6Cv
1w0UaQ2HOJbsruhuQ90uG41K3BxdtrrMdr4Gh+iv5Z1Pvw+h8MQ5dMeSLLsl0G3VKF6oJkdpIIDs
cYIlaFrhMcALXGvIDILz2iNPwrSRHZjR+K/ERa97ed9G6Uzm67mKCDbemS2JADWofd5FnLrMe/Ak
tXktq6XgVS4SEV10+rjAfFHUOV1wXzy1/xiYC6L0rdIxgtWOLLorNnKkPTr8/6J3fYpUqUD6LeZe
rqOEyP5aMRVeD/R9rSyYR1unWryuDmZDLBMBqEEJoU4E+a+PYvnQgaUB85m8gfk9p05CmMj/ucX6
4g9m61W6yjSowcyYmnnMJhe7dSwvdsGKI5zdmkWg+htDB3nAxEOvX2/dOZEVsRvBnX1ydI8eIw1g
DC/GH8Cympm45SJ07EFk+SIb2GOVHJi3zeGyUS7/7iOSnWuNerp0CbF+nz0BOEcYX8VRYqgixQmG
VtKGPi1G5U6C+1k3Lh4aJBgY7QrahI3K6JHMQmgLOGeIjTuitP9AG5F+WS+CT6ZAwFqrHfwcmqQD
gOz+3+GZd0zOOtfcPUD1aE9OrxBA0bTdi21/7TOTwh8rtAkj7sp7soPK0Q3WMqbX04sPUxyzLhHI
waeg6V6Skg3wfFEazvKZcPCxvOLMBQX8BR+/VSOxz7ZT8ERjDtnRurEzGrnMe22pU5mhkrAhNxf6
TDGbLTmUnFzc7gK+5aFn/6XiIDZTBCm2sMgq1I6L1o67usOf59QL+SGmkTIZGBZx7ZX1dWSzf7Re
Wx5m4DE8V7psxr3BT2i2bBJTMRrG2b9r+LflbkhK9crhKLXalRae1o8mPGYGROxe73fh3y381iwL
l5O87Z8QtXU5prCkWqP4Deuyk0byljraEmBwIvHHTWpbhGIeolUK7Wv5vPFPYsYrcSjHlSOCN1Nj
20zIIUt/knQeE7IXe6uAXxhdXGcMIQXalTseCQmihJJH2YjFmnPGb/1njnmTydFZBUCtlWEtE9w5
AlgglhMKT0F701rcxfGdMuXzfUnFi4y/F//R2C2rhwjyNB5oLpVCHJ13gzRRi1LLbUX0y6QTjCtv
o0jveYlp3+pu3qZxzSfZQ8i/qPGvrmbNhFLx3hDkJG5dHjhRq2be12URXJ+ZR8hy6HA+Wx6Ax2YN
mDysuBNSQCUfNxOA+wxERis0O3yAP9228WZa1DBvOvOasVNMaAhzkdyRIwh+HqpCSL+ngcdIAOUg
Q+hu47EMoPr2LDPAA3XaMEUyQ40EPpFrfZrBgp2O79S3lVGGvpWs6XN5DMFdOTdV/kfmbVVLYwEK
vJSnnNYOKTUlQdgJlejOuuyB6fOVSpQ0lZQWSEic5nOXVwPk55EBHWRSNDi0c3cekl6d68AuOJ18
/n4LkWiS7IkoLX+0KjXMG7l7wNPKbmIPJ/w04OhT0DPNk/R4MQ5rhdN6kvEZV/2q3Mm1XCBX/nGR
WL8dniVBquNI945cXcI+KyR28gFZvpv0/uqkCs8zKhErSl3us6xLcRbKCYJIBcRWV/M8BvNvGmOu
X4Iyw3E9hPycvsdTh1J9iXKvVO+GTW0Br26djU5deb3/8BjUNM3mtekLHvEt263pB+oibPpOxmTQ
Cs5Dff24g1PmQ5Q1leI82V1ARRx8N9YYcp+cH1qWk2i2s7Aoox5Xc29gzjamT8rkdjpKILyoBqcW
cnqYlCI36hZudY8K3VGIVbpMgUVjfEXj/30R6o8u97FbEON1qH8j3IxdUTOScgCipKn4ncPFAAF4
GA4/tJTJoSGOebmUX4LRG8Y3vRm5QixSODvjHMxqo0Z2sAC/UKpQkFW6wjjCKy6dDhU8vgB7MYaQ
y+2vkSxcyPhEwgETWqYHPJg2eIkvEm9zUZEoxVQNuZlAGs4/SNrflNWHFgPN49+H1u2et04UvUmx
I9pAONIqCA61Zcl6UfKTkNOEHL4ko6ylLm/hcoorirT6a0xNl+M6hRNhJHPGm+qqt/gnXdaE2jaF
kl75IkKS5OuOl5qWy5LCxOMsj1RvRDlqgaS22irGSJfPcdlva2WmbojmQTYiHNdF38d0kFag0R4q
R3Sm9OLlHa0RZ9y/og40+vgB5vnWrG/aBjuxHPnAHuMGPPpIVT2IJLeMx9PHfSZ2kPB+eFCBfe4c
dzuoX3I3MLp/NE+XLxrCZDh2PI/UgMxa4IQdoS8y6SWbpAGOKmm5uf5V4MHvWAJLsFateyAGdtLy
aZg2Q8lVYkf+agFUbWOjqrtB4WZB96kkzr8YLZO9RXtppURQSC9JGANFqUI/bQut6EBfpQeOP/GY
ml8R/eu8C/uinLbk36LAeBkpkM1sNtVtd3raD3iaiuzllxAEVXDh7NdKEur+sFYERWzbRI0NY97O
YimlcdOKHQtYA94EYLB0kdErNJXrodN0olJp8Z1xydUJSxydm+rEH5e69oOsudMyCdZMhysd4adL
1F2HVHIHYiVHnyLVQ90C2T349oU5FEmPQJKbvZ6uKwrQBprvguN72TWdkm4ToJdpI8IeXwMI40oU
uPyi2dmX1657qu7WrCoRc4MNY8y05rixL4zWxq9iQImlQPqua+Tz8SIGfboDFJqFaZs9vycrZGWa
0FZ4VDqwUNd6Rruc2yVcO1hTzYXjnJ9fo1adFUX1OZRJu5537rJaD3ins469W1cEsM8PIezoLvmp
DpW7f4eEN6Id/wUJsixoOfVgn3Bjp6lbQOlmrsf+M2XX4zqvhVIjRS2ydP+9kJU4bmJuwDjIDYuQ
4ECK1ihuyTlhru/D9nEX+ErwRsgM6lS7O2afNeGF2fcZUw2iT55NTVeOS2alcZRENd6a0jz3lZSi
FCE21cn5NfdiuK26VUntgj1IK6sMVn3rclfYX7ZvTZ7ms6kPxW9wWjstuSO1zIg81s+MFaWjeSw/
3vaz1f9wWirFCx8CTJXeDFFGJzdHe8LULC1mdsLvT/3i718ps4yIRLn1llVOwy4k31wFlX10FBpY
pFmFn/Blmr4xvUkFn0ksDmhQ0tPQfRyq0uhdPwwxStd4qIm2W4hYJsC2aP1Jay6/cLI2q2bHs7MW
tiWJpNyV3psu2w8MQaFQDnOsscdicGARig1xBd+GFQjwZhaQY+CvQL3n9/cJR1OTtF5NwjOKhNH0
YqXRQnJcn3k3tQ/lxSs5fcrKxpsVRafOY886Hr4TM1TNJt8gukDrZbJEQNlB67LSix8+gtaf5mxY
yqvhxr3raLVWtpSI6Poi+BodcS8sqB45UfKDuwVVR6jEZoR1Qx9LYAJANU3N0a6p3rSwpy9Bbuuu
/dQvVwmeeUi18W+wWbdwQIgyrCPZVXKROoWXzFjtv7s+/DadOJMdbbI9oPTWn1UingfRqc2/ufcs
UmFN8EdNQWV85wHaVU2glRz/nYPZJRoH4nPLqXvwMwdQaLYAc2ia/1l0YWd+HBfem7co2SjL7E2n
1/YpwO5Q/8uKFiQNIp4JX+spbxqmO7C3NgHsUUv/ADT74l4Bcz3yrfaMPx2FNjFT0HHqznk98j7h
644pflG6TnNZ2feFCXkjqIKaxiUJQ1vgFWer038iDeeuIyiExc+VBwAcjmPj9ZU5QdJHWVSSL3Tj
eUVln444QVIyrj0Luom/QvsNzHNxCSCWkHzNgwTXPQTKWCScOOCcNqt8K7ZC4B4SzEzuIcp3JFwO
kjkg4GmBBu2grOfeH3RSH3pj3gpmIuf+CbtzrK9uae9nmCScFFjHUbUNP/a/Z1HllWh0OzSD7kd0
qrRBOVZIF9sd10/OnbBCnUBAvy6V9uzZPvFivCjX4M6vLOa+ffI2Uy+z0bXzExKmgvqmA4Ws8mAe
HgBBqECLH8uM/SdB+7bUCrdpdlPbkZa9bb5WRghRST/7aG+ilJFpPkj+UCGMPwiu4/M8Dizo1bTN
r/iPRF/G8dWnL0SvGo4B2epxdDP2XFqjxByCThrGKgpuodplYJnyosCszub4it3CoDddP0zzVsEv
Kgi686XmDmG2yiaByphVZ32GRUpZRJ92IpdFL3qTXcOD28yOk+sU+8JSa9MAPe7iylYDfUupCMoo
kmsMRJW4+gHweiV+mTTEzzzyYJ3Fm5n2EDlBw2WX4R84UzXgIKni2eCiO/Wn07nNJksEe0M7kf7M
hboY0H4ZGopcmDIabViKwGjQYX3/TvXWy6zYuVWY8MkNRALCkRbb1wLH6B13cVS+SnRM1tUgFjmv
si2gkCg5rjWa9j6ffI03txocK286q44hw9bcJXez06PIzEIGG/rf9jmBgijQ90jUbyMDAOq1zWJI
WI0ecBrQNKj4nvnuxb1YYUcEo+JOiATTZBDdIexRvbpDMIKkwIXGkdkttfCGZnSnFV6tN+DTLBRz
3MZM7pM6G87t02/ZTuKJlIkhypoX6OpzvoDm4SEnGjiZAw4OBMUFTAzs3DuRslCYf13OmoTW2wxi
9KnfAax8nA3Ngenqe3Wc4m9nh7xbUVyRNQnEUa62typ7to57qd1jB6U8KNV3HQPWRAsS0mpl7CHj
Cpn4/dvDHI6TKa5rJJyZfbakerGAdvH0ygHkNVAm0rJuhoYMaXz7OtOFezw1tMoSRHZqvF3BO/Gv
oghluzRlX5zThCtESEsOEY5qZzPh2yAghW0VhW99tgXv4+wFeErLlHlIWPURSOaTuPJJ+3tZ5y7P
vk65a6IbnIN1dlo6Rbg0Mhrp9o9flVQ+63y8WBeWmkGDJP1K2YYNd/5Lcf5u/oye4y8jB3/3UVc9
vhR5fNv2H8IbWl3eeAUzuexflvFSWUjc50Hv3iX6v0TYM1IZb2ihHfkdGJcIY7CsS8hUNBjG3Rxi
edqpx6P00UIh57OhJnLm45H/C2fWiqfLiX7PreNn1EYUBCO2JqmmYJVSAQIYoVTqD1hYfWT5vQZQ
LQuK2LGZH12We4m7kFX6S2XFBkA4bossR3IyG4cfoy1pUcbOg9bFgw/YZyvlX/L6GusIUbclZpws
2my7lYTz10xtQFN7+0g5tYChFpah6nnjaaJhSyUS92K2zbLyEPhn2EIK8v/xNGoEN6B6EL7KTc6U
NJL0IaEM7R8/fXf7pdEVJFI3o4Zvzol3XaFrof+WYJQo9nqGJEDo1cugDhKXFbBWZAWPGMF7sbU+
+5r5QQUJ0qBgTaHbCXnr8xaTCAnTJnRR05gS/b7B8Ody0ZJCpyk4gYvchsK1lUzKCDxpj9KKOs1k
FqxiQT6exFFhEBmul7EDbcDV84HqiZc/mQig24x80Nca8QMR6Bj7KMD2v79Ufw9lseg68VWDBmT+
nL16wRQmp+9Tx/e2nKv5wIMHTJ2l0pf2x/AwZgg1rykRFM6niGe0kVIuFSf5uTff08q3G1zGDY2S
dhN2YYxzxL2xaKI9Gx3rOIbFEbE3h/w5b1M5l3V7qJKSMfeuz7IybcAXkgzO31rSBwPUL4pQDcWY
LA/t/FB00ZjB1CilmepV96RkSXqXashu5GfocuB+bVMCrt5NPN4xD1bfK1G3aB1l7CHcC6uxXFFN
rkpBwFn+RX4pV+ryjXR/0t3XmIIM33TS6ER+wtwK3jzt3xpDmYFbdgAqo+lfBp6gmCI/I6ihYD2V
rGNi3oX5sWNsllMJ9qJYAU7OzerBhDrFHizoQ/NNWUzJ4sLzP/XA18cq8CmVlGD6heC3lRZf/NFY
YAt9R5C35Evk86dThwCcTU1fP+SkLhn2+ZACoJrCNGV14v6LDHhliwnypsSzr4Wt17TyaFf14X9J
WhEZudeP1JemiDtl93b9Isf3ungjlDpNPXSYWvnmFHroC0X5aEWgYBHqVDqobvBN0FVKj5EF2htG
QtUT8UfG3PTlvbBWmYkE761PA3wUbS3IOt665WWT9X8qL0ylsCavFbdbknzseI1SogJJ04vT2r/o
omRC/y4jRlGCW9x29Duc/0MmpL+ngebDiMS5pPwjkX9ly/iNz8Hz2DgEGc5qHdGVBu8xS1vvVl5v
W/sCTCaxbqnZnbr6xx3DVVm4kAJMkKKvFZVNWYpmeQWlbz6TkhsPpWuArRUZ/nUfZLeuwAimMyy2
X+Bd23dPmpuu0LdKBRnHB5vSjFZQNkLHz6wGyuLLoipugMoy+gxVs4l62cGfVpMXS7mD/HmPB4PH
hvIMBTc96sy5YSFde+DX96tAABlKozd+M6QdIXMI5qk/w0OR33vKhYnBR/qj3SGtuu8eGP/YXik8
cDB9vg1yvXhU6aO+6RpAcl3ewJxT3p4Xrq4sXdceWLYHjNa7KixSb4UBIKJKqCfYP3T1Uj+Vudje
CsWAXyML8P7erRRsXAXQQ29wWLBRIDwaFj2QIClWeGOtgl9PbpMYCfSLfd8n93zpIRgkwpuuAh9F
hIAfEfId1Gx82+yivr5nVOyXV1CuHon/KdUECtb1t+pW/mCwTIiUomUOGBUHwy6twfBwXgk9qLj4
xz2kvUf9L7zD9+KVKt8JHYMfJl1TlTFMQofSLv1ZzbIbY8yYKKXb7o+48HnUGZN14K/yeHGICK22
OzKVsN11ln+aS+jNw6hqjNDUtz0H/MxcHIPGdV6v3H8+FRGfya3z96mFLBXqWoLoOVvoJJrlLe68
KztF7nc5SF4uVEq0JkvucXdGyAKQKNgKUCp66v8/fpykAo5aIEv+l3jnza8O3g9lAgZr6hePHtEu
efBoIWhpvgR/sHgrgDNYXV5I6t60ZLK7u5RRAd0DxfykbL2h4okkhnazWFnP6vvzIdl7q27qVfqE
sgFj/rIudndtoCQ+imhS0gfsVWw1P4+Df3BipnvlaamIXIyfg2fK73UnHfdSrXjRdLNMQEkycSG6
rT1aYc4s1kixj/NoruhM9j8OZbIM77pnarXn1wg4Yn0rrEut3blkIlKymeciplWOTbJA2und+Xn3
O2pQ0pgd+w/avjzM1+GiH/eD5YYKALnpVQwFmsseV+87fFO+J0ajYd4fvbyMjYRaq4eXnl9iS2fL
N1YdEZBXnCvHalqTGcv3NZe5vVnCKhlJChOLADsjx2lDjmBYWPacwH2aN588f92QBq0ooXPWKalK
OqV6SaqaIjl2LwiFzY7twuVun/vhlHq+/dzTnVUJr0wq+e0AbyMqY68/N/AUWzBlJ5Jt3hSMwsf6
ppfSlAZmpmryg4oOeoZUGpKuzrB1GR1R+ujXziBRkfx3yqTBb4MmM1WkGKYXRss1NmX7EyJGTLvw
q1XtqGeBZm0K0HIIGKSpC3/CSVq2s0xLbrb8RrQPB4wne3XlFF7T+51mohqvX7Y7Aqyh2IH8FkAb
XDyEgSS+DkyOS2dZgjxzj8gni3S9pMq7l7pn7o2HENJZ6/gHV8eQn/tjhwRE/Sm8t7s4mAYTfkjw
H1gDGdAX0oHMYSBsazAvqeLt5l0p7Gxmv9ZjhByjp2knIpW9IuGID8QmnOlD+o85DmSilYAwyYG/
Npc9hE624P6Tq3UXiVKkTZEXaJ70w120os6tmpOu7pc5Fk9cTL8iM9CDAaJCgKQD7743KXVDsKiP
CQUPq5mM5ZZ26lJQOfcVnHqPLqcGFeIReVEO/2yPqnOhOvS4XGUha0NnScjr/j/2T9ej7KcXoOrk
a3bpBwW8L8ITbkOIDRijOnGDQrOwBD8YeZG1++TMW8oBnwQu40cOV8NKKzufyOf2viZFd/1JBAIp
nuUlS1f01rb3i93lxdWp1PXvTeI2JdEt4K0jFy2Mdf2HHqybJ2g0K8bpw8fVm6VUkEWWZRQMHxqM
2hZahIIFI3F/5JXkeSHDUunp1TDblf851ewnPnZJSatRt2/Wqa9CZUm6vi3DnWgW4mOz7hM+K2bW
mAmFNqzSy6EssajL1ynFTCnkZcaRtwIXyCi9sKGvlrDaAPLGsWzeFejpOxl8j8+glvG/fCUZeN/z
3uoVzMzimT4tutI+Df6Fbj2GPDbAsHxqcziVQ9EW+g8eg+mltEwdPGM25gdlXghR91LxZ3mQAFHf
L30EwiDdSwF5olr+skMVwMMJ/c85sf7lnu+QeF6pLMvaTgK/3Fp47VhbkNLNk4znsqrDdMRQq9Z2
plOna3WUrOXypQsoxl1CdcTo0NGSxO6nPWTcwAhDVnLdd3wmZsLEoO0XFWr6ACyVod2Y7df7/O94
vrCAjmdZ751sNDyo6hH2ECgYbBpqp9OMxtXWroaVyv7ctI6zuqmz8mDSIshwnYTvXjgtUiTuu/14
YdaWhWelsmzV7VrUdSl+9z/Gl1SZ3hkI76ekmkjbrSHjTLR1E1kJ2440Z1yldvnDTHLYkf7Y/6YI
EMc8NArBhQWw/bokWoknardtkDZ5rcitLXDdAOKRcQPUsuOnVa2uvm+h241sgNp8PCaD3Fu3BBD7
jM6DH0FjTU8MDequVdBrdD0rKWgbn4UR7BYV4LaYGFc9P3Nky3nHyeulcRMgzLsoEpxVevuQ7S26
svNDT7Kh7kd4Nu9kmVFfBOftIUI5tbpqmT2NrRWEJSpd0XX64VI9G/tb88gUdHhNCfB5DQui4VCH
2f7NIRpvL61521cQ55Ly6nN3oHTUnjiYj9NtzcLhutztDPgwD2QcwFNz3+8pd4ChAK8IkV8cv6ZM
lX3IfeCAoTfU1NGl8X3Zn12SxfpzOlCNCw/meGZhrKUkNYA2ddLLMZh+gwDTsEl4XJkCYPrkhYjW
rQwvGEdDgzKQoA5340uGa0BMpxZJmxxOBpxDfT+afmrkMa9sKO5bbCs8vG7S7zpFrMnZZLTpoj7G
aX5GpdV5GZFmopztAYBt7KRUziffxi2p/FHBhveKNAkfP4hB83WtVaXNqayKbW//+6a/KIzLrYSa
RJEQuFdNI+GzvelEM6KncpFnxgRuhS9TNnsiNewVw62a7y1PjUWFIYGJHjytR7nOgS0YEo0EA6n8
Ykro7228PguVboiiwKwzqP9gu72q7vqL28y9UcN2UrGDZZASl35Z6RpWNQaS4xt4AnqJjTyDiMyq
9wywmoSn2w0ofzGfmYnfbPwsRIXv2heIUqAX5Xva/ASLGRvLJhRqUlGmlakiqHJWjjb08KhS3YJR
wrzG+sFerMRju03qJgiQSBytpBS19UzxrhDo0l1gbb/sTCcjIv27JjiI2KlW6U2wlndvhU1E5+7/
48dam0HETbBaevpToUDk9IVYsbzCYI0ID1KOdToMwdEvavPATo74OoTsWQoE8U+wZzB0Ymi4lulU
wqJqXHWGonx4rEsDfwn+QkLvCt35b2flKwiWh+1i7IM7sht7T6hvA1SSF46ha+i2cl94nfBwXCrk
m61TJpgfgXVDO6R0PLHdugsOcrzqa6+R1wu0q7y5hYXcOIGgPKcnEHiYPeDF4TqEm9SjvVQd31p5
aOS+h7/uAVkXo4pUhnXanwRHhFrI4zhEXuwJtx6R7pxRDoKjhQwl7Nigw1hvxRfBcRmxMbMwWRDb
EyCHDZoh0VviiFd0ye5VkYdabT+dRvp9zwoUAsscV/SMCX02zw/AdJB3dvoqu62nx1A1ooMbMdzY
skA89q4OfaowSIMkWQu+VeGr3jy5k6QehTDfwEgw+rHY1Th3YAeVX2z8gl/IgQks+g/v7VqtIfaQ
kpB74d1Wo4wwpZlBTpQ7f4+b20c5DrzIhqkoXYv/KR1Fln49ype0zG/Yrtit7dkF898iqrKrt332
BAvc/g5biCWmwoRskjfltOrNbcZ9Th/TPjEhzjEwTIXKBc5CH+4/A1LsaJ6C0IO8JMm1Fk5476ws
YMLeCYC/XeFTtddk1lP7OosGKutWejJ/2cPPC+Mt7O+F/oCGiCrCO6SXZjFTKKHA+jE8wlxlYmgi
GSSs0VHxlZNal3ZL374F8lVUH1RSChw1LVcvb8/K3EWI9Q6BaauvlIr8zC7OLDxHSCyXhSlngNYu
l3n5rmaS6bP6Dzy4xaPva8KdxpUh1CXv1i82gyprUMzxG2KqzPAOydVggD4nUNVJXy9jCHPaj4Nr
bx4HMFRQ/zHvZwa0DGeeWyqzkiH5nwpXMTuWEOmNDYAgxC7/0H4fa6IITlTZmAcClyfFC5krefBn
YQ3m04Lcy+Xrq1lYS+dMLSAPuhS949ddt2e3jJF0UxpOWn4cyicsd/dlkfYDS1Gr4BH3s9gy9j1P
S39FYqLGaTRStV/fXK9Zc35gLZYGHhpUBtJp0fZfiMXGwVvsphIVYLOWNNIEKP5cp169PJrpp6e3
qy0VWdC+QpoJ8/gr54fLblcm1zpSBYunbhQNVDxIXRu5PuyUixPeUL7T4kKe9qb10usbOcYt2dN5
Am9cPTLf5W+cFpCkaViCFCD1L0kdIN6MMoiJwZEUn3PV1+yZqfYy//ZrdKw8wwOgkbgQAYE/6/Hb
wdf8FMEwe52EURu3IgPl80Y9hz9raqp6UByuPTn8z9KrcDIpw4WYw8sn8ZUSQjcOaWN9zfxAoW3n
Y0yOBz96wca4IKN3Xy2eEc4N4eeI+WyRGj7+Ch1DYXeL/yy3iRQUxgWxTH/bfIZwwYgX7SLm3dP9
//yGpSvDj4PO+VsIiesaIyOW7SSi4TZog0yJlXtRj4DUIm8KPPW9wXAhZf93PE6D90u0sWt/sRyh
Q3bALI7fx0Rrw4LldRacysi8ZTNtICWZmaGr12TwbJkt8e5MSXBCB32H99YuhKIHNiI3ZyFl+p5D
/BiJSUfPmzoXV5p6XUvG6iPjwcdlNs6i8XNAQ3ayhsA0RR03EeDxdW/TpNSewvawve+pDc7nxpaF
OVoZFdCk3m8/nAPaOeuPQhCDEwopVx1tfxcjAgYH18p0GZTEl0ZHAmFPSW3wNJ9C4fGB9yyVFXrt
mfyjzO9vC1OuiGOV+0SsoKrBYO67evTT6aseAAQugP02Vxb7W7Y0DRZfa2KLMptkHfRaahglvI6T
KiIQ3VIpvlpfpX7LX4nbv9d7GHTgfLNCOxakNzYVJxF+JPojiKp9sjurQyOI0/oxUlDT6L8vSCTz
V9JmoWHqCs7uO6deNR0WRODUNKgX1smsCuTDank37Lpz/sNIefAH78B7QKRLgTM4xbHofJNTO1VO
t+R34VzZh1cqphXIInahabcSAKK9xRYGDuxc9tx+FHqwHWgkCbPflaCvRKOy7sMUBl5h/dGa0jzl
WQefB9mg1QIN96elATs4+QKt1ooNK3m7S3DtEuEW6nI438WVeyT4Us6FCsOIlv9etkGt/Y7tQ/Ft
VBy1s50lgLjbXai1QROPOQggvu+DET/sr7CNuvmtDYJrimAVb3WXZO2+D5Vk32niegZSJzGkiz3i
9DJa46wKw53ZwJovdeMrSolsloP87df7/18gV75aYx+AJYot8yNqAVvQeFEaQwOeFjZueLjlmuqj
uOKg4VLAdeB2CmSZ32heHTiuJzhlX44tmDX2PJDSGC40AyzmaEo0Ctu4CaEANoswkSmG+Xto8Arj
saJQJdIu5LbZloZ3akZ6Fy5pgtBe3rfRpWx/3a6Dk3gyCyyMBDK+BnmLE2FgbsBUDDaey7EZ9d4g
DPtRJEwCSQ69SXHnOmvLfP3S6K8rob9wHQJSiIAC6rDmdt0lDrev945HRKnbWusxjTLJNEodZaiO
zC/G5XGMTuMfY0p38RGOXtsrzo5LwzcgciQf0crl2kvCEqeg4BynBAsKEIKd8P2TadTaVF2YDR6V
6k0dgUIpSSWudOEKtx5LVQBrra+M7WkwSSeBhGn84u5lpCFz0V1KDxNU0QEBsPf9DaW5mt0WP3ie
2tX6cUlfweLjamUl5fPClK4kgt6fxHTIGQZb7LhhOJZux2rVfSx+XbrD3t+Ne/qlztrnY/2ezPUD
h1jpTeQubQpnvoUD39HWsaVVDtdxMaPPur5SQbRSaibiYAjZ7Ji1u6oXFU1txiJ3AKJAg54BZ3G3
gBwQLHjnY3lKVbpSYCHBx23MjozUcMVwNeF/XIZC7LEA7BaCtS1B2bXmzP7f1Zhw0AoUu3wIe9v/
V2MIdqVDNAkI1HzOCo3uQ9kVOxlxyMKs06FAcdoHdfCLH98K6uI+9v4moX2EhqOqNWREem/pnpDB
47WrEH8LBxdJzwBVe94grWNg02uKrMyPZ0++CQCa03c9RpPCgXLItjfs6nhJ5m3GQPVbbT1dvPF1
rtz7SC8GECJL1R/yRL3aGXg4CCVVhhF4+Rjolt0Y7R/u2W1ANEtKfYXgVWiv6fYU3f+LSln4jvpJ
MpAQw698jQ2ev0xvydiJEfJ18HUYrsgSFAWCSnDx9Pq/l9/fP7yYY6Csy0D8cK7Ri6gRvZ0ub5Un
mZo7k9ZkbCSfcImLJVO2RHkEtU/KyxjRy1DgOAgWIpw+JHFMvsrqdkHGCFa4fnqIZ2bFgAGi846A
0HTJqBpFbP8eccbgdpzlgsug6yrkkrWlMQRZh0erbblPk4l7kMkxeQIthLGVKhg6qW50JT7Czll/
sF7NguKtyfMN9z8v2yWu2bG76WzQZDQIFyAHU1B1w21Qe/aQCvtOaDdrtLsFpsomgjs1pg60pV9Y
fq7y3DVQHfWUMZ4m65GkIXZheeXzH4S+TNSx/unOZAEBL1QaXJm9ohWCFcwiWU1nMkffYD42+uO6
BCkutkTkB0nkaWwSQ3ZCCKyHCZ+cOMEwiaJYfsUZAFQNtJ5ausfXhDcddWPfBmlHnMjGG+Ks5YWv
Qr4+5GY1rKHGzg5HsNDIlfJUHcDqsI9F6zgoi5PBKPoBnHd9t1Nqq9qAibCzqZ3V5TlATxdEY9PQ
AwhSWjx7Aml7qqwN92TWNVA/SeL4zDMqK3NC3hJCEquFoKB3ATsFrcinx7GoNrFIq6Ute2pC/m4p
XD826wYr0Sv/L94AsmxYmkgSEbhk1kVOSU2jzuz7KX/NQl4QDgVDxtCKDOIjJxI/h77d1flCcSNO
YRK1HgChO/CH318DSEEauYnMH1IvBLkjF/ihNyd9RXOTFe4Pt8VFlDCASfjIn1vlHhQIPjAZZzGA
HMJgIGokGe2rY9WBe7PJUo0jls6jJQ7x0b974rPLS+MpM/2WHv0hnouUUHFL87sc252mfjvb6dmA
eLkDvfgJUPxCjRASzULf6U/BSyut4HpUWhXhsKw1Sy0f92VaAhMQdd+edmucZ0sF9IEgLKcOLtff
zzjyY0nlaHfGZZyWrpBvBYiZRZQCMWjkE6ynIp2JHSouUn2qB+EDsJ+T1rd9fMIFEWBPjXet6o4g
qP+SZxFdx2M5yxrFnHg8bSTbaFpD6axUm/7iQDap/vcS+WFopZNJLNBIyzoRLO/3wtPA+SDJFSoS
YUDZJlxGg99Eck7O4Tsk0tcL/DgyobUda0x4Aq8sirhrtuy2lIiR2AS8BRhL3iRBNgusg4Za1pIc
w/0brxG8Q4+RBV9xBm1qiqdfgmj0TTQkw8ZIpEmfX1YnGrx4pVc+1Cfa4NOfSMSwPBv1qJZaT97R
oNatJ56uwZn2p/t7FdsOKqI4wNtS14aZjS2PaSCSS46Isnn04m627Trj8AAhl7vTLE1Be0TKNJ5J
LKTOYw+9xy1CE5UdBl4t68XUw5mp7+fQiXhQU6SwOpm7a50zJMWGA609mv//Gu3Tr/3AYHFpX7zt
KaQS79v2kcveh/CgNbax/dvbznJKx5R4ZonR0MOxAizk0DtCzwXmffwq8AGdfXbvUzh3zXR7KJic
XlNoIdOcRB1Y+mVOaoEKJgoSDVsdYAV7UuALdF/yD0W1VCIx77QIcggBWIXQhEgW6ftaFHwcCj1a
8+pqMNBrKPcIWqMXVCP1QOxWQJROejMfZkBo/nj1H/AfHmcQ11468W/21f1wg9FaRsZSb5L6MybR
MHTnZITJFJ05+B2DmnvHmG48YzxqplQCCksjVa3kGBqli4g12hYAeusdsz/DIe2zVYNwdNSuW+9t
3Yk+wcAxEeyRvxyVHAlzyncbdIfPqXAAJ/CBbbgVp6Om1Ru4Sh26lYnghIgE3NCnJuk7/itquW3F
KVH4/5hhx1G4O6FoE6R3BeyiEhTlS8FhAFIJewIcEa8996UhQIArPAyKIbbwcB2px6zeB9hMcNA3
GtYGv5PSHxcT+sS68X6DM8ZOWaZMHNqaXe+qzts2XKPIVUh9mlNQB4LL0The5CKQcYmH7RkGvb5c
eItZE+ePUuargSJxo0HpWiIYDttIUqOUo2U5DqQ0WNlgS9kM/50d0fuVvwZR1X3o9uNyMWkO3Xh+
uWQJ/xMXh6nyurgmxNhdNI2XWWfnQlJGkNK1W5mVm39UUTJj87u4nldqJh5F/m6FnEBaBc0Krkhd
DreTcTUk8QpEeFP0cQJnMvqxsRyWZfGPCtbDZfnzf7SnXF7hlWcqbqei4OOKUz2axJmxAZzrlVLA
F+YeC1WKW4pg0StHoLCqGpbmp3F+8W2/AQcY9TWKPwnpXeiVcAYszva+9f2c1QD7+gKiPojV1p71
5RVYobDVi7lXatoOxaJazOWtksYRe1MVEw1kxJrirmvY7lnlw6lHOGOm1DNRHacMSctjHPYMCBUv
ojGPtoBdiOBCtk3NmKveZuIH7v0ec45QGhXNXATtegXIoyCVFy6h9eDHBJZb/1z0FaIJ+esEeqqM
ZOeOO9tLy3hZ5kG/P4AtRQhzK/ws3R9NYdd46H8Xk51jJNA2oz2xo0j/PJVRy3aw9878GK48qjQY
p/9Hx7t+lidsVguiuvkLx7cyTIqK/xIYQVkypZfRhK+BbkM1nla09SF+M2xtA2J3qHpPS8qQRL3W
s1ZP12XMPgzbaQXBhxjlDngLy3Ok96EKfOHLPlVU7NhaBrDMyy5RVeQSQRoq5ll6SozVgNabU99U
FlyaNK3z16KPmicEWbWfabeaRMnEp3QpqSjv6tuc2M6r3IUcLI4hEhVZVEUlQkkTPMUIgANL+/cy
OGyMFNcNnIndtyEJfpQoCHQwjiy5k9AE+aS4c3xKE/C/aOPRQfSFD3F98tJ4gTdiqExh8dpRL2zm
63P1pFO1HXkJSqi7E+XrYcGAJJMCvXprjYpwrWl9f3JfZgG/CnJfmZv6Sbr8Whr9nAYnvL48gJ22
KqGHN/3nMcKUR/in0BrCL0V+avMJWEf0yM00klYnkQaGYqO28WioUZ9k/rClPbMDQTiI0lTn4isT
1yx6p3rDrcCPj90NFZqBcIp2HAbyTiS/e/n4oSp4J046vlHaFS12jpv0E13hscSiMHpxAbgCirm6
eG+mpeJ/t5gVCJSaW2O9NssPGJkoTRXDgaPmbnUO1THcP5KxNd2ntmc/Usb1iwWQxlUnpIEpsvab
G9vhd6xgr8pI7EfoP06qhDteiyiTaPgFXPoXpeQKk2yvS89aGr772k8yBqb07TVBAwZ4KiLCxsTG
DEeU1110rs4Ox3nd8BPY47zqJGf+Swj4tDX6B0+cChIMy0/7lhBbrbje5bxN/yRilPJx3hP9tgTm
P0eX0KhflEkQ3v+/utrbGe7t/iSGMD/jtDZV+4VBHr98wbl+jB1MnODtIapsWyKfhBb99/5KRRD1
drp54aYfM48hHzMk785LX7vCrdBLgBEGg1EFOTC8y1ZwAgP9OpQc1/qGbefvKCZVFtejwDViUbeY
+OlfEnugy/XvhswaN5BvzYSkdEpXoyCC6kO9m8scGK7aFtfJaNm8j6Njq8cUZWSHcxaMy7E9RQu2
6BI2UVEyGz5aRaVpI5canay7TZY5LgtPfCFtKrbWxunXoh9lMPJPEfDWALGLbCfAc2bR7QTxdeyb
wAK2ridYUZhmLYN3g/NWtTIFoI4yl8/nj9nNBoZjbB2PuE/TYiEGgWtdG/buBuSkh7/eqC/m/onI
mjFpTUKXnE8Hv5+p3pI9JHCS/nM0L85G2MJP7gZ9tfjqiCUzGZBnaI0svAGVCfmMRs2SlUh60jVX
0nOtUnzAwOyOJkCDCSw1Wjm/bs8h/fWU9pL8JqQmbhzfbUIY/Uj55qq8xJwvnNteUuGka9xdxrCt
1GU5NJGeMbReAVVvj11rmzJi/7DrRPcMygCi7DPke4qs6HcfEX7nswihaSkeM29LnSIwA6cfdN6V
R8XZzAXT2sjftSle3jWuin6IvsNCaQtV9ChDb3GerlZ/KSK8IwEhi/YjIdYtipgpPR7NLZxBvylK
TE+3oa2cjHL5cPs2G+H97qFtg/D8nyaW7lvYs9+qma+MvEzyrc86ihttBMXXIz7sFwmGmcM8UKKY
jpUoQKyiyO02KdwtjTh49iM3w9fCpRQmFdI2+Mwg58pKdW3faG28SR0e+Ja1Z/AcCl8xkxqErNzL
aO10Tx5X03M+Riflsb/0///qHsP6MGP7cubmk27vaJ8hZw9NrGFNw1bkZiGPRZWIsnV7x2Du98U0
xbM04LJeAc0Eqh8qcoBBi0FTde9NRidATY2iMURtoKIgHOEOzBmKXYNU5tshK4ftd733t5qeJUTC
rT7ZbNqZP95+7Gp6VubuPHoszr+egQAg5B4ErHQdob9vvRl7C19JzS5eV32MuPD47PaFFz64YN50
a2ST+468gwOT6uZffgH22tJt1I3/q9jxaD5zwBZ0k22yffPiXmbuZkNMCyj8Siene7BEwRGCuHFj
J70nqjNfg9KHfVTABzGpKgNmt//C5jn9VLrIj6IKxecdjuobcN3CxXirkO7mLtIYt6x09A5HHyjn
MQ34gh7O2ner8EdJaR4EMUXBOmdAG9s/3ty03kyVMKKGjDLL7uKNYtRpH5aUzrDpTrwyKnT2hs0C
gXeAGX94wixDNcONiyRhJdVtQ6PXV01ckWJamh4qd6/NQD0ypGtKPiagvAB3uMHJnA+/wsCohMhr
R7UKztOLWsUfpbldtRLyEZDwXsuXSWKQb+cgplF+Pup+J1QoiaOjzku1AG8CbbxQufpbGx1Kswaq
nXJLhds5GBx0zSBHa5VlLfxp2Mg6nBBA47M8XxZPX//Agwu2OlwGfxzCb30hKm0qxHZI0LrmL0D4
zEEdijhDlYEkQ1vyQUqZo5lxVMPCcIN9eip2b/bthahFuTQIvnz4vym1NFUbQqtS5wyfOuYru8TR
q+26MfIZ/TsXTniexOBSKc8iC7j0Ya+9VBoQuU/ZMRa8yhompstugPtzmMXiMOr31fiYZoxLnPRX
5AkZ/Djp/cIKW7RbR2F0TZM2nC7JS7+dwcFRkUMPzpbORJwCmn8g/KIWMirJRDKIJwjeuFGUfrR3
NL6H7YdBXTrqrJL15SGR0hza5S3T+1qK+GQ0kLLL0i+XO/Hhoa1M1D3LJ8jQH6WgrHIyjjTyM9/T
ILOiTsuz6calQONJrVuyJRMhopRhYm+TSqzlKUWpEei4LKKSwW7QnyKc+AFlDRTxwDm6AVktiQx1
i3DwbwckgYD0mM+b67F1Zj2qHvJlLGipVhMiO4ncoErgaZMBOk4L1cm9OyUKDbeT1FMNZ7xWz6nL
c9pvqH/ipktNswICR1kZlq4mLBBTuQeMB4wvGbM7EjKEBs61hGrE0jUvPGU9KbxMQQXiiH8jhLPN
Ekr1hFdemx5XaZw1Hks0OVENbnZ3Wo6jRM+MB2COu2DszEARU3TVg/CeYEYR2zheOKPu4XFQJjxG
tgr63xLHdugb/0i4o5rrt/BoOxSYzZifuOaagqDE6GfNnEvy9/MuCvT8gBfpbQ/piYNg/kZWX8Te
ETd1UpHFAk584lCWhpay1KFmqcMDVhamsDvJZJzqAt7SixCN99YObohwc7E6VUVIfl2Aa2pDIpBY
iLagT0N/2KM5TpN49YmkNfRgMcqLqqOt96wKKmaw4GRwtFIlgPgs3x77lM+Hb545wv6s+pcS6tIo
kqeD4omNK/9vgdZ3CTLCKUjjPjraHQk2uFdt2zPjbQ/UhD1PqDPjzhTyCauOlxcxb8nFBCb/NQ3f
6ZbdBBnR3OqqkCMBnO6QsMVlfTmyrc54NwKwoxfyvcZXOzwcsjewZG5oZ/nJV4NowBMKOJ0XvN9f
W814Lvso4drdCiwTSvzf6YsOmjYubBotO8niFpZ0s2DX+fInSuErFqCGwTuUb4eDQwxjksRIcC3d
Yx38q/GGZFkb459wUkL5B3PzF4MSNT6WA+wwpw3IQCTuNKlBLQMNsDEYoN7aBSbpf3vtdS0KxpwI
F5RRW0j7HQwJEbgu7Q5eyDwtwIajAbUHbcKacytVa9kcRoSo+b3qudX/9LB43Cw+Db3EAoMw+Ybj
8+77u0z36XJZ9e2gAKlYxTNE+37o+zsrKH73j9NU2VEtyacB8ZtdMqnYAP4aGtuLikf4pkUPDyg+
wM9ZXC6YtMfBv+yrmvWc7gTz2JW4jmowA/oro05MxAUzU7jOxN0BcjIPvJyVWKlYQlrGaTDR8CS/
UfzBrofd77oLH9S6i8kc+2dk7RpSxIr04EJds6YeUuIne7YJm2Z3FAT4QQti8hM2+WmLGhZ0+ASh
2zOmHHsQ+ZjGOGsXi68OcEbRi3tNkezzne25QA9sdjStEvXPcI26gAJX6PibdkVYP5FDNUc3AvMZ
GosynOv/REfT9MCdmYemGal1+Bh3FQtaie5VW3gK0gP8XCPAZ4j7TIWrk/qqZcnBe79mn6mNDlyU
YwLPGZ0ARKZAO8DB056IjAMnYZ5uDwgG3y11/GA1juNCvlApVnoSIsLarUuXm4VBQBMzY6XyxOGq
tksX/AZ097Ko25VEYwMAyoNXerIpueiyK9gXN37h66L8M8Q8QLm8CRfaPODrEJ463i8q4oSnt1YL
c0UoyPGZSDFz+LP/ykZn+jCARF+w91rQV3WOPWM6NGZxZia/LDlG0Qxu4JoauattNPQhvs5nsZJq
0/OTPWSidDA5Loc4WcniGvFAVCebakanVYO2Mx8Y/6IVkKxJskzCvxxPVZSS0qBpS/0en5jOVSIz
4E41cax1Afb9AQDc88puRg4fQhC18cqZN6ArLPnNva7VnLQdiBoILcFfCSQq6Q0DvVC90cW97DE8
/G7832/7DZdUGrO9hMCgegXCvvQjRRFTSg580VOxoj5zuztyasKkHU9BnmoNemZG9vw4l8R/Oi5x
8VHj5dRlXKdAB5diF+E/EmqSB066yOwwiFRft6pcN5fzUpN4RyKpCctfcztidCRi2ggb/HomegSv
9/oX4uzPlVtMo44UBmfXepyddDf8wfbNr646ssnOLZTddNGt3n6rVYY/J0/QFnWdzS1Bvtvt0RDr
KqzlGPuxmdx+rMTEQ1ld+UCNMr6JGtsN7Q6eA7nE4gwxRbatTApaSX7i54WFinf3hw1ojFaATqUm
T+OpY9WqiiWFv/6Nbi1tIr3H2+rXhdmSR8W0YoddP48lDSCZKgIYTWrkXA7+GM9FkoxVj+U989ej
FbJ8KguiVrxLiYn3AesJWeBRCtHlK8dT5LLWxQEhH9kMlxmLokTLElEQixaAxyyxK13nDZbfmkPS
Au5R19UiwI3IBYbq4E/pbYZ6IYXJyuETBYDmqE8qsjg6bkx3LMXRFhdfwI2UzPjACcEBeBh2EaUA
xNSBETx7kc2NUvMixpblweK9zqOvVmWxiV4WzGsBS2d1g8duz81K5oVgWxrJ35TZEPaIn8V9R3qB
NkAqpx1zcC2rlxPiqUyeOzQrLB61hs8GCW1Bu6ggcYmdXsP8CPo4r2l/4AeFpX4iEqnqoz/6Lhac
EGsSVGn8oyGVoJgC+Ot3loEWZwylt1I1iGtu6u0QtG4oHbw10VX5QSEzwWX40mYuBwK//c4IEdxO
YgqnwN2cVj+0S1mKKtAD43gXctPQSn3ph+JUeEg+xjy1y7W3T0mcFNulOOwUS5Qctam8+ySrQ3V3
MkKrR2T3KRh1i4rdUQJvxa8IRst0UL5AgTgNdxLzQ0wGV2hqH0e7Vd2WMEq+wyBljJ3cIMAt4ogd
We4rUhxBFzPK1TGDkmOil+H0223ZA4vE9UCe3MzEFaBbMHQsUtvbyt6QCatbYZvpZIhrf2ZimwPI
fZ7SoJeymeD4tmXjw7SDn3IRw3I4QBCBJLbvCqGPD7VEDoumNXWP0jufTeQg4nSIvAGORZEfix49
mT9uJCfRAfFF1F+dPlkdVq3TSGfsekZzVgRBfbov/l0trIc5NddgLZqcxG51Xz1C0Ah6FUr8FDTz
Yhukv/iV+NnL5qT3pH4nFt4Exq9QwUWIOngBUJrFdQ9ypmrVk3fjuEGoQom4kvXSC2u85Lle8NnT
zRDi1bWjgQDdAvF6AJsuXOwDp1ReNwMl6q+3LZ6fghItzJwe9Lcw1QFLqHtEckBp+bT27xYbE0wc
79bYQr/iU+/4tzW0Mb1GCBmOScZJqUnbFM7uut0bioLWunbqrmBPh3JDGkrz2ApAH3vRfHVGIqgA
p0RU+wolSsqc8B9vfsaLUwliAgQEAQEeN+whXdHpjZhkyqYPwzNfkpQAESQ+IH28Nixal3ygI7M4
KUCNnCH8rlc3kT/eZ+HpDAnSbKoBDdkeI4+dtXSZCEd8SF0ijn4SKInQI+7Zpn6/vou9p1BPWYxS
xgrJDS4rC0n5mz+Pga5ABs8XiMin8q6cPUZ8YGRD7Z0fOfgsCiDQfxMOBve6YxmgTVhG+OGVRzIZ
5AOCrs9thXQWtwwSd02/aQ48BId3h64q7ppJ8AlV/MbdA3m9PiNByezSThjSmW61SIldBtLfndrY
9NUALkW7SDzlVaTnBerWX/i/vu9emmOa3ZltafbanzwqNkbCbdr496pq05VWpKg+enfZgTtu5TLy
AuW0ZQjrN85tdWIlZLs2T7mb9JqKbnulyOf5tQzfZSa4JtJWVj/i9vXjHopXKYSRXXJ4hYiT4OKs
XpXXXyE+DIhH1Gd6AF4IEXZLxIq0P1N91zM4yR4ZUuGVml0EBOV2TovDklQeG2SUFSZnK4mnhs5h
u0hYdI2v6KPq+mDquAWLhZb+lrPhVq4tygXAq9ErWYusv7nAKPfw5tigBPsPt8VFx+LedZlFidpM
/02HH9xvGWmVzXjVzHwRSE4Lkz8fIcOIlzITcZUboY/kK5CSbGtb83WWiySHxshki7y4vCZrxcoG
p1Q9S/dWpEDm7pBlA8UMI3fX305qPSwVuW4xUfqK4U0BBxtmShrPvrHXwvTsmfD3hOqgiLarmiH9
BgEmpyhWi/Vk9Po93jlI61WRGG9w7XxQBB8GM3k1UBWVjBD7WtCbE/1Ezk0Jc0avU+SrWzSEpi0C
z+VoqHOVOlfu9uq0Ba2VP8FD1s3mYdKKw6A4gd7i4qpZw3PxEPm6lKYGotto96sQn0I76SAMb27v
c0Zg4vgrpn6SF5pgnDNqY2nz1lIFYl0CqWTUrSb0yHwY8OmJAhvLErBCUTfNXH1EEaBRl5U3iyxq
smFMJLmMviZ0a5gFV9z+wq8kDJ8Lvu9h47aP0FVv6wDOIZ0hL3bBrmdeKPj8RyG4yqYsv0ORNpo4
l9g5Dbcce/pSVYbn/BdDv7x0To5mgfe4MjOqC39vI1fL+fw6avOspbCXnRbxkK8/j7E2bT71IuQ5
4busHs9XIx89HvM9W8IjWKF7YDc9wwAzoQVJXKmlIIGwfxmr/MkYvK7kFDZgsTAd7O5aYoihzvPa
/SA4Gpy/zAwLPVQSzK78bylaRLPGqRChd1Zoz/ErOyrNd7mht7G0xSEGg7PYc7RRz+Roq+6T07B3
z4ij3AeGql6D9FxySt97ZNZzjL1Mdp7klk/XhkK6V2Q+vFwPcs8Nrs3oAMyYTJ1YJJIFb/ZgY8uo
cwOhYHpYfa4blk57/+sSwM2tvx1u11nx9XpvkMEi+mKBrW370+1yyyHx+xUFzA+dHadh/prCdtJZ
MfHTPk0wUM5eMaTcvYBMJmQRqgzv6U3OKGovq/T7cDs5LzkO3VzMvLEnZy4KidMLv0UMxq1zsGQy
eGd4Yq2TYpAOGtyca8+jjF7LV2AN7zJdKoXM8hDJIXCEVRXTaxCcY4d/yxOeXV9fhWe/eGXpSoIq
+8xY780A5jYSbdo88csq/OY3yYgLRm5Yo4Z6G+kK0pU1BPA8n2t6JuvqipAHtybiSUN/AvVnLySl
As4/WjbJiVWNECJ52jKkBbFkz4d/up7LLJ2+DYEHwuyvNjyIQKsCNFJwFwmxEFCOGM7PLcOyS/x7
U1+gq2W2MJEPDX61JJP+3yVr2Jysr+gP730wraXTWFBTl57H3mkoOihUrvx5Zm6dGSJmMxuP3vLQ
ARyVqymfJzOwcyIaQmwcGhecZg+L/8b2/h5+TJQ3GcuFa3AKeOIrm9v61LvDZhpHCelHjWXzv0Uu
hGNJob2zAUgjkeMdeit3ZNH/3YeC563czcqmcuEzbxSvVy7TDjNmtDJ364EzfLx06VSArAY0AU08
M2yXVPqd0pTbZBewe5uozXczfCUQIHuT6LAdI2IpXmPE3KQDwtNXZd1IhA++S8pZ6zfuVTHMQ8jF
2hlj0+G2+kbCCylkr2cqBGkCMXmHF31MTD4LEWDD1Bd+O6AexWVlqHahRY0O5EgWTxqE3ifggMsR
PYsmxPPxoD5NbC5tQmyZerFObDJCSti0R3rNoGToq/XSSZeiFCgmg/U7BNhcVPeoNdidA0dfRhfV
S73vuWd3xtGZTgzFBh/F3cByiOqMBlp+GEy0zViQQesE4mpj0mkapZIeoinjGz2gzPOcr6yxNH0n
tg4rHV5bw2i8O8rhRFW7MrhiEmXJyrGet2tY2uv9d505m54DQWW8naLj4p+76k312ncJxmJzzmJa
79+dC8qfx591k1qDFiiIb+c7rOisFofR81/4+Z6YrWok4QA68Z/hHKIbo/NigSQUnkWh+gyv8x4Q
pptRC9UKk7UxRLHu2BdkVK3ruuO7TSsppSgAcKDunYhYGmCYXCci6g8Uuu1iYVsvTC95JCRBFZQV
WlBeKwrajbGUivntPBK/rux2EO6bVqsUNmCKfzI4UtgaIXBl3zYc3qfCGkkNUWV1fKQmdMKwMAtX
5yrGsYEZU2sGYrkqJrkIsVKdeO+e7dVY9traDk4uwTJmWs/tDDKmGQM8D8feLXiTS8X6Z9by2XrQ
5S82VpeKaSzuyZmdxpTygQQr1zxfhONENfNVBbf0eOrBrHjftQehjFhuK4aPtIJO8W7UiTx7coFp
vQbMqf9ke8iQWBzDZTYxdZk5F4CVxvqHtVg31JQK4m4kdZrIwVokl174EMUfwU7dBp5mrYxhaJU5
Zr0Qug9wM4uXNjJGsOTRI0VwNIZv1Xq8wJNj5tLzJRlMqEPQCXQOLHssdz0W36aMMUPMMCDrCPqc
NSKwHnMPoXh44JU47soM74CDUk6opXZhmrSH9UBfVpw5zYq87Lcv2PXlM4hhWgvHxiNjd+eH2pwY
iMFQ3Ss8kycHkHGRgSHg36kWuqneQ0a1q1Py12xg82LTgeB3DwI8a3O9TnzqlWz/0Ug3PwwgaVrF
4sEe/Jonx/fxRhG+AcyDgZaI5NjzfYMRMBaGLf+SS3PVfCQ+bwUydGUftx83kj6q7ZLqAqzQ/BHv
z53QNMIpTVUIVqId37YJw4Mg00LNNfCR+ZwBfkhg+bUv4Ch8p0NZz00sxGVVwJr7mYYsKIyywlc5
ipblKZaLhpRkz7OEuCiiSKiI7J1h5d1DZicgQ/M5nAK1xrTZzuliXwIeT2coumf+X4Um6EMgq3jx
B/+wtVCESfzFyLQ/TOSPm5KYN+TTNjKHlvCkdRdZqnYLVWvmOXn8BXLU5PLbbWkmJJtlkw1kfyA8
/mToqhoQ8CA9QMzxWODSXoqK+9Jd1qI1mFCsYikz+RMjT03/rbJdo95KMcQT5/nGj8AO42Cm7RRD
XeZ43lWq5BXjeALHAn6l6pwPg/X3E+6H6N2Pqh7mkzGxrdIGk7F26A58H0SjOe0I43BF127gW8PO
BvKhn3UzKMt+3mPx4nkpWKH1UqrByFgtEVcYgvpisruxr08aeyDyTQOHxEb2ZUvmfAncx/F8Frr+
mke45ONdm/E6yvuxr6SqJabpSp2ldUnRMi/FbJ8IEtDfYGICbR3bS224pLRIu+soVh8n5pRgCQLA
dq/kQaXi/CmUNzhdxg8DXYqESqvIpnujSMp8vs5Py80razuEL6K0GJ8sqgTuY4DWTE+KYw/sVlb+
58xzG4/R9NhHCIvTkWbqT/tsd3LyhVOq6ZyjWBnt9KhoUT+vbvws3wdqod/xBxVAHrphWMNN2YhN
VXPdRCq7X7NCw7W8aXO00FHa2iomhgGLfEpBCQpMZh/Jmtqt2ArB+XgbTz/rq9SPK/mnc8wUdk8p
YmV7GDV6YWpqvQr+vq4CFa56bo1ws4PPNxXAqbtNyjxvaUjfpwQBaUnoRxNYsG2Ss0ZJY/5K8oAA
9T2ch5X9DUJjXFou8SkoK3kp5V4nFxx8J9+V8nwsOseAPIadn/BsvCCvo4gcrnzwLxvYO/8E5WBw
fttYcTrP8T690lOM9nABQHfO66vkBbZKEnJ+FZfDmqB83ZwBr556gnjyA3p6QfEbr9ILCtozvaJP
z98Qy0iFA1eYd598rU9jWb/yVUVw1I7MrttzYkd1Xf+9MQ6nR0CXRbl0lKscPFAzWMyiiguJQC28
Vk0QS11VwBSfg2dRtHXqMyq0dcotszhUkSLIe25fmdqvAxeQrwvFZQR8bqkT+gE7JlIiV83xXw6s
xzksKt5wlCFDd8EgI3vcuEYSlYDtFi4qlrYADweandZSXfdys1xMLm5wkcgd+FfSfDKoHD8kbxNf
9n0fgaKic/zvtQXTehOqoUGJ+Z7+vBvD7kjUh+xZyAKOE3qfJb4ZaL4ETPblMPF8qUfTQT0Ui7AU
4kx4GjCu+e4/bkkbgnjGUHjnR8uho7KKGQfp0w9E3BlmDFBu21S7z8/q+1FqU7vPv1vy+LpmpBvc
lLB0Tjoo2XuOJC5u9E15Zs2xge5wGtz6twE65IhFDdieOAWJ976x1kgVaVI9Nci/hsuGd7iHRn1S
5dUmBcAcPB12WXsBwoBb3HoQF640uILH6msQDkidvKcEj3Q1EibnNkm2+SoOm7GOL/e5r9uD5VBW
mgDQkdzHfhBhuFuERb3W8jTtxIYQFHbbbMq47Qxoyorxy6pZc4b27jg4uYOtUQWyXHDkdg5jnoFY
8TEiSzGlnGsRBRprbzS97DiTf9MAtFCkLltl9TVDKJs3h7CNoEex784pBvzVvenaKqXlh6K69/3C
QWbeBTyOPjFX60H/QdEVXT3HxvotVpAxwhPqurZjUWWEhhYbktsXdlQGJNEwKxO0lpB27+48BGJ4
1fnr5SI7kmFt4y1HUzPxtS0GJy2iCpdOZWAVHsUBK9SSLCQi7+BYWpi7d3cEYndws3dAUAq6wTfr
YZGP6IHQtScbfrHWuXXP3JJV4Hb6mHFfaVkpjOAup+54nUt9+9afPkRSpuSaUH35yc2MzINx2CBw
kCKGjyfmmkeLCPCnDCxP/LD6PK+IQOUUxCSAYzCDDFMAcYMj+AzULM98XGNDhKrFiWW/9JdQXmsf
BwOc6RXx4210S8ZoHbqtHGhUF/M2hvmHQn+FByJAwl6+Gkh5cYacZZ7Haj5WkR+gpE7wg9tY3ddY
5OaUu7JQvVjEo+SZAZr6bYCF1F5NZCSpIF6dZUaX+0MTxwZVx4/UWQCF4K1ZAF9T9PLfSCk8m6b2
IJod7V1+qXXNSeXRUcpLQvuQew2blk8IvqSFjxK3iXGqWzS+g+Styfhl2PoFuI7CeS37NopLbYtb
BByzWz6h5iMkQwHxeZa4/35IyPLkVxGekVT6N7N2YC9w7G7jOzG/yQPS8kgrpL30ck+MlQTaoMXb
XTmv0N7gHl/+LfOW5kKVu7QTVGvsYKQHUKPedq0C5Z6j8+c9PMphz4g6Lk35tE0EDIdiVtFLNlNB
d8CbXbYEbLNatd1vh/ocBsPi7qBbnl1rn64z3TgrT8Gyn3AkNMRhW0MLGiWhDR8uhg2Hpsb0GUqi
lwrNz1LsE96YQoOPKtSZYw8UVXazPD914rnhgeIf4Vq5ZEQc3JOD8o6pdQyl6aeXFH4B1DH4K28Y
/VgBT2VVY++80pmpbV5nim8S4DPShCavrJpokJAS7oR1GbGZ4cMmuA2xplPNlPs0BdhpWRFQvfXh
zXxTpc6Txze8XrG2RbsUI2o95sNIpVFs/yCFatEF5iyCJz3Vv2r8+46JmfJCiwJ5G1L0yAiz0iW7
PAVUrSMwmE6xMOwLl2qmUaEczzkFazb+CLR6KUkNWs3s2WUBKyqjWvd4gBGE+l5EU0WqHzgLnpnu
qBBXxzgGgww1EB/lzl1qkxJmoLsPPQt5G5zn7S3AjGfT4CnnDeEVl/KeK3T4MLXxDCVSQjKwbV8J
R2zLkskvjgi37AMkXv2yI+qPofmeXNfk20gqd5Qg+uLHaDcljwijcS0zXcmvZMOb4QEnaVRyYDyv
C3LGA/cGeHODrxp0XZRUsrEUq6dqqGD73u3F5epz/TcFWOL7HEuYTxEIXVymclKlJ3BQE2caGJhD
jhCVEiPPWEDQcTsD5yRb4Ai9wfYa9djT9/XzUM1ZHaXXOixcpu/03dyPmBmiPisk9v9pVjUQ/lLq
5pThJU/Lb0hE3o4EMWM4KPrthxTx/boOMcuZ1EptXsdCN17GFn+W45Mb/VrRuC4baQrTrAw5nuLF
Efnfa3N0MJyz4w/rl9tmA291IkghZEDsKIGI3bdm2TBs9LeZFpG9EKBkxUt1a2ct294tbouXZzAj
xHWOECUXuwV6zMUFFUBeKR/m7z/KRefJNIw726bIJd/IXOZYguUyaOg5DNhYbsfaDBmQto7k2K7W
rmDzsjb/LsBWOGnHwosgURwVp8oo5sGHm3CW29YedyVUxlCOzp1Y94ZFeu17LBQqwDYCSHuNk5hm
LvGa740Gm9qsGnxSXQxT/XDIDLjsYJpuJqh1z5/Ge1LwUK2fnvNNNxp9LJW/KnvGG8x9kdxbw5le
0i0GGOaWZz+ywEcwwRxichAuMj9gVdhmaoXXABu2IOUtDGlA2xP0WAcTYZMOTsQ1ZyRL269LRxLC
Q0StUlqN7jq7Jd9c/+toNoaf3ngaRlUCY+M63kM22DFD1rpn10yyQ1nFZmA5ut4Tswnd2nfvPZuz
Jr5JJ/fYw5jzZ2BGIjIqTzpTjbXqFTrJgLWb5axFJf9Zpsl/8h+yLO/698cJ1nFf8JR8yP9WHCis
SPgB78zJga+UVH8OXZrIGQ2eztrDOZ0PSoWYo2R4Bif/XdZxTWLxDzfsfrxSPkk1l+NoeUTq+qIT
oA/S8yyukGLaVGRicwZEDztLA4jQj6O5BwkG95mKMVeVl86bC37/Fz6Zafi2mhrzLhffxIKJeDul
l3hLtvrfnkfHeFTUPGHD/SnhsVlb9LLE3CMj0DSTDywGbYRVkpFxNen9IJFlDc+gMVY6J4R/rU6f
V1nV7btBoCdyd8G1RuDvVrzFoUfL5qqpguf15OBbabFSLpZDOGZ1bnfmE5+n12/2KgQAWNz/8uKY
6gNK8BRgll7FQGaHcZKseVKCsjp1D29iD4gvextPofJwP8Gw4tYHsDKGySzpE8chxF56ZDBUDSlp
9fcidmBKlApkT5j98QkzED9PPPoygTtsvVhpovVqWMLtsGGZWfVB87+eGOcvZpukjbLH2a6j/6Lw
AjabfX+28qek3z1T4Qu+qFB98hdYX2F5/XW4mGFvbug9nWgIKlNk5rUYyPuQfsWsS0xX6C5nO0Da
La06cYkp6NyQaXnRCCjqRFTrYzafJA8MT7+LSW1tacMn+pcgKw5fk+tCkY2yLZVvuW052fkYh8JQ
AlMpoCnDh00VXbDeBxI2e73dbbKfGP+YIdBlcFxLxQvKUvzMmF6aYkS/KjgR1XMzKgLPmsvXviPH
T8Q6xEVw+FEViOe+i9i6nPph4wY30Ab8ZNbC3Vw5SYAmDNJxFWmgI14iHsc9sAGJHMs25ps9waZ4
xhZiAImnSCY8YRszXiJ/rhN5c+dmngluX+fFkKOIgC8VfxgPRzCgOdFD3x0N55CClAaWBhumwmSh
AI1taFGb5tUr/g9y2RsuuBDSzjkTGHKGw6zneosxQmKFhO6nRg8l6kUm5tJVI0JB7YvE0Yxa7A1W
T2NnJZlak3nfb4ReTHzvniop9P/8oS3vAlmqaJIjmQwrTsa5nnWX5xBL6HdfMmd2WSgomYR3FvJU
cPGFC9K+GT+058uLxEakGiQZLKetURRRQ7mx1/oeOW+3y5pyZrmKB2G4u8W5OHgUmGH9yD0+3UGX
IiNBtg+nqLMM5mQ8xEBAyov0keagNSb5EdQuV8YW0svpyco3ytc8RQsPsxqJ0Aed48TK0ddvgWvx
d1Hs0KHPqFj+QBT4QmtViQ9XFEA7GD5MYLpzCA4mlaDFlXRkHexHIbUBT8PCDZVbmlsPcL4Ndtvi
gcxO/vW002ooYJN5od5Ckr1aV9IgjaLRnelWHBKxOvmeDqaBYLmUQBRvFDJDWrw8LHJhOUio8fYy
qHhglPDCrOhfgdJTOkiirpLL2ZlwSNgTsehi6SkH5u0kIWh0j2+Vbhwjfx2830I7ESYyRy7z+l0b
wz4pNfdJ1EO70aYeXqx1oX5DN0JUdWQXhaz8TwSXQx8oEM7s5wdcTvTb2GH22f0L5v2sKhtq8bDI
Ok+ztG8+U7cXWcH5lR1Q/eEsFxd00Z6gQIexGPwiEQR9FReNh/W1MCZs7buXvBiXk5mrXOc7EQpZ
iBabelq40hR8aSUzKbet+mfJaK3zFeFtxH37JDrWoakw6ZfVOJiOFfiNvFLUBtsy+ZTpQUdO4Ys1
GmBcH4iFQy3btRrFL7EVaA7J10aPRqzzfqG/8HmHU0T3JtSgbeoF/V+NXjduKz+aV4f3vpsoKSuE
JpGBJ16+oU9i3cHPr8unzNoygl3INkNTOJNLOdEXufk0JZ0Wuohva7EDa7sSgsjBElAkcZEYs9nS
/YJAILpr81RyOIKYuRSPf88/qdA8u+q7Nr5tKJgB1HcPKXfPXetkBSi4kuUjJYIsGiedw2rrq3+1
0aznczMF60VJmqQXxgVCGF3qK11H/T8eUqQYm5UXI/q0zGU/CkJhLmndwu8o86ulYiQIsBVhzrTg
rMRfn7GTugu2+OKcWmwDa3Tzns6IhwYBE7tZEKruXS2+u7gIRn8vg/d9XtROlMWvw5FYkc2qzuAE
hRMBimlYrNaEHx1H/H9Bifv72RhZB9G/CBYq9ATfySMG7x+6Ja7JlYUOrxiCJrUA9mdMiKaDth4a
k9pC7Ju3L0MBgxnzA592fUqeQE3H6r1qykbsslFCRq7EApE/GfrJgTi2zeDNJ4hcukDGZaRAvZGO
5/5rRHXtwiiDKQTJvljS4dFPJWkFAlpykiMxmsa3AsdGBeUynnwsAhYWFHuiWg7pbd2Ox469hoX6
2onKqt197lW9wBPU3NhBytcoY3Q3c90mKnQSPwhfvPIoKZkp2bYl5fBN5gxFpEWE81EPtGr7x8Yx
cUczDtCd7HzgUNv33Th3E0iFq1Ea470q8Y7ADz4AXXUJAfc2P/YF7SvWLedklr8KFVeLX51gNTxr
UG3UoM1NR1ZJy69spWAe3+NHj0/Cj5R0VCPszVzwqYmxCfGRbr/YmQKI/d1okDqEnzl3up+5Zjeb
8Ei8AXvGvdobgugxXscP1g08wM/Rh/hXfAvZBmTn01ss+3dLeK8W+u7W7BpwTUx2rIBoI8cpJuuO
L0i6ge8S7YybWsipAZqLUhBcpokN7dLosXlD3VcK182VdmnhoR5pAiWOiYU8zTbri1Y93V6kZvre
WKmAovLC4/KgK063FYjA4nld4VWbWTK3aMmx8/hluHVcLIxTPUtFuVLGavFl3p4Mx1HJhRG6TiWQ
3o9FsV+TI3nvZdGDeNXcltuDYQgBHg+WrIYEES0AeyWiM/I6154GHRRSqEF8wxWsI0snDQBylRyK
APAqkos8Whro5z045y1nBdB5FuD6n0PWBuV59Tuln6ty6a3UuRdFxFfjrLGZPCLqUm464CoBH+4e
0H49O4BXjRv8/xJJ2kxbdCEBrz1Lml2SWYpdTtRlYsAlifc3Kl+oWHjP/ZOhZFENmSp2BKOEGdHN
49uQWmw/j49YZSU0a6lmXXvDHwCCqp5wS17qqR67nrpJOH9u2jwcJGiF30xhB9djxxbvNPb3ifKf
gEOe/nuiHdFllfH+/8mzA7GOAozh8DFTopQzRSUurteZ2I0baI9hqYRaRPboLOX+nud9vQKvdQM/
3khvChmSqi8XKEESAoQ1DZ9FYmXdWPk16dRSgyvRdXfL/XF3GXk978V+treO344/Lw+BmTKFqmMs
mCZ+ChvE9tRhKGuFFeNbU143z6bAVnQetmYFr6iXr02tbEZqZ25lb3RgJkMW+tODw9D7lHcCMXYk
fOf6axw4IzsdBJvWcc+LlBt6ZqfmloaDDXTFt3eFgL678lHs+Qx81eFlyHaOUIhbj0tpNHpa3Wm3
yUibRrKUX+4bdy89Gd4msOKhjCH0w+TQx8cGI0059q9LlawrKyHKJjFCMEjogvfinVk0PRfs7byR
9TkBXxLaH+d0dU6XEAMMs8VtPZJnc6ysGs8H1fWrkrxa1fN036UHZrSFzzL59S9a8hiqxLgsAj/V
dbQtvTVCaaQ3obzTQZIw047ETynzBMaPpdfBrCDEI0rk7+Xx/fkb9+HlYC2T77SmBnCmJd+fz/5r
65Mqlm/sMyS3Ng6+HzZVqqaKFJKdgFnzLW+iLDf66GsFEBAt5Mg1uGpOp2i1RH2rczXHb1ohuwi9
noB/W61D5Iqp0X03+Tq9SCb5wP64EPL0BEgEDL5N0kfBGXL73ZxIbZGpMOELAxth2oNAY7LKNoZz
Mt43T7HbSMnzOXg+FJmzw1xwzZQeBD5aNUvDA6ymv11TzLlkddwo5c4gz0fmagmycPBYwRC2kdbU
mTcUH/cB8Iq5sjlucf89x8/wL+5CVgPOxh6Flz8IH6uhogTGGeADJXNBHz5ISErINmUoKlpgmhb2
0xlA6ZGxsWxEE/tQPj3mL/kT4suE27WVLn5SrHF+jFZeeA8GhuAHjWb+qeIU4Qz+c/tkDDv0elqX
hbYfod1jYHni+cLqQUiAdvLv1oJzmHI9bFGrwKCe3M5cHvdT6KrNdpQErkTkusjIP2h7LeL83tOK
9H4qqtTBef58T6t+4vC61+Zs0spksRPSXtBchMQbFvQMFuj3o6E0JAlWghAORAqx/xqim7m9JsIm
4LDyoOh2lmf9QDIS/PLaDKpy3UGIUZ/uesaPZeri9m/qoB+dUWH2hzTZwdTpPTYcElllQ2l1HF54
Q5WxnbYODH1jimHJOqDgsRF6nHMA5s7wlzRWfe2bJ38FUbI5zQbjFRgVEhO3nRPznrmZhM2SJlLS
Bq/MEOuHrOYg1tYAPbgePXuKi92N0TZ/qB9rVT1YoHiX88yNcirZ+rlYAHybLpFazBeVJyVcqpGt
sgSYRJyUoOhQ6FT8WJCRZBa3XVRh/bwQnJiPo2cAGzYGjTjcF+/GtpKg0Kj4nQMmZBOwQn09xL7F
BpsCiHJupfFANdAlaQHl2TeTma+d3211Xc3rmZSd59qkrt+wDsj6B1An5oD9OmgBwpE5GFHI9KDZ
hczGWervH2slIMoQgsUnYcK/5T/JlbLfUTyYvnGxIRdBRCQdmWFAE/1/XcUh8bPG/ZnorK6Umb1v
HISFzPCj3mpsMAYu67q8S5jtnZJkv1bFJjKbUsQOX7TFb1/BAqO66tfZqynbECOMbDRq3PNbnz+1
OsZkOdhrj9REh1W8XEglnarJS28xeZbBB+1ihx3b56P45KNJtlxkx2bu+GknzPMxINYqn6MUU1hQ
XeBHr2z+rRGS0uS8n0kS12YYmcrG+7ZlXXX/Be/1M3CsiAtXhWOBRWyuJz8z+5pzQFmWFRSUuk6v
Zm77Gt5hteFtquRGfUUSeY9E//6MTPf8iQw9K/LXIBxA5A10X29QVCwdfGLPhZ0EuJkjIIQSr29j
o4onYL0qQ/+7Kplv7RNzpLGNuKRUB5aBuhp4fxubCFXSxieo5qLsQaJtkB3Ay9VYFqL2v1D3Zg0I
wvWpoAkRDrql6s6HTuAgHPNfAgLYgmg68A+k5MJLCLsdY938W81k/ES52uS/Ng+FA+rrL7cab/Mn
KMbjF6MkjZ6RC3DU5R+Cd/yD2ALvFyvC4KwXgfXmG5b6QsiBGNt6/txymb24Jt+LVtFQV/UF1yg7
Pp/dwLw3lWksJ4aWnubEWUE3QsUs2KLhr6eDKtzI5FzIdgk9zXMCcGbN1hM7FRthXlwAMUvu75vu
/XgvezYLXjBKGhcAmWMIhkhq9/0oDDMjDrHTb/GhdYymZZXqIG9AY/IqgNbwOR2127kVv3P7eM9s
fQhUocGJL29/kI5PVy4pbeeg4AxM7hKFNR/lVOAqrYNqPFWp5xTZxe8G5SWyIrk2PFeCF3Ov4nsl
9Gt97tbf3LbzMOQaNaLAhf9hGnDTzdm7lXkigDCRB+Hv5eAlN7SNdN/SsQXA5Nak93YIPByE800y
9HB3yl73kAN6ulnGIVSo7ffUFv2LeXknIa4ilPOeH2ju3l+tR4RxWr3ScvJbyJzWxUxjQo9KZwR1
taYOKxZgmPdrsex0Eemtqg2Bgb1I1CAruE0pQQrZYTRznBjz3fLaFPz+ATEPBJm4gYOdFEyYFBw1
m2wLC777X/eJHsx2TKFUzoD43nLie0pKvurvXaiXnxLeVXsQEnqxAx9lB64x9/BpXFnAzwPTtcAf
i+XlXCE/lSPtRgq32w8sY0+2UidOOnqZ8AbRXmJMcgnJmrbp5vUt9haHMkts82vZkIkzhU/DUAxl
GaaoeQ3LdmuYMFXVfgjZ9ihWtWseTJD0FoBLi5NR8ulB4MvqUjO/OayXHcTbcWaBlBUr51KYinIw
EjxxGSuPQjIT7gQ8HUD+IU1Jv5JVMNO4vfD+Y+oXx2C+KU7ldojQ1V943nomusrQf4JyF7/M5gfv
k4o7TIILnjl6lHLqd7R6sVPqO4nBlTYbDmTDmgkpWhSYqgqVdfRrW+OwaZTZBcdLEACER1RHonZn
TxbIFcYdP8jdvrQuIu+bj73yAikQ9sBNj8ZaR+xEjv9ruwEKNO6fmpKfCzdH7dbxX6yFRskejH1J
wN6+a6SyH9IyCB9m1L7mk1lHAlFF2cJtvZXBVgunXtKN31rktFGMURLmztJaZ1ldzTQoytAKCw+k
bp5cOC+4hJBihfaGLLWY1wmxWdQix63QqqEQABMKl86Bfqvb3mGNfSYMFLeQC8yjwklL3GNLSbA2
CjUZ9mZmy0L9hY7JgAD4PhFv3ZWEQynoCrV8+7xHuYNJb24n8ZsdO6j9TFobal7CRgmve5PrSTGb
MXAyzNZpnJTL85kpuD8XuRrvahhrERMNW7tv0IPwlPSX0F8zs9UB0Ye8IsRGB4Gy6QvZDEud59dZ
VhZXUWLbAsndv/Uk1E8bjINX2TJOSfkCNekJoxeiCm580+NGqT/kwLgHSxWbABJKNQM5w8Vu0lif
w85nccimRI+LTv1649hInARxtv0sesVl/WG0Labng+Nk0SYQ2CsQG4BsijwiZUTPqm7ctPd9GU4E
D+da8L8jvkZSPKPHqter0JOkBL8fUWPPNQq1Tb58bufxQvkZMxfVWjjyD1boFb+dyIwReM4UsJ+0
iEY9k6tKH0zgI4BkM9QGSrozeBe3fNj6iqVSoViDXhs7XkeYm6tTcJkU3wovgMRDSYyojq0+fM4s
eDPabf4LQRPkKEeWmMJ0m4snlHLY58LCGRIH1Wx5aqW2Kw430Wy64pW7JrZQXfDwAG/g2EdMVXKP
myg5SS/N39GlSA2mPfHVbmQ3nWbsqjbXSrAZhcOL3FB3nI6yyISpFTiuxalHKvdyJS440eC/rYWY
B8YQpHtScpFUhLencNZkWzMB1HYcB16PsRKiuS6CR3sBdwB3NyUllYNBDmW173eweP5Ro3h06QYK
C+apgLGeJTG+oMf1qUW2SvAWLJqtZfhYjwS2hM+1OadQoCuFFRKbs59rnhd8s86qquFf0+htIyXz
CN06zBrj1BWftBiu3V4n6UlRDKv18VOw25MsO6hxPXG0aT3ollEunX/IM7yJ/B4ggoWugF6kus3G
mpPzXax2UOBcOE2QPxCdGMFoNTdNEh7VNe9Zu9UNjBgIXVJ+pWssw20ulphmh5TYu+9l+F7IxEu0
DZq1szGGQPsKzJSj7z2zsxkp3a1/mqsiI7oliZHpQVN/5dy4wG+0nIXaiaYQcUxqcn/BZam3ytcH
3B1vu04Xh1LzWJ1SFmBJRUvhfWoXKCQ5XpyCA/64qbUT+y4MGdYZSjf+aa1tb+fMA7BA/LpP0zpL
6ZnyJblnr4QEK+6zchjvvnngduQJaJ3m8kVglFAhMZz0V9MbwKPeU+3Dj7kopkqlTFo8/tA3u8+T
cpq4LcNCFbtVi4OnImnAp0f8aE5ivGgIlU9gJzc2BMGO6Vs/LfEYyDyBe3yAVWa1LX3BTuI01VJQ
+NIS0Av7v9zsf9USCBWCoZ/b/PZHSjTGLNjz815zaDf2xIcj7cvcgiiT4SiO1SfpOEKa8L+QnFvB
TOtBzuLzUsnrbLwxIQK0tPHf0fVHR72COX/b+wl+p9VHi+Tsmsf0Mg01d5ieYJXktnp4BamUTZsa
JruN3Wz1uKc7LotWn1dnt8KWomHQ/LFUeHvBNYOEsddoL01GmdLHkx1OvAdz/zctbSwVyXkRqW1T
/IU8vFTqQv2UYfLxGRcO+20a2VI9Q6lr1vL9rhc/2NEL+g2OBWwGJkWkbv+1jKV75FcoOAUw8Iqu
7FoYgJChGJUNDSqips6X6btNKO7ixuJQct6kswoxfLPmLiSKCX0lFbZ2Mo+cdvWBkdXo0OjwX3Hd
M0XXfGCxdtXoZUnuASnHBsOOdk41210TUEMaXF+slU7b0eVpPcsgOkBc/X3EG3YeWKKZYrU6kOpE
2JTCIQC85bWoenlaHn/g0Z6Ff4rkwzX9F0/XaTMq5jWC0+6iO1MMjtf7opxPOOXMme+DXMWDFNeF
TAUP4o33q3JWhATOL3YPwVRBD3V3O0w3mB97B+mGt++wBO1bLWw7nGA3nToqD4WbQsLtjH5esGRl
cZ5W7VBNYCwYQIyfZUdWS5aUGtQ7yC5rP1DP1yNgtyVb/Q8Nv8DyiRMyL78ZmPEL96JoTztQ/iJA
Q++E0DgSyIaNTOTv9/CzF0exMPCDfmmMvd7Bm4bD++RzHT/ub9XRHvi1BzeaCLr1SEdHJRTsY+kG
S3T+/gpX4gJntQU24ZQfcJ/go+PrpCOde5p81vTHzKk+83rVSj81W5bteO0HWhxbYq5gzBtUPjZg
8GhpqRBGA6qhOGNi7pv9LpYmfXuMro+7JFr45Eyu1marr8cq45i7MRTUc+30LgXNmKxcDy7X/J/r
OGYja3WnaLRMgA3Nb6wcODWyrK+ustZj8ClQ3/zUIXU97Hdf6O5eodGPDyhNYci92At3+J5kiwYc
cE++42TQJiTCkpuy6eluvhOj+lXx6ALIxAsZWc8W5hJZbHX4MMWwTWoJwsDdVtwTfcgFTfWT4s29
W9P0zwFTntwiEXCEw1pfvb/wZyNz8P9Ce4VtvP3bA1U4PzL6swX0iWRopN8Ivjjr6ZMmPrhjoR7Z
kThC5OFQhwFh/65QYpAJBqtIiNdVehYInxx1YCGrdetyFTgAqY0iE5h5j3UTn/EbZ7czKhoxPSZr
pwy1prMeIThQmBAkg1EmlCokEvAmv89kBU36dlt2OPeZTPYtPlIZcTUbslfraMIxO7pZ3dONqNf4
JPRk0AoaMEmlBRD364hqTPH7pdIq8VrbOygX3tj4j+B6HNZ+Fi0sJiJ895UMWsjeIM88Ynwcsk7z
+SsH3FwwQcFwoiAT6mnke+RqEzSAnvXKP7wsV8CTs0jRgwO4Djv19Qop+sLwBNYFvo/A3aV7m8Ld
795ww4LTwWLW+EY7V7NZR1ZKQJN2xD5A8yPLPo+aPRQY/jDQayAjRrRtMrCRRd86H9glpTKyvMAX
Za+OgkefCB+dk5JHT1dfWk/WmQjnsq0IrOyVVl3RxsA5GIKcY55MeXGVfNLLwLhBq7Zd8oXhzT1H
S6z/d8X9Dnw2ridkA6f7r49A+WWLjsYeajZKqIHxo1VxxPPs9dln2VfwR7c8GFHqNbz3fftEaXGb
W8z856u71IjEaHTdcmwmHBdf2ZH/70haqb73iJE3SSxtXBSG35cJpXVSrulAM7vXeVMwGFESDJeY
8epf2fSDWFSN2zVF1NJWslzeARMjtMn8QVziIczpQnhEOvUFuqYurkCFJ2VCTMQSRxF6bneXDGuX
wDDYFs34qLyDiypgJEmHmRXofj20ZLYyeRv6I6pD0M37vw8XghcrIHvd6woAFG8EIoqEHJBj7hY0
I2tv4JJxRbYeMqkBJZAtsciUBKpS59uA+PIO6IsAXIYNv1tv/POG2znswlml7/J3lFPmL51Ptztw
V62+dZmUU3vHN1L1K7gMUXNHJvWRZRj0TSmSiA0Ece8uMGczajvA2NWkpjLP0M5amDicTKG0Z89H
coKpQzPJJTMSBTSZc/Rj6eM88g27o9dl8B822xhTIwcW0h+gsYcF/74/Ve9M/T/idsXQ5AHfI+0l
YFJTI1PNOLOnxEQPqdRc/y+W9hdqxuUMESisCuLDkIHMTTlHRSidyWtR7FmqCYrgl1E4lLvH/32q
KqErGhwICz0Ykxb/qtDLMLz31K0mKOD173BQ4AKlbSA6V601Iged1bSmLiWN4JefLoaTwLPfj+o1
Z4f5KjDCtrPLKqE/oigbZ2Y9SGhMEhds3y/Nu1JLCRrd/K5emMaskwWQRegTn2Gk0Yox8DdN79YV
JqrVHwgT1EbX0mRxhYPaBqKYvN9VXDNvaDgLBEeTEuFq7Jy2dLxQbCpZ0l0yNdwmSu9xGHHEWk6E
7X2tiu3Ul3viOM9H8LdCt4bY+B2VJeNMkI3ewbcMyHWNL5jyUoDNEz93d1aTzlDKGQWcYWWZI5Kb
jKMQW0xAgkIGmBPZ/Mta4WqnH4/MG5ZuqJJVGwKIxptg55FFkUjr9+3Te093qKbD/d4jIZmZNde9
aGr0KETHRgZnsdzb0ULnmNBMgBj+WV0FKObawfwZaeHq5+hkZxo4ElxZyMUryJ1tz2V+VEVp4mt1
hZlfs0cUfCQHm3VmmUS2y7WVje8QVKCCmCgnoDpxLuK6ahv9Kg08Dex3LTqfaX0c1lArhi/0mgA4
2Tpy07OYc70koJkeHxIGjlzAytcHagp7XimiTcSoe8ETKBhb+cyQ1bOnwLgSnRP0iOxs0457CQZa
q3qgron9X2L3RJ7iH2JTHjiASeGPR+9wmfj78yTvhTLKMXJ4wvk2XSAkcmfAYXgKtYb00zClaUSs
U7GVKBuIXxZQEGIJsNedcuWKDk22Tll6w3tSgRyqBxjursUfbQHebtOIfpU1pTrLId4ph0D0RRc4
RyDBZONMkoXsndRHati7amOvIaMyoW8yxG+PAmuh0gpGsv9lJj//CxyP99CPX3lU5dmPU4JlQIP5
zC68JtXkxHfE1duDWZkQ8VqNVGJ94pI8KeSRWpAYvxUj7/zDuSPPQufDRmHz5V3o8gxNY5ZGgO3/
w4gM24MxP9Z6ap5A6XrHOtbsuvDVK2SWA3zQyTPKSPQkkEfBPeUH+9+XCzINx9+lx3IIjJUo1J0f
u9GZus63HiyPtMKCk8j12IiakWHfz8Lqw8N3wIpIEdZWZ2Kq7mEKSKPOAzOQjvV5+Us2Eot3ZVTC
0c3HvmZlueYu5nL4HNdYnh9dWwaGVAmGs+bqT3Mfz0SImDNNZg7ZVZilaAfK4pj1KTRg3fpJvL2N
3hlJonSpgqTB2apAnup0yXiEb5vhfyw+6qiUSHqeNdmU7myrwWWvzVU3p52Fu3esXuQKYrcQz8Ir
C9QM/zHNfsvTZTgoko0bzrK1lD2AwOOOfi2djtt61ez69vC3AAAE82SJ8x8TbHxoDp/dKESdTMqP
B7RvgvB5hqZVuFQ0LKuaoCogCY9B0GgSmjiaFEAaFqND0Le3oC6F9KhsUL96IqV7YgpSc9jwqtvU
Dgp0f2KMeue34ZKyA+b/5zrg6e4FvKrmFKnJe51OGMFqon3eyk8tZTnR99WtLQcxjf1+j3jSTxe0
73Q/JVjYMTCWdd9EzQ0uVQM0IuJCyPL1kT6UOXxaCCNHPIFYvVxvLqM8DJs2FDmldB300GnNR5b5
UTQ2n96Fy9bdPPAXX2KWSWbaGiGGYc4LhKeOE4L/LNmJIQfMq1cKPslyHmgxIxbylqj9XGspZ3zf
IxlNivDEhQBfVjDD5tLchHV+qmuvdiEitU8tcw8zrg3ee3z6SMkIhRnUMFKW4HG65+V8tyifdlz5
IzpV0L0vvGKWjmMBRGBImsSChYZoYM7myv9cxh2jJXyBw4GJ65NKDKP3dqdgCrhjPiGdi37io5dp
sTxFPRCdY/oHepLjamKPXA3U2HuHd46wmGwvk53aPmrXf2DFJiJPcUqrlsHP7Fxjd8o4d/por2U8
wx9/1tYci1kRU10IBWJcm796PO3J2T3GVISPHsvHXY6zhpQXWAVCeEPl+2xAw+JD7m23v65qnpE2
sy1h6iE0HrFvYddJLGWde6zBYN3MUWC/IjzpSX0v4vQqsuq7C0Pc9jhtzST7IQQdRr+6NMDUSrus
Bmkqdw27N32G7U2D+luANhj2BDpV7lpxHeBP/wsWt9ih4LgGIyG3Cc4HuvuEmfzI3Pf9rWiLkWLA
FbrezCPn0+MhsD0o1QOvOSH6KuFUvwwpO8GeLv6dIi4aXW1yjMzmnV6eJshhGYi/3xxNeXQSKqA5
GowaqfgKXXxCST++4r4nWGvdvA7J9SeS3/wxEIoL/DPF/oZjQVKwOy9VF3FvZembwjNbgujg+lUW
RUlCGAMPbQgosC+7oYoYhuP8o3VfILENjCvOEzQlD5JgiPZNkZtOvB+5IzaH4Spxdby7LE8HXnjy
mSDoMtcPBj5UrlQ6xqc2FjiSVG69PE3Q92cNZ6KkJ977tQ2dehM+B/wNwyLU7qtP37wXonKG7HQz
DPc/tAhx7RVEvOm7d8//hlEte+6By/hUvXLTsPGdt2oFjjN8LpEa7LFSdpQ3cdd+E6dl1I3ZvgSR
k0wmxg71+anPZhPfX4P8q7CqP9/u1+TUPGY4frOICuuGIkgTdpjHf/J1YBHzqvQXnvGCuHoiwoc1
cpmVWVkw82UJWCJFaTzhfQyuU02ZR9jfSQV2ve7Vj4YaWKOWMJwW4aNBhoO2o6VT3SA8jmqywgiJ
9idtU6XN0EFPXnvui9XczMsCxvngS3h0pW6DFGHWVJoSt9sUSljzX0QVSW3rJrd6xOSL0/M6wUhv
OItMDiG1Bei4FmlwCbSPQUCvB4Hv/aKVC2B/TJqwAarXXfWqRCQfphMPniPLVZFdk9jKkEw6vm1F
ze5JnBKL6ncVgw9CKdLF3W1znkby+IUQRgUcl3QnkLmMI5vZjF33u/cr//cyE4Aoi2lbjSl3DRNT
D/YN1c5b05/20iw+khVHatP61qQXI3VdzfZeK5O/Xn5VIOihhuosCwiGB6mbLt3lNQnzK4bex62b
RJYyUBr3jVOpd4/SttjQgKAQ9cbAueELTzv0a/bH55x2sSrwK9gTdaFOpmYhXrKSyKqrRhHRHiBq
NI23jIPVcYPnOCw5yXCW9ikOeHaQcaETg7CvDmdekyp3FR9QNAKNMOrMECGSPxAerorfAC3ItOXT
4nvUQEc8mAlZkRjgNSzGChp4lEpNIpBkg225QOrBa7HUrwTktX9jJ2nKkAEf9FNL4s3nx8bGJ7Hu
NDwuzqTG4OU6LUXCAeqb4phGagVpmEawUdkYXoNs3nnyc74vyWVatQu5NTduGsj4aBr9sddy37v/
Zq/JhpBb158wqz4WUPCzGHAK7ykipmj6nriM5PlSLxbVUurcoM+yCzigRlSMesifXCYuthAJigNK
IhA6MD6FmfwqKIVJN1+5KX9gCfJz+/6XffA8iDdHsCmNS97MV0j8H7ye7LDi6WbB/rs3nMkJXmre
MvFXtaTcLUi08/G2KDSJXXOtXI6Z/7xsdZ30iXCi9cnX6HOizgyGfZX8pjEHb5PBRM8nhuiPbuy+
ALst+Xl9HTgJAR266+dvpQkvezHjj5/UZcyBZUBuUwjTb7sz9qnafXHOMI9H9ranuMCnm+eNhw6m
aARL5k7kBB+VtZ7NlYU5NNOyNfMhr38NgEcpEitbys8rwQmHLLCchItnaG0JmZvG/MEtWfsIxIt3
RLS+oTmO30H3yLUb6AMlgrI0dACbnq79Ic8IbVJimHoNE0zrngoNmIaxVWwcu1Ct1TnVHbnqckWx
RqA9gaFoq4ZcA91Me+hZivmD373peSnTHr8jHg6mEfvWvMqWIlcb1flKC12YSmLCJwhkQZ55Zpne
Sbuf7boKKau5n0OQ8AvDK6IOrdpSpBVx4f7z8Re1OJMXUeIg865TKk1HraveeB3S8eNqN30KrwZg
+5na7YH/izeOTsWkO2OapvItX0d00n0j6+1GlKYkePbMn9JMwNWvirxLQrLZ96BjZf+Jg3PXVNIN
OD2szbBXeYOCfUWH6mBReUdSHKVRmba/iHlOsef7wfGQ0jOH/fJPHEul3P8PEW4J49anbcHrGC4H
NC53l4Dnwzy8jwtbDb2xa1GG1hM07o3Iter+n1ysjJ54023KaWnX2lMOJnfVzKFC4L/c/LHQrdGe
A8NFFXyr42UmY699UOEG4DvmiklffJv97zvMlC8FB0nFXCSnd+axxgwAAhOvhQSNWMb6tOt805cE
r5h1uVZ+Gzrk218PHvmzt1IUYTpUcnGusMZ1rTSRT4P1Tg+x7gyDw2FP5WpF8SSxJi8CEBNxMEOd
Knf7jTgR1KVKal7E3P31fu0JlcdDNnkq+dA3mRAFJ2R0OCvNVusukXyPnPKfY4jtBjcyMkwjM/20
oYw2XLT+x+0Ap2LN/2K6bnWMhXOvBE5b8rM/lalmenOqg6QQ7J8KZfFFDPwAHY2v9zpZf9MK5KW+
QroPmly01DqKJdKg4UDhN3iN5A5pBs7i2OZpcDCewWxoVk+qmHj5AOZc2nCVd9+aCB3mHccjRF6F
fxl1WzToKo84CSxggzZEkhsOJ+6b2cU0FUS0BQCUWMRxJYMZr8CwuHE8ljv3IaKkv3/0LR+8dmWD
KNhF2+0HUW4KtT0+eTJqOgooWmrnJtRNmxG2dHj/scYFFzTU2GElWn3UrsKklekmLdd0VV4fUo9A
c4XgRdMpSuL+DgDTULbqiBSMZ/i2YzGxzsuNjWS2JkvUMaH8yb01wxGFnHJPBGFr4yD9z29yxEZM
og5gplGJ5gIYqgq7MviR+AcTfeO+BOom4Vfubx7IETyuwKEYkmZvS6gC+1D95z8aeoi3N442Ektg
INfedyLc51P+3bglQymjHKHtdrZ0NNEM2zuuxdAqapAXim24dtuZKRy6bplLXCvWecfPvg/U4w86
IRYsDJF3dBNXPNZYXVGU95+YcDhhDg4FdSgLPlzYXs9N7nYKJ70nDN0eM/fhnpQSFMLodrO4CGbX
blNgNfNWH0mFgg720/c0oMvMRByqsMi/hfWc7S3q6ySVxvUHaZWJLifcl3nPUgHdacEIPPXspAJu
Q9IkRqpER77pzVcGpgvJGSfYfBM/LooYebKb07EvMyx0VJ/BYJ82GQCfOhM+ZA2rEUINn9stZo9J
MyEdIE9w3j8V2NM6clGJNdDidSzbn35ojpt7MPl6+VmrLTmLvphRqzeVap5Gvuv24XBTJBnPvRAv
uKQ/yRWfFo/on1LdTq17q3wt0799LzwVBFkjEhbD2Ewrt+pIKATIH7xn0Bygh/FkdTcR7VZAlk/6
WbM+agxFPFiWeEpaAJispNJ2xX8pZsVE6mLZXiH4Ow07KSNg+pS6BnF+gpBlZTpH+BhpRXP4zmur
5VctlwK1WWekOB6KOW4Hl/bCDfQKuJJadhTYzXJmcjQ422hoVlwge4/gGPHgvNfr3q2IJF04/Gch
FkBmZGrHXMe4W/SPeZjV5u7NBvjP9wZY8pjZwVrrAcpjk+JN+vMu0DDL35xdwhdZ/q2qBxPqfmrW
GsPLBMIbT0P9yGAXf0S6n/xaQcXejEK3KMv9DnXxA8EdjuKJuDSG3f/KAXjsu/V4D24vl7TmQvrK
IfSSIInDF8nJEUNlbwbWii6YtimOJ1OHJ34AsQNaWMyhSGGIiD0/Cu04dCIDqjHGnpEpNcHWHQwl
59Lhx9+JPq/8JaJ8c4U6+j9ljn3bRzfve8tbEhC7cOnHLIwHM+nwah3Yez0Tt+uvxJ1/jMs6ttDZ
kpoOeDy7J3dba1A4YCEy0h39AHx6o/wVw9iq3XgvZqboJzc6/l8S7ypD4xsHGuZ/WHFCiP9uEf6K
gpYxq5dMhfrOZWyHknzofxfBb1GYbORR6g9coQ/HwHdFjhbdO9uWaf3HgsAnXAZk6n82SUy7oRi9
pjq3GJ57LW/9EIYiamjQMAEvPrZF2DKq6lklJrUOcpK6CfO0SR4mQM/HJRel8TMh/+T/khKBKgr/
QWWnBEImQzXzo68C9gXFYvR1s5zJ3IOZ18sVpukagBZR5tZ3+8fCnkPTht8aWRPsqM5zHLOstopH
QcHiyiFqMqiH+/qX9XbbVR/C696ZRylP8M00BlUvDaIaJIQ7mXwRJ+Du7oTILqf74tHY2vihtw6s
paQz558JNCffurPK/DEn9ozlNMxmXDg5B/cWDfnLU39O0pSEvFqg5yYQEX8+8z8OAR5Z/jvmmNpd
cEygKfwhlJSbh7HnKmBW1rXpsyaavJpxsMFuy4o6cweUqQgKyVZl97SKV4WUeY8cv5OYbVyzal15
2wWneBOIjGIJXxRg5LRcCkwB8rE6CGM5+OAJSNogWOzGKMaZSneccO7OMq1DEqaS3vVsxuFCPpMU
1a8c3kx0HFWDScRusbCl3nX6INOcizuVWr91gNI1PFq5QVr2nbUf3b9R1M2Pgc7uzrnrbo0Iq7gA
n7FSsQanNQKiGPFyU0smmI5mssFncUa1yHUEc28Q+13XmN91l3iT0isPdi/5LSiTLCsCrQD4y5M6
sLv40uYv581EVza1r+rckpTQJzGdtQ6i0kw8nXlu0y+pMbUIWvJigW0kljDNbcJi2m21/wZOcVJi
G6GgRRiz2G05l/KjD9lq/FeA0FZa2W/OjCOBuONzSVu0zgpQBJKYFQHGiFa+D7stjVFHYY+2IBzJ
tL7mQFefmr+ukCvxAmbl3kFFSmVytQDToHsXPBrDrn6GX6ocMYvRhv9duKuxLm+kC9tdxo1dPHwY
nruJY7nsoZLND+TKwKsWA3mts1UW9mQXMATr5T6F54SzIHfS8POEk6YEmAcsPRcxaWyXqQwGbNQc
Zk0ml7UBzcLpuAYR7hKDyxHUtvsmc6uiOuZZDdwE8dlaFtZr2WHJMY+NaIwaZ6Gudn4nWOUDGPUo
yrEdLvKMZPaO4p3Sf6vla6AupioW7M9p9DSDQnQUYjGL0glTJk+kmaesNwN6IAJHv/vE/eylbsQB
2JVILkmyfH+hZWq5m9am1aleIJYwYOQh4YgwZ08nHSzgW/O5ReEr1WD9B3+sZEFr8yQEGRXOEAdy
XuqDhkcWq279/pGI3ancjJpPRJPBqRVPFhQPbgq39nyfGnRgF4aewud5nhV84wGnIGTwAbmdXHQd
PzFF6vXAXwOzHy6DLx+9odNKcv/Yls9pWIJ+ssTDVa8WbP//OR8W5KPMWL80KnN5MHaMYbi4rX/J
cTnY91z/ibh0FKxQvsPRpQLRBfeWtezFpVIdsC1H1AE+Kk631gjbbrI/30GV7NYbRoWjWzkFbK8h
Z1xyWw88FKQUmboifmBEVu6RGJwlponC+pWVRAEytXerArqo450J2NCcOvUfNYaO9nm4/DCBZMSk
fIfwZucZJ2yBREMdz+THH22X43jbIgyp1eZUxCrtFTbpEuo8G8/xb+B6Rtc2o3D/3QzwqLAyXKap
LM/P1HIHmeutZJLo3pZMIdo7mm2bSNM2VgAk7Q2AVF29w30d9+XzB7bfCwydB7Jx1sSSqcTTfNq3
zmr3vK6i0KOn0P6r07wDZm3xzvXY6u4q58WDZ2daYeawXT3yP6C+q5njcURIIF0QhYWFSMo8XMeE
RX8iVUfT6HDgt7KLCMo6L43/rIkUfrHt+UwxsRThgK94IJ5agFy/OGvRxeaOHs4ir0kp1qc5cLUE
hiVN4O10VL9mfI5m8vwaHwX0wdKqPXvgm93awmFxLGMDaNF6sUjKVRevpKqwP3x1uDRXYDpIvF8H
jG3tTNulnJRBklYJWqtBHn5EfcHxaJAaSzRpVl3xKxzhBDuVoSBTTs1j0FfLtFCyTL/PXsTwIVsX
ObgadFd/6q+6ygE4JY5US6y3KLVZOtNvRMVMwRm2rOUaT9uU7peofTzUHV7gWXojekP+lbUg8Nw5
VeKiAxHEzGFKiqXg3Jl96O7sHrNl/CfYdQCJrkJ02phIyrKI/t82fg0JKsXYrt5byhoKp8VQzS3i
8qUOPEKEY30sXkGOK5SBec1+0rkpOjdpznYMkaf+nlSSf0pEhQP3VA2v6IydY6+JaDzdcUTrxaZr
SwKi23tHPuHg4xMKFZZLHKPNPXmI3hLGoS4nzvrA2RxNkxASkhFHmIQwB78rVJMY5RTzxpaaOzxY
k0muRY3rRzKe4P8MJdjT1DfTHWQA4eUuhDKmW5sCmPqW4WLFesMulJgMoDvrSH1EXXQ6695VBccj
eVKn22WKkHnPdOKQ95ik2sAcpIQOBb1Xydx8QPogb87S4XbXLg857ptHeTZbwo6TvWkiXK6NnX8w
uEzbyaJuwkyCPLXgivot+M/1CkrYDyhFad1L2aAi9RpTRhUoU8gX4YjBTHTx/rYF7ZG3WdFHLLGq
ZOMdo4cjpej+TQv3bvUSa1dHZTab19qovU87a87tlXMAPHTWz4tjsJcQDrMUzUNFHrTEbG7byXwL
SGj2ot9PtyoGuFOxrMWSFojFBRXhitPOURHfJ/tK/fk8CklQs6fIC9AmDxEN1rpDTZcy1mUko6Ws
TdUGR50X5xAnprg6uhsK8cztm+J/quJNaiNI8qsHwZDQFL+1CanxelU7EFE1lstu3b/6pNoeye4X
FRPC9VTvphs152thuigK3j6K4RcjsQLXu4QncOI/PG12hzf/LwQSHiP1nBRXHe7ivsIR5YMJuFVD
KX4g61I9Se/i3gR0swqeEvD/Ey0Khji0298aWAwEAshfXRNCYZlpCCpMFnt01vpXqXOVjlwrPWJn
pCvpHfjJHta4LFD/7Sn0s/cD8vBUJMJ8GK4zdWwtuNXDLk651jCuajgl0YWKcwf9rmMvbG0AqoPN
pnvVEgFeMsjBZWbiFP5iL2QhqNTLcsWW1USikEN3LW+d/vfmqyD+yJF9zaHq9vw2O1zrE6KNK143
nHkoQoZ4AtbRl4oEMuzbewseuXqZeKaeCcV0FJhd1+xwMmtWkBfW4V1UnYef9tixB1m0dLgf8+kP
AtvPnmXIpOA/UwfzzlPleVObMdEhE76DXKva+8mrwW7PJ6QCVMWYGyHc6h/pp2mDlU+9X7VdBeFD
MCaQADjXp7znZtLi4sKXqtquZbsb52VO9nD9Lb8tlLGNeO1lJ0HbXVDdyPexdMKJXpAq2ZQYuwEv
fa72386uxhT9SE5Sd0EGHlSQ6wGQMng67D6LrTY11DKV6cQ58c5KvFfQwadOEFCFTOGbmgxWuQ8l
A+zo+O+6QIGRmcfMdbvZVm92nKaFrLtwMZxcYFxhhVX/eSb6ArvRovwvBlekO6lGL14n21W8feKQ
5mEk8US6ZgL+V7W2yPBs0E8GDCgArqz/nbAJSH/v7kmVWQ9RhHX0zOqxYlYoqvXZeLjQHL4vh7vY
+HezWx8qX9euerzwSqEku7lmq4yc3iN0cG6A6dwremehB5IQrpebq+NuxGQALxEJV5Ccg+RWaVYn
Pyat4IkprB5fZK37OItSecdxy1HcUtzw8gtxTJ7Iy9bZOQp3Ru8VjAqHBMTK6lYiAge4IkGAmB0t
dad8D3WYUdaIwI8R6kNrCCyeY6JWOqZyS1TRyuDhwYASuKn4kvjmd08qd77SQ6BEr9MRlQWUVKJF
5UCsFJZaTigaGTPqELuzlgIzOyTK7ZSYfrypl6l6PG0xet9HO6y32DEvuKWMg92ZEVN0s5+/jJSl
f0S0q015rapAcxhmLdPpt9GXZRQMMQl6U+MB0rkeEPZOO2M8eaV8uryM1aoOmbSIWqEEbOWMt5tZ
xfqeG8Ed+frMYAnOgpDpcYniR2tshPmSF/b14fv1GD6jIC+8M1c4OYlwbG6k96hWOrzC50zImjJr
zPrV+W8yFNSEKrpOGJ5/NYzrFuTI2575BJLaWcagSrsCPaF1+/6wiFwyjVbAl6LNrYQz2g6IpxJ9
IiJOrsIubEt4fECV42P2dX7n9vSDtmdXnIVw/fj3gjpsflMX154WfmqUYXa61pW3eE871u4kBUou
6O6iChAavzef4EIm9hVHuthUY9XxtvoAnfjmNsts6roy3ejY8hFcMMr+Gv2BwHSfR25bhBFmIENJ
a/5Hs3NDcVmL1yFIYE92FFwB/qMHQgfdPgOOm+jZw0GCJ8WJo7J/nfAXHs0grK3G6j+2jA1PLBR+
J6li7eHLJkLQQe9UJHYB56M1V6hlavZ9pineMRttuLe23FlIYMRho617qPBjVqK8GC47EKkVBlUk
S0e+vTcFH8CA4XoKNtbgAD7moxgHAaQFW/GDBN8wrvxCyVyxbqIm4ePAqMEjNHUmFZ+Il1Pzp33F
8KqB2Zg0Wv3i9ytCagAideUbzcE7FqRZ8MB+OLuTDXzsQrg7F1GngTrBxhSR8hPzTqeVLZn+3jsx
hw9d+cq9sD1kkNVvu/6mB+HplTrGGvV/VRdmRlrkoiuE3GsrcJ5Lxjgxkwp0V9xnEi6aTXblrQXK
MM5X9gMgTGiV0tLr1GLoQcxcLIlOxT5dGIF/OKU4L8X1jb2X4NQtQTvZ4cm6FyDluh5Us3Ncyz2Y
yirRKJzsVo0RfomYGuztGVn1T+qFCDfwb5v6+uOy7uGSzcVk0zIfhEvDbxDeOj/aWpXZelBKPoHM
YdSFyenh5IewtuIaQRD/ezc5xOlojx4eu2mhJ9aPsfjd5uIrpFnGx0Pw118Tb41WIhD0Ic2jEYWf
8/QaegZUrYXOliJKQ+4HWSg7H4sFm8RIY90L7gwRDzEFkOfapiAfoSnCh4VrodACdgL7TlnJYjfL
tcrdjp4Rh1YJzc+u6kOCZCEGPvUUDHzZMBB7LZr2Hg5iayVZfy1s3p8UehYW8jbAdNdgoh8e4lWt
FKf+YBiotc8qSTqBdFabq3TamhgRni/LrzCpx0umQy41vKEAF0JQfhKnegYzyDyTf+qDHxzQbd6s
P+t4upz+VJK4Rc11d+/UqKVw0IHYDklbo5F1CRYwFsUyuh51UJ+JmMbPjBSpbBXxgjaWG5gR5KWv
N3T+qXfvbufyvZXHtg2vMOvFry3LiiCBa/udbjegU2LoeeONoNWLznpc1jrF5MnMLju+lKRELGfQ
fRZom1814n3mGHUMZgiTPhXKT3D+Xupgar/uzKbyX+rVFsNwqDatH9AxhfJwTrxncG3xTrvM9L8h
RudE2BVuzmsumb3m2Pxg6FrISPMa4jkkBWhR7wxNCWDT568sVmgHECuUMDX0BdZ61oih0BD0LBjd
9Xd51nr9KRERe3G+RWI/YKM4tjXd3+p/tawibIajiNwBL9yvvneLebdyuupJQmnUmmXiBW4Y3nt9
/iA6CHpHMw1GMQErCJ2KQunzyZo9bKdSaV5qB65ST1bwYQ5D2sJmnmWfx+/gxx3yOBnDQ2Js6FFW
NmwsWhnN6UF9PetGD2pOO5taqyLxugOUTHCSdb+hjl6GrVBBR6QWSBN0sBTgkHhfAPXfav5r7g25
nyUotMq5fyx1OlkEg9h1zHgiO6xuvFqQGAZAg79Cfaxc74s6wZ10mowq3MNiU7d1WSiSy/4gsTH5
aXrPzh9O8md3EWzZtOLQmGR8KD3SdrbrLPWpX8tVMew1ZJyoeuGnRftTaU3ekD1t/fCkR3plij9F
iIYjW2B5mrG5vAlbP/Lu9Ck18NTmF/QmSEHjXe37mIivqZp8fXUQx0FgIcdr56818E55W79kzrlX
AiyEeHZ4h8bZompmZn+Wo4MBIJPuPF2H2+MEwgb0SECsGlCLm5qoxA9RZBUhdbLI9FgC0Ux1YeiV
/XoQLJ5uK5lQv7OJYnqd1wcs6lsqt9Xn6k8ZcoJdwspgq8Z3mh06tPhgzuqWWMXqdaPzWOnp0Dm7
7wchY7+2UuKCBdBMAd5gSBt9Yeilf7bs7urNTx2sDuzlTMruC/3S6DJZnmGPOzRXsf2Il+7UaOOI
dpTTai1e7sLqcfirAsAr1dCi1thOWOLagY1ssGus9hB8wihkDpUfKyvW8+ErBjpc6I6pHmJaSf+c
6/nCZJa/T2dQ9uemZ1aXUiRdQf+ft0IcbIYIiDdy+QXq9HcUpFV4JBOSgvdiNH05NxMG2llzZWXu
U0FS1oyP3myV58Peq3XIhRkzBXqoFjMxBp4Uqoy2KhTG7Ls5ceGtP3gHJh8Zbx/2/eXRth0z2U6Y
rJ0ZPHq+jQkZnx0TgChKyfLpSTnxVPzVMnpRf0faniaOFkH3gkjWi0c3wpEV9OPKi6kBeuz/HelV
5K5iaUhLpfZCFAJ8NFfIqWcMDI8d0AP04CDy7cI7Po26GIdygExhbmSvxn/jJ01dhZ8VfjT0SrJB
ti0DNMUYY/GraWBUIpX4VyB++wxqdIOFDk8SS/qoZBJois6LUV5rBhyezsuN30LUD4hBNESs3PJY
c8VQ2OYEZE/Bpj2ptfp4o5MlFL6nMjl5+FYpkOQKW5H2sDLjqYtZIIQErDKmGnQWuCz76wrCq3W6
W9wsJilSZy+AScUdQCSSVZ1n4C9J9cs6LypVQLT1lekumbvJe/Z2iaCESNe4P9fMNhLDsLv7AtOB
p+F52iWWPc/PuNOn8V2E8FK4VgZQg/dro4f7Ttzx1C1mO/00+6eYEHMdMYK2ko/kZlGS5yzXD1xL
QII5K6iiVw9QejhU2IAZ02WxW/rhJ01Xa/pGStblZ5ZkpmdircYV/FOEj1VgqSf4u20Jc4F+yCvH
KoidZLNFncgwYgJpjGJuBjxnYDeKWyTuc2OaadHNYuxAaAWZMM5gAYp+X2ER+pE/QKLPGckPXYiI
HwSJOyi1Rtx8DfCsIl2sXhVngjTGbIfZM+ZueyT8PGDSOATClwpro4oiktRIGB9SVT/TI2BLHw6C
/JWhulZVH6W4YB3GyVfMVQknB8zGWTMqqY1fHVCUqSwJVISp70Xm5Mv5q3y8YIuebaj4rv/TAu+I
qy3Fy9HoOSO6GPOiehutbLDIU27autzjGYvTmHbxJDSKZWyjae4DfWtC5vtPgiFne2XmgLmVcSXX
vbroa0h3FIqKsclcbaDTMh9dqv3WLZK+wfBN/8VVQkP8ie/BnDvJn/jbMF5jit57WpAURbNfWygO
DjqhRkJWjtEseVloa2NLk16SYi8ryoRQvOi7cSRHoRvWFsJdAsL5zpccJ8QC8Y0KFy748dot+M+G
sAuse7Kyp8Ma8rwnYQJjJx8SFWF4LRmO4R3eefT04VOhOcJuU+Op7Gn5B98CRGgCGShnkLwd9kP2
CI3d0rPQRremvZ5ughad+KOxkKJCCVylx25FiH0vnH5SwQfY1EyXbVlpIG78QmJCmCknHd5WQi4N
ZI/MynRqTK5BXetNsEQeBk2guxb+z7QnmMdy7hPyZGRKp3gKMQQc+SbUSZsQxRni1PF++FlUv4Th
xM5zGvqiAjz2FnWAA2KxzrhnNDwho/22sqLZdxQbE4Y384LZKw5m4WHi5IcO8t9D0Q8G+OczWMTu
qrDotsPYWa6JIycDXs6lF6SFNYM2N4RFMDJZd8lEukzE7JQEBlBaWruQkrnGkdsnJUkDY/9G5jrq
e8+MpQOULAh07DJC4DlzvQhHqpTPWphCcIpm8L65rmfEDnh5QF5uecxbLBfc6iSpjyhV6xwPZPfs
nKD01eMHltqMFPBI2qOVV8O2Zn9xgk2/BC6TFmL3oHgLPYtynzt6x3Yginn9k1zpEIcnhn83ideQ
brfwTPDBXLK+Ls52D3NthPvO6G4azpnDMGsWWY4VDraFLukj2t0ysCXL8K8e7rS3cAbWFBoA7eak
Ul/jUcJ58eZ+vGKiMNbXx+VZpY8C38ohrmrYBA6Qyx+VAmtd8BHRMXVElXSXUtnQAC4k3YGoioZ4
B6tsI8HuvxU5p5q8lu6PICDpmWvdBadUKbZ/xme/HbKNFaxhSNQv/+1nzXAe/ArI0/RqQUpz+CrA
PxI7WBtXS2oA7f95B52449HNDOe9EKRMjnI/Ph4sV3Cs+8ViVlevMi+0OON1zZ+OlS+Ho7FIrdr6
tvZrnWXL6klZBI/6cOam1GAzKsfdgTtdfEpPcae8LUdmmCkyp1Wgeadk/6DinUOZeNHBsrjOlLC7
1uG2/WWIDRgaEPw8qEPuIGsuxk0liCbPJsySKNyRDM6vM6vtC0G9CPgRCuYE0Je0gMrjP+XVBQmb
CwBSNPsnVm5KO7R5I7rvxtRxkRVgsagf+Ju4EnJiah/iZzSaix+OVdTc/0J5IA/1JGV+6pnSGQ6n
1Rawm2DT+0sU8t1KAJYS66tnNgroCtLHZbX5UXoPlt3yIV4w6h/TBRgjcaZhH9i2HbDNTW/LjsG+
t2tRvm2CKnJfv8BSqCFGz3o089wGaMrbRW9nrLEM7G3JRz1R5/y3nN7gQL00gARo9+elEQv2U4eK
/tGD79M/WiaLAaAP7lZafEMAGZluoN+l7fRgP6TFYDFVXd9ma65f4OUain+wRVWNAP4UluJp2DSO
8v4nJ/ZxQ9h1iIb+VLNC40q+YCQvP7H/wJPpBchT679fTLeD/ThJVrFNomyD3kRBmykYxPLYS+oq
t9LA1fNddPox/s26sGoo/g+vXgKi5AaGNucUsiEFc80QPQZH6qa0lO2ONHr4kSAcX8Ddrr22tSkV
jLnrPM/LSeznbhltpNRAwX/jeCuHtJ5mPz+q1OgMQ9Yamez6397e7kkeLIR84fb6x+wxwiI9reeT
Q7jwO7Q8Lqr8AA/4P3KN65jzciMMp8JDSbZzXet9nzI9QbPYi8A9Y+HaobUGElOehomlmLziqtxH
ZYKo+y7QkHA3wHGPgoMYfC624zARPk7vMElg4HHF8FRSu5KcsMMslWSGtFcA+fVcOHYSNhgrkDem
8frUwdHVbK5VaMVcchaFndEJ/gkOchfVPnqO3N6Z9ooMqbXioGHjbYb7utlO7t1FMdppsUeiPlw3
REW3ZKBB3HqVrvTPmFWkVrVk666PeHvPBetm1dkI7dl6ZTYUlUl9D4B+76MoKt7BTXQQWWuD3VT1
V5KelJluLglqIgQfugqlPGhO8Ng7QzF8BMuv1FVR0gGQPNiiKEQUsJj8ekQg7LJAhQWOloWU4QHE
PnENP7+Wena27j86N/j8MlWl8mkPKoJijBVUIDN+xvvc2QwnqkYNLvsYNBrd5eASqIhFKT5Y71CS
NGDNsEMP1+m+Al47HeE5DS2l7uqTudfmrg4uR3Oliyn9jm/0RTFvggk4n2hIbmURU67BeQGnAGQx
+3/Bl4qFCCaZMPTWgTv1e5XuoPAq5FgIno+yhiFnlgBjWbduva+Taun8hEdnZpR4lC4CCDQgPlgF
Vt0lTjmX30U7KQ8Lh+rSpIeYRxCY6Qijmq33pKZMbSMHo4qYLz9gBEpuZX9YoWdrqU+vRmzRsP4P
LH8yqajAsh+laofWgiOQKVeQUrkv5JSY7JuDVhUHcTQqMKNaM2W3iqerOwFjZ6xvAaEbYlnuHdOW
Zh8c7K/7INWLoJzE4E4ISfEaew/fTzuwI6k5FgMc3sS1Z6E7FqJF6hqbK/k6906sUF0H625993Ml
oBXaalWoPtLy6c7vjrduXxhYGSGFjYlqkzwo43OrPiudnqP7nFF3NUOd/GnrMXRYqdyQUo/O09Tn
3BULNMdY00LW4CleZpymM32AbXuv7+N4ESQZDbWdqV1DJ5BHtG4/jDM1JEzWRiuOHAE0Bt+xErqP
mdOYwaAFdBy03uMi3JitNmlVhSxCxgRswFffASngbF0iEbj2MkR3n7ph+I2lU8GaGrUHEhlKTX/P
0fhhdRnQVZt9kju2yxgqM/kj2n6e6W3iWRn+lV2z7wd6X2U/joucRGW1xbMMBTw/KCwtj9YRQOdt
qzLgyE+FBJGBBUXuUH8dwLTwcsQw+9Iry+tSlp7QgXKRuqGPv+WhwmRgdyHV+i0V/Y38dZVQMMs+
BHPDJv+eHevgHwShZxUphBEywVp1Lmh/ov/NjiKNs652fXyaJtcx7GBwFjiWKtkTzIrPuT7bBveZ
9fYgxRQLNmipU3rUcc24vMB9UM7bD6zQKp3FdWPCGQg4rF45Ptj5rdA0gHsMCjppxMS5QsmX6uS8
z+CrENuJmRKmMtMVvlG2gksOJB79V/Z33NVmL/vJpn4TmnsR37ECWzHJp0VoyRJdJOrlcKJCjq6u
SQbT1mY0+CAZ1X/grmMMEgv1a9CotvpQDbZDy3FbElEeI1lmeNy6lEokayAeaelSOP35ozCTLWg9
S4+9SHwb/r4VsqPZ+0XKBwdfdFDvCOP4mCHJOxY9U1GO9ES83+M8ePu3YOu3OVBZnDb/+QljUQ8c
56Y4b1VQtRiddn51Y+/qrr6MlFPxqIm9+DNKydB03mFxRiUZlADDfjehRjtw5hLQ/68yQf8N6j4P
oC99PIJ8IpsqHrkXZrCrwTxyoujUqRfbGUkTg8P8bVahJT80oLMSGrHHjiFsAWSHf2F6ewP4lMnw
1H7TvFDQ9KFOeehWPOvtZ6zXuizn1H80+iWgLEhvMqSDhWo3WwyFqQ4mnCACmGhAPgclRM3+C/4o
Sd5/Ae1aGxPVSU0PPqAUHDtCaWBEK588ykKbzkZ79zMR1mUXynxgWlyfSCZ/nlBuwOIoUTQEmng5
GnaZ5PhA78DEQWuhov9DR4494LWa4VIBdHy+yA0OFkZ+S3PbCdd7nKl1nmr0CPxJ12OCk0p+bCQQ
3SJeBwethF3Xzd4UQCzn/7w8gZZbeC1mIkdsHlPIPZdMEsYhLFe91p9FXnG2gybfQISOgVfA4dRY
p2jP07buTDLWcSgqfQ9vXpeP3LzbGKI5grqlTv4O9+Pj0vt150ZPP7RXnuH6LCcCZ21CmaTymHWn
gKV9QhIR/08J4rmaJJDbFVLLN+C4wMLytD/cFThYAojuvPAa4Ota9OvDDZcucZqVlTNqNK6HwY7I
DWBqDOs5VDfubn70+zu6tRQPhTdPNTD9NW6thJvtXgnUDo0G2xFid2Wq0zXUSziNhZ5z+l1+jNAx
MpeB9M/rNNxWIFBv3eWxTT1e71Z7wJiLAP0GEns/EqGNMRD1gqgW6X3KRo/V0ocJiJN5AqnzzfCJ
IBubZI0Bf8t3bKR80eM2AEEKyzyfkAj3i5N4dKwJSWLMdKArh20wNOFWFQ4wau2wGwPBVsyZER+h
USfYwjqUR3qXytP6s297Ty7NG3wrsmA+sBoWCUGslXfyGCInfs/b3MC6ylJTcRNN3c7KE9mQ07RK
+T7YMI1mpue2Z2WLPNC/gSphhhHKSGSm/q8i87v8yp3w3/V2O4Onxcvvueof77xbYSWrSq9hsHkG
/4jrXM89XOt5/ZHeRMdF+H+wBNyxAtovJpHekfz+L8WXU46KRk2W71jnosPKH+iMtGm7jbm7sGqd
8Bhw5qI47CXrnpAENOVdkE1aXINkAtc0WnxDtejSn49PaBMEPRLFrmhsDuW/yqJxgN3ZyM3VWT6x
idClmVIYzg/xNUItwr0pPOs2/gZIk/Jsn476UU8opvvN0cv/86sJ7upTxUgiTGRVWSkmHrWKRb+n
ruaK7z8yMeyZSVCbNq3WWfghbnF3f7HvJWfjrs9jYn0EazC4T+9Az1az0yDMxX46cWPlPJ6l6at7
FyapQtEZcwsLIKR2JzA3eKzwImFkFT3+/g9HPPOxtDl7DHW7tIiwZsAhMfg+92Z9FWXWPqPv0jeF
oqR3E8+PmuZmYK4/Ki7ILDNtBvrAuZ4k/QeTdGky9N7k22kiX8MfPfEettbmzPftRBETREQATRvT
GQpafZQPtIOM9H/Q3DognHd3jW+IDYV2PJOYqFsgiiPKYPvenqhuJn/R79hHIvdrAgNhr+ktYeNK
kkJYSW+Tg3WhNMNQsjNKNpWlFMI3LA3WBWEJ9lNVBseu0kcFAlIbkpwoFhOEAcLWpd7sdUmSETm4
i+T+eY8BGHR3gFj9NYL8yytjo3gNeJplgogxluw6DEP5I9iyCY7aCqP1zmpRDfUYaIKfCQJ1Z+0d
WbNtqxamOxajYvWIYExOogRvMmCFRK6alZ5xgtoTR8q8KttoP7gvpe1GYCOczQGkBpIiGgCCLb24
649e2Mseod/0L0hS9OrDNXjWGUMeBBYnG0XKXbYcHSplp5yefFH/lY9eWh2YT5uLNs4McrbP8z0K
fXPoILfdFAVzPAtLJZQ4txRE5B4vZ36KqcotQ+evd0DQQ6GXL8kx4hm3n1/kM8BWRmZfklaiTMG1
j3ImFe8hN9H6ENalbP0g2U6YdI0rPVInQ/J2oIqGPIjt8vUebPNfmqCqMF/ZUZ7Ck30/5kSPnB0Y
ZEXu42DmYUtbCbhQ66wGGr8qu9G9rVK4319RNJ0HxwmqCBm9uOApAjxT5TxNQLX1hG+sUkuDSHPV
IqjF7TXZhoY6MJOAp9ju8arCC8TqjnrLXkxJm/oVvftop+jKxeDCYDZrpLuxHVoMC9oEbME6LtMy
yoilk1AlRegwkiBR0yhLAaAnVB4UsTgT9K5H3cAwiQws7VCqp6e8SZ2+B+Y9f5PFMbLEcEtGBrlw
Cz1o9qUEvqzTMgTDJtmZ1MqLxX732ceAmZ16FXfqRiF1+7oyLSdegoLnbY2UbM01OZf60NnqpzHw
9D2R5FdUGYWXQ3wy7L0SheqgLDD9/uGLxWOBB+ARIk21Sg12r4R1ucaMLiQ/2+exHAYH8K68INmD
3r8I3dpqiUnMftxMQqAp2rdQSYCgP4rab7Ua5QfbLGSJUKUfqiZJPzpBWPNQQkddHOer2J99euzE
KC4ljgvjAuddohtpOkO0hlHZjfbEg0iJQ3W0c+DkvaA/Un0o20kfgWQcCH8fIQc5/KZ1BNWZ70CJ
eWKcFkuzjH74KrjRtWUK6/eBB5jDx2SbralE6ESKPJV+LvT7xCmHipW4GpxmlgL599PxkVeyLK3/
odLAvv4ETj06MnOvcmfEPPSB6/KS//0Wn7ymue0I3InWQiHWE6Z8ew0H0KsvKsQlH/uE3Wr82zQY
Xt89895PiV7w0bKbgm2ziSKlypgLiURDlv45Unwy7O7CEqcf41g8MXQV+BonWiwr26fwFi3k52FP
y8po7uEcUapNg6nWufzepSoqnjPbcQ7snurdmCAh/IYlWXHhaATSXBorkfoyuW/3UYny3fbo6rhI
LkqpIGTta65c70/nQWdRACCxJmBl9oB7uzNumWLsp4n8n0c2Ts//1iEpjwH6NlzMWHxDfcbSJiOR
Id+qp6nTcCdvajdC8+h2KkoDbe+i2Lj5acgeYud9hscMH0doWovOc3R2RAbLZfLQOTnIGIP/YfY0
bOqiBjgPdVlc5FqgQ4f4hbARGQQL7gD+f3zQSsssgoPK08BoD2Ht47AITDFyHmncZmTvzn2wkrS7
jrh1kMPHcTKfT0XBLP2okmIop9pWKq60P4rU2Xm+p+9aqeKJ9B7tYCYLXJ9WKbFJtWa7hw+tXOfo
XvsK+XSdgYRS8d5Lis8njatJrsquuLk9RyU+P7T+FsYFMjdyonBbyC1D3R/ygsqKx6Fg77ZAVn5E
2Mmutgx8sYT3T0B8XoBDR20im7WI++yu5kh7cFyOCzyuq+NfsxUh0a0rfQMhTFzjMFdmMYqXKqLn
tlUmiO2wpzvqK/AYhxx8V76R0+WY9/SNfpJslBC0SvIRfZirMxYeDlfTNoQMhNDjsqzJgv8JW7lL
p9uqo/yVzfiPAjLJeHgJJq/1vrbvEitFFeakQEY8c9MU2KK/mIKtO8Zqi2VzaS9R4r3tnkPQJES2
LHxBMejki5mgjBfkG74KkawWdfAhGqeKcVb3wV2Dz6i1R3mkVNsfo0zn+A0vuwU92ryYoSpP2D1h
ElQhyAcNEptn7hMajIgp/t8ww5U5Tt4u5E37JrKpYB1wQKgNltxinZbddACLquMYFjUPAWFLeIQy
EJECsy+PjtfjDKjnkk8neyGND4ftUV9MopDYCY3NwhKZu2VoG8RpB3EPnd62wTjCXFzl+4xPmZ3/
NGV0Yy97mIeSfgakUvuO85+RFfMFTtZ2lu2mxixvMqfFy2TfBQfipASDs13OPDIbFSZuKmBrBEmn
S2ywRwzXBKzLXG+9gr597FWbJq7b1c8oDGrOWZgAnxduigem5ANqc07SU0gl3MiH9eSlw6LyL/Qb
Tj2rrDUC4vWjAclxprDd5EOIh4KJ1ajVIjWJqybe48/JPSK5JQg1ANM1Pr7HIBD1a0XebkuiMLu/
Bxu7gogCgtU4KILhsbY2XLfd1eppfmFpPSbnemaTliddZ09tszZypOd+j3jl6p1PRTwmupX+fDqk
H0YFTFbLI+LbBO9ANyPxZk1JU0Dz/+YtG/Ax7HdaS/6NwFdy5buKymiSKMWYL1ZhImEI9/wpWUox
nBkirDkv6scrCCDfpPSR8Eh6zF6/ctA/E8C8o5ZmOL9C0bzr/bbxSJn3xH5NDtn7Za0oI/LtIurN
FoAdPY1xRfhaCOJirmOOFuI4gvmZGguLtbUqQc8EzAM5cmzjTj+H8CugP57i6eV84Y98ikaEeSD/
A4kNCObMdHo7CCjF+XQMhsvdFCxeemJRWRTN6sls+/qBay374lc7s0iBmV0KLouxOzD2JU6h+gi7
ov/TEEGU+EifHqsKRpCWAunKP0JrCc48whq14xwUYDc5v0xtB/iDeay9NyNOsl2C3sv5LbNJi+46
mQeGmD1MgvYRgI6bc6xMDLV6GG6KGs8Ofc2TwmHEc+7a2qLy/mWZypf+6JjcI9fBLwuQAsl7A7ws
r8uJXKxUO81Mp+uS/+1UA0Opr2pO2krMSplIVZdapuAWGHsBPL14HGdT1oCr6j1yHmMiEn4YmiyA
MMVed4vMWBDm9WoS3YjlxziqyYdOtmldiLThM12RH36zTmRHe+auHvERgKEQlhcRDZp7anHi9eCp
VHjFSH64AVnZWGnyF0t9mYitT+dObRkkTsMq2FkgIlYbJZV89jS+T7xmeYkiR0lYfvtMUK0j9MpC
mw663wWc+fuhw8kWvJW8f/ebz0XfwzemTs6Ot4byeRwYPvL4L4X1V/Y6IFlWS4GB3AL8pgkHA9Np
D7kp8Mwn7fBijdxVDlODJzgInVy1cM4nR8KnCz1mzX9YbYvj/j9uhxjSTIfCWMHYjL3+zZEG1TYy
Ljpw1n6X+k816FrKoJTAHg4vH+cwt9JCaDPGm9KeO5tzkAJBG0eA4dt+3NNr8baJRmPm+CF9mWMN
i/Ln5PEhYSDcdYsBVQy9819nSXCzJJzTSbccGAHnhGx/HI5m3jmjpbqRTv1hZEDOhLC+BRRTBKCi
I7Bj9iDu6VOjZ6OIOcY9UMGTP9ZLpFXl4aGh23DSfMNnjsHXuU/22JPKLMewL6Ki9XtuS48lm+qZ
kkQXKV5l1M/aGGwjB42WhLRYKOJZ/dhZwJOPvd5ncsaHmPQ8hL/JS1515K8Sp1tiYDEg85UYGmAG
/ASFlQFBqzgXF+pWA6X2QtxAebUPyMmlhfgrBStHZXnxxfjFOmNcP5TTLluUC2JW1MivRg9Xrcax
Jqo159VtE4vk5fCAayCSYzyLoOCFVzvttEqjTDImJaVqPA0yZ51CXtLFZz8uafX0AsQosstFqheV
K4fDxY+lNj2NdtXqMxp6CDE40L3SboxREAoLUKvicWVGxDu9WqgVzajcm/hcR2Q52n5V//6fWohW
OOPHycjiX+tw0vNBc8tl4XGcEzp2DDgVqq6KDEbqRaPStTCiDMjwGGKutUz6oSJ0hkHcdzIXWIc6
OHsOVy0JAlc3ekZqmvrwq/WFC8RCahPTmmNokBlUqVR4WT6rYrkX+vXmyDvc9epPgOiaA3g1FjTx
ILzddKl8bxLlSin+jkpO1e4lZaBjbITulVaYiOtuifbOaCVoe2esUjgbX27lUr66L91xUCepmJcz
BGiOM6rL0Drc1eeFZyPM6cHn/MVGjxHoEK4H9ErVXYtCV9wXASuGgFyRDGCRG/72aNi3KWf30urf
V1Be6eo2mHQubM97Wq/xUR7jsR7B3N+QmDQawQCc8DgmEsNz3oO37lztOiS6ST+UmdH9NW08wwde
IJswtEnSPHSaEz5k3M20kfvyWhHaGsi66fDs9kvKGK4yKF38eKzpNPEY4Gy/c6chWFC8yQmnEwMV
AnNVlwK8V9HR1P5bQssTwaZaR67JGsBvoPYS7X2iiaTPD5Fhxkgpxp/d7OIpbKX++1uERrDaubEe
bRSjJLEvR2muFG3/hnXfji8ZnuvOoHGbeMWtsN7SmRdkTsVB6UQ9ysgjFTSgJy55Vl+mIAGKTStU
pqAE8UOzyWz3A1DOI1D1CNuiF6s/tu/4gwCXKDSEKAqyh7QHbiwSWtbCZG1GCGINfveu5hG5BPm3
GBcRx28YPwKpDq0jwgbqDX5JvixTag1nzasXzFkO7t9ObScBfua8m5YEh2a7JffbCjbGdbDzBWnt
iiz2o2IZyaS6Mm3yIZjIoLfCjUYcToRlYjRbfECxvSVQSD/UvxFoM2km/MahBgt09YzmNaRzrJ/U
K7xCDFcG7uit9SQwfybeR/YLkfOUKUuoR6P3sPgmf1PiH7YSMOta+OaaGC8BP3PqCiEvN8gN3shz
HUcvjBDQEhB2R3hYGtZIY02C4TfADZnetZjkumXNF2TPBBeto+44sZkEJezrcU8+JtrFZFZudSb7
kt+U/x1CQhhtKY85kkpDqq/dIr9RJSt0xxLJ2ZWWQURoeI6fk161sR8xHHnb9Lk+UBOWZze0o86J
dIFtB1oIGdm8ReOtQs4CTF7h03d2W0b6GnK3dbNnkoMck+VsGUUQx7+jpZo6WqmfLWioHWPFslqG
cI3chg7H+pJhisXX+vdt9uF12cHkfAGyjcjBOydA3/t3QvKyOpbnK+mZU4WsVpXFM5zw5iYnWxqR
dk1lc4m3GXWZbA27XJs3U0jlXmxsa5G3jxX1Bu2fDMZg3BYsjkkMKlFuMheAlIG0932DnTbNu0TB
M2lHyrryQYoroH8AOZFg7lqGLXhmGwgWaHXipCzjwpcygAhZs0bHO+4sT9rKDjg01KbvV2v7FiQ/
17PpCqJF+lxjkZUCXlnqhLJBNfQ9nr8OGg6Z9PeQS3UqWCY8RSWOHOEhG1V1SLd07g3t588Yga1I
1Hm7LXhiix3XIHhP4gUqizHWKjjWPp+roCotiWTnX0iZyHEm4jnWmcexGANRa0hfij6y+xABKAjA
UtG8YT7QmQEw52ZYHKXmwx6MqAfpqpFpLoapdnWay1Rm4HaqbwdenMWG3KuYuZIgP0NmLBouFIv8
4pa56oXKV3mp4BI0u1YF6eKWAUzKWqySmT+/k++sKRucEhaZnWh8yKjRgZtf1P/RlbciSMmvvdmP
05MiMm87oiBSuQvb3oN2SuCP4C188farB3M0sVIQGzhr56T72MAh8FH6u/34/4KmiPfXzt5g0eLJ
ByQkYOan8G3SDWEc3435GM+/h+pmRMHo6s8/1HUmRlAVDlQWb/wHRBnePUc0NnSWMV2JE3Uqyxqa
V3mkgoS7LGfn2Qq1JAw6LtfcB0LLuS4FF+ZFbqcEPsHoUTJXC6j3ysLLomqSIA9Xczl0ekuWiUBi
k29Mf9GEo+2P8py5FuK8c3kJ1AEnIjh5cnVbKWBgqmGjstZRNRvixnUWv2S5tb5L0cuY2XSWeS+p
nEoY5Tf4dGelYwzqQUjE479efEQevBcy+2F0uXDUjLEsiNofNMDD/fLS0UNKwbvmYbV6NzzzLoAW
HHIFdN0hmd1ojVIa7h+XGyxa5gefvp+GJv1Ap0wDOrQEVw5e/YzrT3Ash8nLSCRg4NPCnIwEgOCR
xPxSDM/080QnkXHBDocURUvPwYQJvq7/H8rE9Y/VqfYJoRIFvAjRO4LDAPCboE20dlX+mu0sF40M
rpMLbtnk2z5slL1L2QamlQaAm3plX5NvXydE8dhRJHAte2pMzKRXy1kVFxIqCkJeTYgWRIfchD3S
iT+OdCFg9efPL6Ytx5x9f+L79veJb+7DWymJxbwD3MsLUshI3+a1/XyQ4nxKQaUxy/OGtYm9vp6U
EXQfZsHRSlAnxBBRxF8ltzkM6f+aWOpTl/DmfWcbUU/7qdw7VpUQ42ttvkcv5txBeIznnSTeNyvT
RHiPjot4/z79ErgNCmPv2lKBVpMGJg8RM2UQNgbVdNssVwsr746akc3ZhLUpVQjU6AvCnAiQuPwG
xPzwzH6ztOc6OpkNy+x5vHriMC3uVCKK5gNBKX5YCjpvfrZYte4ljevLC+j/GBAZqQcf5XwPNug0
PI+nSCGNoqqONDf9dE56MK9cUyU4YQHiBt45gdT6xx9yuiaAvTs0TdV8Fq1gkeR7BbzPQLwefvja
DOBxt5sGiIGFGYE488xkRl1PkuX+F4a9R/hrbu0vMm/zlSZ1XBNvf5SuBN8cAOorwiPYzzWMnBs/
is0uWl3h5tgRCQEo8WgL0AKKE1kUI/N7wZOW9pn7FToxkR3mx9GnnyPu1my0cTLV+J+V4fhMPfZ1
Eh0AbzS8rGtIKhKkW+yZsmt1aU6n3AJYwucjE6/grsfvwsnN42H+Xa7eZs8rC9AYbPVaynp32Rpx
N0JsCYX3l9GwoVX3A7edvQSnck+5mN4RUY97v90l3BNceqbJ6GJStZCzJqXxaGRrVp3xXCpzMK6P
si/ej5jhq+V0YfGgJgfZwQKsfDby9T+5W4NI3N9jbbxaYNLNEFp3w/omMUT0I7+7MlkxQ8mp/892
52YelCrIQiLt28dgnl5obB2QNTne+NYf3TD5F2xuKbTfneiy/p286l0yTb5U5YEF5bBA0jcbQHSl
Cg8D7dk1F5tZViZ33p4WzYpQhefNXiphgqwu/FPXEZqzIRNETwfoqg/kDmNHyHLYK/rF5RpKoIuR
pJbiNbXsSfl4N6vi7PnNbQ68NvYiydfhaJV3p/2VSc47sH6fQOkmLkDSyqJzanFAPiW5ouaASgy2
sNc/wV39jH8RWZel8R/b7Jkmy/rpdcnr8n1zYRbuVoV44J86z9soLfpVJ8W9QMwf9sGDo9u8syYI
H8m0j5leYLpSm6pSAyAAKNiGo0wU0y04Y5+MOGeufw7gJVUn+BY9Tgl9clfxpxWBHRtQ4oRlkh5n
EQyLb4MwER8qvLuzaYzAnrPRc4v6d/TFIT1h7iUzXp2qZ8wSPgreSijF3lgww0/kcyCyLnuPzqkI
dsMKGx5Y5bqyWhZhrGYUe/SCs0x4YeEmkX6qnd6nLZKHOuPBAUnBw/GnD6V226J0m+x19ZuVTpPb
/qwjb8nuLYEgEw/4gvmiK6Ef4AlvR9uEl8Ay9ijJz3fKUt9R7wwW6QrxOp8tMz4pQBaj2KAYp/IH
Yy9aqaA3VT6S9bxHm250Vt9eEsRmLsmp9TVTb0Ng2pc/stjj1wxMBuE2YZJNwiRqycN0XTf0IAFT
UGoGoB+vdnkIZWZp8mFUv3iXGgp9Y7YHqh2ergLyEZaC6s/7BjNpD20m42rAcNuSGAjMYgW2XtgE
OYgox1zpTocZQDR0MwO1dHibOtgEmuMBnox8+FMBJFFSm8tgo651G6VIR3JOKwsHKm5zf5dAoSkP
pQ8p76UTXq1OOSyAF6dfFNYML2JLv2O6OgBdoRiWtlwqUnTryZGZRfsI+xZWgLwnzlROVpauDmSk
/mFvG82TTVihxDfO7uoU6i6KzCIagsjmyYL+o5LSwfwmYAH+5zO7JRt1T3RlWEeBs+0IQwCJrwcB
tGDvcnM2eWccJ6GLV7SPRH2Lgd/w8sXn1rFGqnozC75KJJ6stfbqZ4iGAyDgRZEdO1dcP6eWrIb/
odJlcwdlDcaD9yre5l9HE60fPQIf1QZggJ+LaaDD45bO6k9bcLnJmaXr/tn2ydz15UpDvm8895Ki
iZMh+YAn08pT0/YAI7ww4m4vtGNZFH2yFvY3GoV/cREQgFMgy4kMQbm0FDDcVG7UPzl7/bil5r8Z
hM3mZCPmaZzMiQKSANuUaFjyzzwiulFrL+hJV918jmSuHFDdlmtUvKAdNc1oeIa3XOkqu61HLhHH
vHUxGuwL6PhX30x5w4gRu86ETEA5+peGVPhChbskPlicuvIzk/sP6SbWmP1GPLnZKvgcXmAOOTt7
6ivsJsHeL/ysBGwLUFIgJGqUrP5LIoscmtS6uiAhR62dGbSALaHLQt0e+u95qDzOMS2QE0F14Svn
g++PBreYjc+Crz4EsN/+vlUdI4jPQgr3hEEoVHQfiWuJWO4U07XggRb987RYzquPY9Oa6IRmjaiL
m9blZDPrSavb956jgn2JvnuFRw5avBVU0l9ycUKtLVLC+Yy3HrUD9pp1aY4sduJ8AhQCLgL+9OLg
t8k9wEr7pd3hObOOzB4Ufk4d14TVpBJ97EUcVFgCo2JjgewdwbzdQuIisx7wy8WhUw9d63BsplhF
XNBfmZRVKsDMIjMnkgXnRq2uXzmJeinR7ZlrZ9RKNfgAO0HufTxIyT+/74BTy8zClxmmBGVlegV+
bMpG31/PiSu40zUm28pH/OsBalc8eJrq0eebdh0VakgOywzqv/+nHD4FMy1hH6mRO3Eqpn3fLH8e
MfEOsxr+ocR+qujECZCYxtLx7GrIIJBfAC1vCpcKSQ0ibJrxgSM7xkuOHpsDNSybyPRvQ04BjsS0
q32qkuC4B5gV1uHdund6KLmw/m3wpuL8l+bMLPvxBe6OjLa9T9NUoKse2AyqquviaMQzOeGM+GdW
hHoWxQk6GmX9l6keDeFU+uLDL5WyxOtG7HVEMp7PG0AZURnmbqg6q+arymJ7LiZ/PrPHfS+N42Vv
cQj70Ou9w9/1wlbnwbWnbTotQ9JKswCWwJyatUYYVN7+bJ6FcqUAoNKN3t4XcEzTPawVlRP1s5rr
uk4JeTbChTkVZnJDbD06eaIt8OxengyXvoOJa01tCiAU45+VD4I9PBIRV8yejLCz8oZ8ZLlkMxku
mWbbCs9Uzb4WVsATTRGBfH5tHVDPLFUptMK0vZFXLX7BOV/8FXlUTmjwgBpGOMi/pfW2gYfkFBTG
5N29rwJ8LYVt/7xkomkKEzWAjnr6hVN+AwsJprY9KEDmWnC+Tn683j1EeEo4Fr1oUgrYSt9pIBUb
oRTcC+tM9uzqlSLVz8R1FmRHKL6Gwo2+Krzj+MIyBYya0qHuqgrtSl7UXf9jDVECYsOVCmW5VDM8
UsCMbIeVbVYTxYY4rkZg3XX3Gj5oYmscwYjGBjIzbf0ZbY1v2R+/93eIgEkUigQYatXDal/tE8eK
F1gT3SQZnDjVDxhtywcd9XwMIVxGzmbM7P6tYhj8xWXq1dBudqqTEeDxRkKf8XLZvS0R4f4g4Go8
eCZkuVfvT4kXxFQADdYGAOdirGZWsKEtQbmvyBu3315i6+9kWXgUwLJcQDXxCzqqtaGQEqe5Jlis
eKppjE1vhEtU9IU3W+jFMI/qTCoKTRpqVe3VMjpQx5Rf6CIvu3VM9Xrvqzbs4WaEg8RnmkkBTHIN
H6o1xPo41r1csvC6MSTnzY2djvhUlRr9Y9Sc6BLPyaOH1lZamttwMrfSx7z1CfBlwR3JOYHN1oSY
vDKVhrqiVlUkYSuu42l6REJjl7V00dlTp3PnvieJhbWqlWepsOkWcD3rgduyakPujph4lDYXMOMW
Ej5TVNd4MtkPW91Rbs+NNKzZj4hZPT/MaGb07oRKkfOkOTP4Yt99zowRYbNnmVZDqbik7T2fXiYw
5znVWhULbZLwQibli338QzrWGFoNnVkambplL5kbyNCWY1gbo/GmV8CB03wCQa4hVoeqyJlhWxTN
xJw1ozvLDprRRHtqy9B81ypTeNinZIdr4bvXPB0yKdrCx4vSEUqlblu+i+IrugXFg7az0uOdzP8v
dQZhOl1+t1/rUocYrjXokhWWanGMDW5jQPdoOFDb5u/UfpU6kmL2lNvG/h177Rdql7UNRgaGiZER
BTHFjUgyT15lu8EjqvT5VIRBahEdIwTEBIswZpi6EulVJnHGLzFB7+eUfOFvwGoPMHacBTjQmHJd
a2NymSBrwm1w02fbHPVnUt1IH8UoL0bq69zpW+yfYbiaJgebaw9yKdeifP2DMavDdK5/uB60YV9m
uE2w9mLytvTPoz1jpILEJ0lHxWkzFQclzgfiixuv1PSfS54KuYTtNt8LZwuVY/Ts/lKAcL3DX1Ig
l6+d1T1zLQdqvLAhKStlW66jh80V2eYgBVKazGO30IamplrPf3HYUj1kXu87dSPmvvilg3nu9fii
q9RhyiDv6b3pKvEJS1P+/CwLth7/aZaoP7eISWp3dJqqYiql9qV59k6zR9hHLYrprbr7EFK8v5oO
se0l5sJxvVO0Gm9qgXHjM54eXuxSOnqpk3aO084Rric7Pq67OFKfUewWFT3mHFYWoxQ27dIFZDUp
k93+53eocyaO5rOo0ChmoLXk7+X27/V1XruWOoeTjaMqd0EuNoA97SLF9RcrE/IPtLvb6Vyvx45v
E6jJkP2wyMpeJHzognB3X/q6pmiF6qkl11feh9aV4Pxjo+CTDi0ClaUyg+x7nMb2u6fkCeRgUHHD
aYw84Ev0JfcKV76rKlU9+ILGg+tDaOCIv1uRsqp8kS+meaFE2kaXCqFhZdAFVmKxBoML/yRKKlTq
csl2dMT8tSCjRYgN3AgLSTXbG1cEYI97com/odsL+qagKY+2U4FjDY5HIDx/pw6C380nCIwzl2vm
Vn0lzOQoHdjscvFWKDy/vqLYmhANPVxe+atgHeBhTg7NYyDLT8gM3eCxsTcTJLGkhdrPskUXMyox
NMgd6+54BPCAJaCcD6mNJlcEPtqPn7PrpRtZBc81SmMyQo9uWYusTPjRV9MT2Iv/a0lfae6QS/fR
alovMneNSxXwaNu0WNRNSdp9l5skTuF+IeYQhft8xuJujzuMYWKD1E3dvd15YeVCA2Pf8NbNsD9S
ro8st3lND0hpRE3CRmTPUuUDbncJRx1jfKG26yD4YgPsJcCPVFQbZe43oLXXSfC5R3bPNHR9RwLQ
4IHkBXA34hynJVI+KfPDA2aJAjBvSwV+q5XBllayZLgRTbcNnzVeoA/N33jv+TKOs86HmlMCaZAY
ZrvRLZKFNL97z43Agd5BDxu1acg0ZukzdNRROYfx1knBUtFv076KNWt9Jay0mDe0jgKUAEh2K3mO
joyIX2vpPGx20ZJaP/3i2WSlshgxj8UDzseHnz2cgl7uC22xTZ88c9t6IFwWM4XkN88GKj7lgpcq
kaGAfG4DhyDCHmC5JyQJTuutQM38gveNIh9BK3/q41ZDwqi/VngncSEvWXOpSUJdX7dH3qe7DCEj
ORqi0ydBvOjD6BAg2/pZ63w90HvTqSDdZ62zlU71D9jJc4nHML6Is8cIs/q6rt009GGfNTXyslcR
Stt9mpG1Np8pxSOFgnSrtFDFHJAi22r1p/sjgJba7p7UEtVaqqPg55LsEyWTyCbQqYAbf76t3a1r
IfBXWm4JaLtMg1wvstMSFnuq0st23z9PhRwGNJ0KpipM2Njoyji1iqfKEeDWuD6aU+aI0NkZfhHt
gg04RWCCwtkO/8qsM5RHySvNHZi3oWL7iBGqM44e/A4538jL78PtfkQnV7QEh1h6QqaLsfT4Ia0Y
qL4+FRnJhgLaWWhdYBPxFCqJxhObBliQPWp4SwGI7JtAmBvg9k9dUmVU8vJJ+fRnUxK2D+l3hu7W
QMO00/qZRodou4x0Wa0LhYNPyEwAMhr/azFB5x/GzaqiqQXnBXIuFHtmbE37KcBkaZWo0hpgbfBM
baPPFdrVi2BT3OLCQ6YKFqvpNze8rWnT4hF3cvkSXiyRW7S4XIaYdRRNaITx0Bn985tKqm7Vmiho
8uYwmO8LQxvuHhs2/xqeuFZacCFsxqsTKMdL92fdQt1yqkF46Ct6On8jc3UEdg3+plF9iqjn5EGW
BnYIYARDoRMIHi/MX5mXD9NaHgJEIB/Q1bSPKpi4pupPLKWSNk+A/XP+khYSIgxhdUzE8ifdvFXK
TNIw6CFgwKZGXMRK/etBCbeKfbeSWYxEvi1f0hlcHwRpLEI0FfsuM4RD0t37wGkYF5Qu+mGM26os
TUfyV5WHdAJn1PBkXUZ0DGfe0Ymu29loJzS3xJLfa+CSYsBaVfDpibZ+cx9qCoIIZ1xwr0ihJtE8
XLIr8+svWtpcmTSd5ibAZFCtvYbHWHC4IvQJKrYW4mGSe60Vklmb5KLoGwG1hpnRTWdcXqBk56W7
u491is84OSyucM5MyINDQP7oJUgbsiNxGe6VV9JMRN71l5GXLhWrkEa66id3V6SBRfy0pcoAnpRt
WKmYIMLwo6SFIRx9rx4aSdTPwES47nQ4H0G8YhYZ20+FUpbSMxMB+/Lxa3FdIorSNihXudvZZolY
Hyz7RvQh9ikYFk8klSPQ9WzfPSM6YDVQOqPEUwhBWXjLH2aKn7ancKR4KnqhQ9i6F0eGfBVRJhup
9qi/ZzkG18Ngis+f6bqOy1jmg9H9kUsK/EGwRgTeypFrRJ7so5KGZFjeERPXSkKJU0dumG9l/NXJ
OFzUDrsrQqtwUf06AdeAvduRo41nqH+vCowzCKT3UGXhgECBpXtJ8/gg78dsFf/icSdC6+wc2en7
KbDAx0H91W62+WGtjs3aH6qR5Rw+HCMM8oa6DL3WnMT3vgXetI7W3KMBc5pSDCZCsEba/VWvwuY/
Ui6O6nmqDAouK5wcQkArhjVEG2BiZb6uMGnXKlmOMJzka3bfqKA5YDFFXeRFYR0pUSqHzy6D/vc5
6RbPUQG/lIxpU4hCg6bbsDRDbVkL/Za8FkCto3KZax5iFE4PKB/kSYlFqKtP1eNj/Ho0reFXZKSz
hSSoYSZJ+tQUUmU6WL0Nz8MfchGwSiIGQXo+6VgfwCPhI2+SgoLM70+eR6xB49Set32mYgbKeoVR
3R4hkjnHlfWtvPi0rQL+Dx99u6TpLsJ2bwlT3wsthmoFsRI4jNH0XHiBC5ZheG2vBr43mDd522xZ
lvVsYdGyv6jXW5Acfz3mnHoq/ZBNf/Z6lyA5JQaXtcNaIc4pwa+6P/KHceR+c4vKU6gZZMuRZ89p
bdJWELVPlRtWcAqCoKkKXKxrhZz+/6FXAjgX+KMbJ0wvKlEH7CcYJmvklNEKoW9V+WNa2QLvPA9X
xv2JrQxNU4FU21vWGI5sidk44R8waT2UVd2UXLvwI6c4TLQAQ2KiUz4HXcagMdHEnrWHv6B8nfir
bzByWAZofLwvDgQDig7e29wTuv+YxHXB/hlHfU9QX4S6LCGhOaVumss9//XwtusoRKdq4YbxDxma
SfYrwXhD/eFqoXdc+FBdR6ZyAtnDh0WMm083OY0C07W0XP58WkNRjVcXKz0ZikfcKRY2MyrA5lSq
twguDoVlPREDGrH2JqPGbAN1VQ/HAcQwKxufgMPsPuTVAr9gkXZRIWXZ7zmsexihwuDHGN2YF1jX
gRbWftYrumwDhqrZsYMp8s+pMtvbPl+NqIV9c30TQobkf1XIGmu5gDgnMyTvFGgZEDN4pPxtanv3
wSe1q8sW17nef+m8csGeA4z6LOAddpW03HtLC9nB7jnYThlsW+w8TJnH9Wtd6EeDAdUgtI0VFVgK
eWcBFi7JfGZffw3hYitFnsNuITGdIgH64jCPCLsJ7fHBNGxjf8UgFLhZl8PFuL46MrK+ud9rIUyT
p6vZM1c83RzTu7qboYV1jrZYqZ2c4HeBCX5Z3OZOityAFMILph2lLp0xC0T6edm1QzZdRmkzytSY
WEJywH1xXjl+wwdSnpn8Sb8vruaaHn8c4IJHXjeN8D+MdSIgeeF6JjjOu1VpjDSb8Vb5dT5aH4Mk
L2HrFSon3tuZQ6UAYWw9FT0YGWvGWnhI/dP8HymJ0fAd7KpyTzGDxIS0MHbSgf1r2asRIemlRXjS
zKExWbvsZly15SSmzPQT1ZDwMcF2u2+Hw1/mIqCE2OB84lZDQpxL1AQl4VCnvU1kZ//zfcB12NcR
0Yclc+RcrILCHhzvTEgc++qiM4bIuW/bkJRWawXKA+enUX4F9AITzFJaut1LOkSm7W6tKI8ks8Q8
1p3y3VmHAm6l9DUWdsZVBteIaNExawIUUXjWQGwgXmig80GzQCzc3wSTYji6niXVGgFDqfm/8YNp
TUIDqzu4oUhUp6kR/RrhPNQ/bQaanSm+Xqn5LOybZARQQWY53NgJGaH7j62ntmzxqJb6FHM/YmT8
XXz6r8UzMaK1ISTpp/onUWvnfE0hrhEj02MFXRGu8fhudzzroECKMhC7KNBwdsiZ/xS/bgVJKUc4
yoMDHVNCGWPtnh6ESnOedSWZ/aDP9fQu/sW8yeIBq8/PI2aAQ8tMFSHq8qEXml8S4rcQUSPNIX1f
ivzv/flj47XJBQgyQ7CZChqsV7QZ4G7wg4WQ8nUPkTPHZo1hm3UHwMC/AATDfsrod+BnbcJx+l0+
LH64Yvd+KMo8cCyYWe+JYm6tZ9sTWZv9OahOdRDaEiNEu3Aikvnt//81D5Dw4OGhIpIooSRGa2WV
0IN4mTN2+DIaMQEwpJO0LZTCgBd1qvO4b2o22wPluegUx4wQB2V0awkGye2901RvruZ+FigluJfh
CNNpRvJ9/eSrBA91z8TFjYgfswO0CXFZYXo+P3TY1h4baLkuqaqruXTZd68sCqm8sD81i5S/xwDB
eJwrdeTofnw+/fRG/L5LdHopWRcPc12KhF9JyP9zkhwNXFoMGm7xeTcNgbd889fAfoCEQQWUotxn
rKrkcN26DK8H1AGJpkD4LMzksRn8TeHQGJkQxq5+dTtSKddmYRLME+GjUpcEP4lTYnlB74JmGvpv
e56T6bgKKT1SH7Y6Nq9NBruU9xe3BNgirehV7XIEFdPi8NGvHGXBuC7UwMqGxpjaQawRvNinbLYk
UPlNnpylfkWvV+lClrYbOa3OPVRHnYLZqMg9Kg3LVLqnsplkhfwzpEkAEhOBiD1yQxhZtI4JizLe
jRiVAS57BE80fY4DY8VF3RlmlwbN/ppj04I7S8m6ZEp2OpjZUlmwrFUvQOWZfB6hWgPybwBJj4Pt
Rqe6O7waYB2DX6xAX4MsxX/vV0FKwg/7Vo7k0K5y/4BhsXSD03zFL74dQoHpREldJ/zqlY9GihTt
oD9gnL0Qh3MJ2lSrl7SnINV5HEYmslosx+Y1EQJRT8EVEiMlUKDWkSLv8NHO813BT5oTUNj+cFpN
Qcc2vcFHwvcGdK1AKkGTlhjZhG2+hQT7Y9d/Oq6keYCMIdRRzBBxMVvAzh01uSgp0smVnwT7+QKL
umvJ3Mg8v7eihRaiATqx+cPtrIwv6/XNlBuDZs+9PXfNCN2kXY1xW2Tpmiab44i1ZchOZb8x076Y
GIKFqu3OyxVyZ7RtcNLkxXHBMdNi5na/hqrv/5AcoNufbLyjumDUl0skLszypT+NDgjCG2ccBgWw
uVsY+9+jjEDFh0XjEy330O4aqY4qovSytGNoPTIGAKIVPgTEwsyXn29AoS5F8YdYWS8lbU1acpzk
8Yx112spOCidisM2Ey9uNgDRMvUOSBkqUGtV7vpp1yWzscL45UCcLzPYeu7MAU7QJaXcAMX+5vv9
dLZWqUMgoXK0GOPUkwn28ibdlraJ/3tTCN7AnqXyK67O4t4pkACqCHCgcCDp20WFnYtKp4w//ty0
mD184wYS4qAvpVsQrWv20JVmDEKBSu7HSbhz2f5Sb7mFVgrlA7WgIYCkzK2J7Ft6bAKca5w8Tej8
FIfFPAosPCPis9Gf6j1rn5dFOuFUqghQGM857zQbYPemomimdHFz5rAw/OxrYtIprDPrlo8jjnW6
BVUEXgWnawhTQtX8IRLWPQN3RtB8N9NSzH/GcmqKKDcEp+gyox7G2LLM9Hy5bT940KjF9HFy0oBI
2ksxrWsUVodwasaokzgXJOjHfKwzj+4qvNtbX99V/EkgGlq1MatBg10Mqz1p4aCp6W4hyUWVwKcd
q0t30PRR94ZYqcO8U6dQCXDoJH5twTY5UdMcNqUpycMdxF37i/07VRJPdqoqpdKaWBVmz3ON5BLq
9xU1Ih1QCVN2FR4YIboFOVzhXBlsabsapB04B0mIS8YEPp/hL7+UnK6OmzwHMUptsuAAsZx26MfV
ODNRjtuBJXF/BKTOexDVsN10Qil0petDPVoNPFdtLCUR54orsP+av7JmHqaRO3n2iIGYGHtTdNZJ
2/eoAFj2JKJKFAowr2EByrwhTblWCkjv30a0GSMHS+HvBOMRxZIJnYsjB6r2UjTuOeyrAdsRRZJX
thFluDWQCtPAUASZIOgQGV/deMdrutAQmWSDMT7Y0GmTCJ8CL3vkxcNHS4DUf191qe1cvOGXj8F5
mGSqiB17lAOyoKZ7grQx/p/JGNDtM0ZJz0tkJMQrT+V8zI9uCue+P0Kxy7QKkQEHV1tdWmNEiS05
mFt5maCryF5sLaiR2avgh06/3ixQ37sjj3AjcMAQIrWTFxMgo3jO0YiwDljPSfzKmDqIZ6pdSabT
lixSMjXEmHDi8nv1h2bmNWr+X5TkJ81IMgiu8/PRisTmamQDXa+g7J/jIG8djQk3cWMEtLx9W/HV
OkswfroVHDSjXtn2avROGtPueIIVf+s30DT44OoEeECsgn1On8SUPBiXyXWHG/hQnv72hjrN6J4y
FeEeiGsl+gQlO313L4UyiAGqvEiebk0LdXMCVHjWtpsh9HflGRpQ+HNXkQCxokGfj0U8my///KTn
XSVsqnU1jqH2r1HqC/BhfXD2DhOJZRbeohsvCDQDwLQVytjpJCfLES3TDFi+aBZ2KPyovocQqOan
os/8o1PMLf2caHFSBpXt1o0Ewmpq7YcMFKdKmNiDPa/g10G4FpshQ9EvV2MRbVXfOTPRWbHHnz5l
QTvbIRIlvilaGzxq53+9QqTi3JkJArmEBKM/zjZdRWDf0yssGq4asaTxm/0RYPdYcKSe/5Ido+aU
NhJLOKEA/z2vOq/Z/ci5Ys0x9ec0p1zrukJ+sxjbAj4PBjPgSJqWAF8uroNL8jh3Btb976qHqQar
5DOtO8B0cIpQwwXKLckpzdKnL+bB0Ftq0xX++q4RLBzIHCJSmLXBWfkW9YqTdUAsv0Js+RSLgmAn
ZpZHJyEFQKOff4ybih9iZqTmZcGXyea0VjEFLXnJX4G945UiskNVe0BP478xjLxU6YxNQ/24VI0Q
LTQxL3OSjpTNOHb3fMguQUx8/OULV8i2ABgpE3NFps7ebVgDEY1w/w48DxE8hYev6CFdRw0D7PY3
6eUAo4Y11O62dSCZMT2hILRM2RNd94l/RGgMR1pHkPVyYWkyJDqxhCsDWMFF92QDW/IX+uqQEuIb
ZdAYDbLlOK+2H04irINwO2lqJXP0mQjLDRicPW9cWCjrvvYQQsUGWduWHWodfRe1/LEqgP9SYE1J
itasRYK8qX7G6bfUFxD4PAUjABn/atYXE7yDPKr7rRIah3i9T0WOccq9bfOlHKxC8gkLn8iWpW1k
st10nurkhxFwKskFZnoO4Q4ATz8gYPs3lAugzQfZaDGwURaeFl7oLOwv4mZ5QhjcX9dRHtAmryvz
swnGtmGqkB/pkeKB/VHw80374MEB4cHP3pZQnoreA3fHA93E/g+cE0v4178TAtG3YXkLTdM4vRdd
xYZqrKSRjOek8heG7iXafbsAg/U/O+kLVbP7AWTimL64yZ36cPaPWXiDzU5HI26ns3A5OPSxpb9D
mFEW8DqTMemL2Ek8ML66tS68IfBJG37x8dJ6fCID5JI4dHcGOJAbM7vSbuOArw2d3DI5A9bTdmcC
iwvf6s+lUCsB9E9vFLkPR8CdUSARdLrfunWgH14crp8tt4i/z3/8VcKPLhP3Juzoe+MHdPxH+A9H
+3CGv0eyu0n0JRwVUWqqxsywh67iM67Z2Yb1NNnb+TJbw4k83g14Vwzokh2kY2hJ2bWOowQFZMdt
Nmzc/zYTUD2DRuX1i0xDJP/mhjAvivkr4HznxX/yEoNwBxmCx6wif7pZ3c0tqUm7b/5xmVe7n7T6
eStqsEB0h+DyWBHa6Z4e4LJCohecTx41WTYrIjPKdS9VH6soTJ491c76wntAqI5pCSuGtmp/Dd3M
K6H7rwcwcMSl/IXrTs3tykuRl28G9sar5IVftbuYdVuB3jfjG0Zh1d4O2b2blYIZ7OQ2ihaJt2y4
RHXvPxG0PCgRyQSQ7avkVPLA2BYeZlF23bA8LHKTa3xODeFXmqzOOdYORAju5baCHvo6GezkIEpn
5wTHV1UlPDdTWMnMx+oYhkPor92OhoE9gLMG3Ia1CYS8PZkBSv7reGeR1c6HLPr57gjgCPJ4HgqK
bL/CvhEbfSfyZ7SdVT8rbnh433ydrEtZR45gEehBblLbdHotzcCKCZdGsjRtb3aww0Xo8I7F/8QE
OzqK2PVJ51pUP2U6GfVcbKfXrjGUGKH934l6tKRVGGmhf0ZrA/CVddIz/nS+jx04LEmWrAzrSlJN
ofGa9TvqIXSuBlJnIPKWJDAiV0JUIJ5aeWprMSvDbz6wXaTYxYLUAXgICwOQ5HYaUgJtaNuCPZi2
LbbLbtHnNIr934wP/pTQq9etpIeJuQVm4I+Z+IowJ9h/jBcFc/IN2ski64PTLszqwt2SIeoO/JCO
EzG3qdaqAFNKlYK+Bz9ke4vEElRWM9w/EzwAZhJmRfb+tr6wBIFihi128HB2VXDs/PxREg4YwkD9
kQbsUWoTNs2HWLWDGlWMuRoPzGgtrQffH48mNtGB8VxY2wuTGJT2JM2LbVIBjL1VMMlb5/mUiWqj
PvZLQXOECqpVG+s+uVMXqH9NwZ6hrhjsvilA37QjrhIGwgLs/7m7KHsdJBEHicRLlvNJMLW0o2lE
PnYOVR444bROiWRSLjkhdHaLVLBwW8ccgopfx6RsiTN9UBGPXICX59Y+t6E5C8oj+yF6YlQ4s/U0
8s6F7nFb2LoyOVsmKUAZ6EfdgCYeYmqSPj9jHMWMOw8uG8/jKCjkuZ8jFyRySPzzwdEqtXEgCzWa
uYQpfYudAh29lRL/GvOfhCG4+ZaSFXugbCAEUtphJRfp08391UtxyHl3tL7M5CuieFkm2FxJpZ41
w1AfWHTYSWbQ7oHMd3isiaiPTEgVeEWi5bMTXPeBufqfbS/ALJNX9+MmOXMAIm4+G11k7/T72HPs
8Fqpla2sqUZtaliidt3l41eZ7Lv6DFgTrRydBaYmYVONibBqBS0A6l4O+6zv8pOzTU96bcIsQpDE
M7XtX60Boy2nPXWM5i5Er/eun3NU7mim7bkJRiDvrHxYFDEtndbsiznNN9NOjizjMs/53VwooLjx
f+Cz0mmeH3DtcvX+kU4lYL/pYnvxmm1OI/ug8Lv6cvTJFwkhQl4abl0Y3q7cg6Mmgjml4btAVqAo
Bu4Wygadl8RDQ0YUihC8LhUvV36XwxzdQOqqb8T7KahnsdQ4ZGxrM+TVE4jsTFNCZDLNa/1hW9mN
CIBPROEx3PbV/3clifKNcu+iX4gkQqCdWyDbgV5lg/qjDHXdvSU4yL7pIAugMBZualFwqQeqf3NF
TxLLttAuQCGMmLXdjlbnqAu6tVGlK/CHKZF/p0L7hCuLMHq8VmUyECi3mRX3+H/szobLBBY9xnje
nznFS2UMozeW3wlNV7OSnDmJDZWA1i3JQ7tmkmPmgjI3lt/X/vSBTURt9qARumhqWNWH4Sg964iI
To4oDJSxND3nZObf84QcUWouPWvZ+QA4bola+zpRxsNCEpbHnSoLtkuTXdcb1f9jAhi5MzLkg1tx
73j6vwnHOx6bcauNSgpsKRUU6SjZkAcpoYZK2LOuPX2E7Y1rzq9DwV9NsqtsZL+Ce1DygDdqFhId
9T70lnVcwSm3gLABh9ex55rwP2CN5r5saQrapZMM8yJxJ2tqu1FPLErRwJMi9ewYM+RJxWTE/I+0
TY4pcf0rRWMNS48b5r8sZZ6pEAtFdkDvbVD1ZGEW2etEArdaNkZH9gB1hZTfP/3Q0ZuQ/2XMXg4Y
Fas03+sJIDvaAus0n8lOyMikBeAU3qkHVHvAYtKX8F785CyYjDxvJSYwOKfswhHqnQQcvsxJ07an
pWIittgZsvsPo5RURCFe11MztH9cvCwN12zob9726BU8cg7NTo+h6gF82SOEYk21NRR4szNYL3vm
9c+sIaNXQ6+HF8P0R6QMEvgGCFUFxQwyRNiFQaeWdIrN+JNEJGGFSV67n6u2gP2c91AMpGTlDsUD
00c3osw7y4F5XC9+cM4nSQ6IPo5gvabxy75JeBYScNL9lGmtPbR466/R11ngbyV4OuzePqq+Akf4
sb/RUCF9So+1Mqn0tEhH5LMATKAtnDe2RORweyCivBe2GLytZGxphYXqrjUsGqqzuZmWLkTN/cC5
qxYqn6K4CxTMSKeJ4XoOyKid7yDBAFU3jZlgd62KvaqiPmy+HX9N9HjUQIv6ZOgGfJuV3KHwTRoN
Mq6Ua+mprxlz2w8NAyfjY3jueShlUE86oXPaLLBvwgp+zOWe27guGXtVOQ6c65xdQop7Aj6phd4R
bnENtDjXAQ/VpEoZruAzdvVh+sPCEsoBtt1gmI8wn0e1F/NzKJg99DX+/S+HybA6D12J0KMmqbTH
SZEYe4AfUHLUYoaZ1Ywf3YiqBrdPDeV2bim3h/GxPKyT8WHK6Ir5NPC63xvKOb1oW1P57TskBrLG
u6PWS8s9DeFmYun77HElNaQOSAXH3/D1oC2dTN0FnJLr66E7qcD0k76QaWmab1+R6tfUIJRmEuds
wXbGEyx9ckGiajhEn50sID3MEoEJHMsVxPnZWixYQApeNuha5j/JsFe850917+gfULDDXkeA60Wb
3AgZ458LI9TPRgFtbjWhI2m+tr3TjePibf7rIbbBbpvA7tVO5VW9fYwzM9Hi0JaO6psvvr9/Tbul
KeDhBnQGqYiITYHy4b5c/EN8894zg4vxbXTYw7+wIfgV3bhfqU1s6aqJqJY6ggWofFFDBrX7jFcW
drXI/gmpsT/qqdfZu6k+iYFVUsMsVYxVAHFa5W6slwroHm6e4dCaK8jltZ61Antev8JverhqEG9M
TLx1GCtChg79xlzdg2vsK6claaiQgXtvjYGx2T5RffuNclYhQecOvg5peFVCjtPg2SVRfWuqJnGG
EhRdxIAd2BP8wLVZMk7V3vLy+7U71K4PiU5nmRqF8wdBK9F4PDjiTEYTu05MdP8P0RNO+blRyT/+
K0mV9ytAdphPzie16gYAPo9NOfM5y+0C5VrJk1vYDsc/AUlEv27a6rVBoC7caNbIOICmzhpI120U
6WRn3aC0gEIX/LWSgJOEvkTO9GlyBFPFuQZwB62Y5BV+S85sIfe/iv2xHCEsyoiMoFLBPTWpp3S4
udcw8L7NMYzB7J97j9RyFEJXj+H1HuXDLqXwY8DAV97YC2Zyh+a6PHb/QezcngINC2lV/XPcMl/0
QQ5RPR8EKbK736nZta21wPU+oBbqMWKdMOADGaHEW3mK8KpOTMOnCX+s8EQCo+Io+rk+uo0yQunw
yhPIyag4iaPq53mUKaFQE2jmD8QC77X3eNFK8MTe6jDwbOOV7bfZcwedye28+1aJ/Ud0XqF3n339
Bd++djmqUwp8auQb3+5hWdoe3y7mMH8FdStQioGb2xpAO87ayMTZa8rxrgBcApDTZ5EvpR/Lkhl+
y+1twT0Mq7hwrqCXu1Veb8csLClq01daiEb500U/jM2bPcC+TpqNDxyWCsxqltb7HgigK+elbm+K
sWICGM0gFCJ84NH/+jzAIC0JK4PiEw3qdCj86bvqNb344mC1iAxqJ7+UxuNRFCdAgCLJwr5vNhq0
CPFf1S0HejZbxVJF1yYwZn2KxHzBPg7FtfzhC98xF8w+q/Gc3TuGtDHkwb4ssdWH5Ujx0riZVuB6
IZhnh/BPGTkuGRla/XpLT2eEU73YcXQ2QE4yLb4y5GAUgwPQq/Ut7dHK5yV+V+NOsch+73LDY7rR
kpFqqQMaTB3ETc5wRA7j/9Pwmi240jZdVQ7+KdY89t3oqm6yjsfcOSrwfP0dS4ATwPvm7bgUioC8
vpCDzTFS+6lKBnYwKoWO4bRq2gotqnccaSVV/7iXT8c93PMaDZTDRQLI4FWiJvROcnbwyWw80PKm
F2vZF8CRu5aDMAXkAiURTKE2ImCKjr+F0v4MfN6f1lYMr+OmbKNXQrC919Cp788buqhHwCr6GMDV
ljnMS01/1n16JjyxqXr9ANG7hj674hh+DlkJf/pjyMZvDw4YYoj3shVhYIZpR5G9F0MAe21bHNQo
mwjnPGlQBBi/kp46k2dE9FB6xmgoOtADXuhP4BkufmSIYseCegNl4IsOqYJQyf9r4nOlwRpV4JRc
KkoDSUdjPhO7wMywu/8aqkc9EGKN8+FFJmCFaUX5Mk9rjRuVEHamMn+mZHVx3vrESvwyZZ9Z3A+G
mACe3ZD09qSakhd1dRSoxFDReHMC6ryPAgM0MJxL9347MkhlShhbcGFZ/zEHtbuURLQ0P8RGw3Dv
RyAwb5cQ4dh7jQNC2axRTMdImYDAKCjsMmN9ut5vHBqSHO13P7jgL6APi/kRRjbKzcm+Z6L86DIR
BrXw0TXQ3J/dryxy1Z8qAhvhHfLnYpVbjpyFbXOEJDLc2ZQn65/CqyRDxayroeSuZA6rPZvL3V63
0w8lSzDSU/f7Id0Yq4cAoay6lKuyoOesJAoBne0mfEqa/ny3Jy3dO21Kg8Oj/Vgv/BQuehQX8jfS
EReZxRg82JGFw4dikk0nJGMx0tjlbuE2UTSWBqNKupZS76Qx/pwdbyU5fiQtRCvC6C3j0zVVOdBC
REklmKyr6cnLPetThyPXlG2J0cs+sQawZOFMHn64wVYXdKagFvpnT73zUdTDrI6FBZZx+TgJ81ud
SrmmW9YBwLCQCyyJXjxUFpK2//hoKLYNVlU8HYL//1yyQxUe/s0BVi+d0hGn6zNOhuPGn9lMN5nN
flI7yjXvfBhghbzOhQ6kECE2X9MO9DHOtfxYdi42O0r9LxNMdXEbZGhWGG/sZwsZ0b/q7qP3DmL1
YtbCJm5F0ncaQHdHKakiMMVsO03CBA/O6Nwtu7MM72aeS4pGRm11pdFJQZXXqAZEawz++xS6vnNy
t8O+AvOklANXVtT5De/q4x94pQ2DHA/73C0izWElvJIezyryZ4na3hKeAjsmOnTZFxHBx6PivY6t
CP+SCdUBiNHSyBVdDckYe8k8sDik4cYIhEsvGppkf/PigHUQRDprL5gKe0Bw/8TTzK58Cy9YSAKL
qjeMZSe8AOHuA+3cxTtMXnAbUQ7w6Euem+C38aQwSzmAUzLm2GtV/Vsa7MkfUqQgjxs1rfWm9Zkt
ot7SDlS3IcsSX7Ozc1VNRqDkJWVTxQ0u6itMlBN9j0lXwfbXNp3KUz3ZajRrMOG1qi5T0ILWdisJ
zVW+RVGBc8FiCiaMTwxcd4RcPjMzVaTyH/anWbwsCzNh9cyWKrWoO6j/AF6fbZexdyw+9avCn94H
Vc/fc1pAPY3KrDJuoI3tkZ/cdFaxZSUymqLcs6vUXvSYNHJia8jluDZ2azUkjQJnxFzkYrA+oEwJ
R96UnnX2FbRKHgZdrxEtTp01m9+ClWv9qS+gZM4WWC6xN5O5YRoNgfWpNYrFhUOjSHRzyG0/jhFz
v1wgSojpM1Sl7uSu/d6f8TP+UUYOKxfF8LdBAFNTJ7FcgzAzHxW5tKVjKaNVd7aVF7u6UQFrLP+L
UzQVos24bsTRe0I3/Gt2PfW36wxSjaxyOhyTXVIuplBq57rLUYlCvh6oSuGo+ECvqtEx3oH0PtM7
YhkIr9Z+cvZRVPc1adZ+JdabckwMqA4hA2OoggvYciLZVGuEUkdnYemyUbDcWmiihqmwvIXv72Y1
CH0SHB3DaUfGvbgYM/vaOIq6jZfGoMHSExHzCn/lkFzht9g2tlY1bBwo74/VSVtTv8Q+HNNOmrKv
/ONp9DnvNZvudlSoAkFH2NBJkRQhl8W98v6I5+jk5Rj+tsiUzMeHsGkKliq4obvHDwuwK8rzk8sR
AVzHOshzmx7K+aG/MlCwoUWTW0vQ2p2eOZYASvWTUAF+y88f0izi0Ao3hxQjovBlkKGaWs07rV9o
JNPA8rJxc8v4PSAO6C2UF3mjTw499g7K+p7kpR3DLXGZxYXORNHYsHtlc5TO2hoU+foalK8zRYgU
SxT6LRhVyQW0ftL7KUMd9sZiH1dXy3eojhq6BfwU5QUUD7av9ztDm6uHpS/Q+JYdDqq13tq3oPQD
DyhSy3t2E9UGBnjOyWu+Pv6pZubNq0c281c0JbFWF4yNUB9hglXTeUfm/bY4kT8X9mhxs10WKcqI
4K6c2xzKLlYOeoMJ/DEbn85Y5BRdHUXzNJ2WPp1LZ7G78mEplF3z27IJqwTqD/FLZtemJQWpHwYV
PByI9gXtqelfD35pcldbKUH4RB+1nKlapb4lRRWcCJOMUUuA2VmFAxw6r9K7mks7unEtp+KIw9wB
w0PgC77opZ7+TYK/JVGqmfOaX3eMBh2u4/yYGyzz5pq+LRgDYvrPrJf68kfH+dJ/fv4d+gNd070h
vTGcLCmiDA4Nrqty67x5irPBJKt0Ci6YBDWG9J0py0ccE/JA9DCLbfdXuetilECDtcEOlp0Y+qf1
qMuK3u5TKoLp1SX3o7YjQGBzcpVgRUUHbljcTSNWv5BgvnQVU+oJngAYCxtivkTjBl/roz07Cuna
4JvOs5VSq+hEted4Dn5B0UwIQ4u8Tb2NOM7nvjhH9Cdfh4mdApqwtH2VdKKEzzCkHglclpIHCDxh
MFNCfw0xaNJwcFbr/Ew/OJ2w7YkbceqJkNkdSmlXTQRoX/j15qVLAxCJqCGnJKJSQHlhFKjy6QWH
R2hBH2jU4tdfSl9m68rzpv/55ns+drz3nbun0HLwt1R1bxEPXTVJJZbwApcgYxsGKn4GUTZ3ERZo
YLfxAk20QxAK1KegywNLqpu+/yI1PWuZiOXPu+0dyj4Kh7jfti+qhOK4tNKA9NOcN1VRW5q8JmVn
53tmswKokk4LzW0GidBlX6Xqgj6L8xr2n7xxGYRGpqbtwwgU1K/zX1m1qHQW/Jz2wvySCbj2nI6g
Prt5sp2dovIIKqkreGAE4Bj0ykd1aa0bNagKVy/B0ZoXsAIDWxMwa5tWC9SS3s3MI9LEmjEo3p4B
y470KXc+EZCC2sq901JWYH8HKLrjHm4toA+k1tVivGyCTD0UoeI3bAzk0nffxAxhsW81VoNT5X5/
m5MsK+UDYUxlfPWtaY77+c8T0hP4l7My1g7PcmcLyiYy8IENFWltKbqpAAe+dX/bjhv+j7TKLPyH
UJMr5VuZ5VSpAPeO0MVsyw7e+9uqhW5DaAC4aeh3QMxOEh94Dsb1+E6KZyscr8sNYmkT0m2yymu9
1P89h8KG6S9ZGaMBqQ0KDb1mvoEw7GHfJVwwmf7RT//9oRSKZnhYWqqD2WxrC20xN+FP7341dSfo
qXKkBqNK/PnU5Gm+cYBkg31AQHyI9gy6gsKjNWtPVAqYDMzFWauEcaORB/wSkmHGUHFZcQ8kYmlC
j6YOzaBvnZEOP2xiapMNEXjMooRNazM90kW16gP9YTiccDDDb7EsOu80QsN/qQttgX0OfSYL+yEh
uUfPdH+CS62qgwkwb1lQSyCyLIvFfH1JQVrRC0zdlKT/NZ8jYhOQXkEssw0/RWAyQ/9zq1O07RdV
/S2fMZCCysUCQIazoqWg+cRsQ3DBPXInMRlyiaXdiPWCvTT2V4MvE3RktjIPcodrxHm06sUzUeoo
JWE6fTvf5rYvpCamaz08CPsOFZQB/4jn5q2CjyOZ4af2M36smjrmWgGEfUIPQJSvzjw6R7PZD8Rd
QFabrSlJ661lBCey4JXarHWCc613afHq3W7Q0pe87HOgVd9R8o43zxHe5fc4BXJxQpPvDKo4Zp+8
cMkKGL0xBfQFxoYVQSFdsyiG1JNmKaZPnjlI16ENsXkbUNxbl/JLYWFCvBUl9UC593lLoyzy9I2J
CuJLdZI5659OSjVE7oom6hiOWzitb6UwBfICBH78+Ac/IJa46EGFYNJztkSXjO73Kb63kG83lFyD
ZMXCdUQaaCa7Fk08UaLHiJmyyylqOtBcMOGpcC20nwq1aFnBBZKZJPXHAuh4FLEGrGJXPk8+3iXO
+Tvt2HCRci1N7lb9eIZcWzczTRk4uhNxnA25ElLiQ/9md09T++508qkx8bdttW+1FMrDUbF5LpFR
0SStz4mmAXgi+uFWEXhFiVpJpt090ngNZRy2E8EDl9czVb/CzqVgTzdqXnQR2Cb68KO07HEdZ6KA
k6KdEwjwtdHF9lXTB7u/c5pp5VHrNPaHSNlfwk4byhU0dCy6pTPkflTXTRde8j8pogs81vCDDQ05
xgBUzFBvXFYKDv+s7VQW9c8/SlogZpjA1Gg9reAuTSKfcE+bjXtKz9eQT077BUggRmmGFdYdomIL
MK/mVrM0DuU9sgSVSjMUsAtPx/vyldkC+bUgsjXdtkk5RJpYn3PiEbe5ZQ85HqzJJy4d+oU/3V43
0xG05WYvo2NLCdSz026AesjXqTxx5WJgCy0eiVP8rkWa5CF5un9F0Fbk/mrXvZiAlUMM6EhwuxNI
PdP9deyQN6PR4mdFnQ2OPbAixI0b+X2S4IFPEhFkeUNpH6YoKCJh8eItUV/KCrvlDhw4OThu/yoW
iTUMPP2MqYCcIGON5rzZLYb104wV+H+wpOIRzutMbkjZ/V0angHb2QSTy6ORoH7IgxDVSnY59ZQV
hQk7nEBTmHN5BiwppimWT5PCpbxMfJoATzvrxA2piw6E6sEaiyadRKFnBDYUwX8h0VMX3k6Vm9NT
JjzkWpD9fajnoyNbn7jmkrYuVEEqK4lhhlCdbXxc8sPJz0to6tUNIo+s3OgDelV8NRwO9dOo2OZu
lZNkPR7/AZ2I0VN0fSv61ceHj3PG1Jnw3+Qngp6Pgx0jyk7MOZBMdUFpN/1CJE+BFFWeBvsOMlVd
F/74FCxMk+/ne1Z64OypAN8nA8+dDYbjYizSL1is19tzLa93aRgQnHAE12afAbt+k6up/EleAlSe
IukwOWFDvKYM36jlOCvkr4rYyKRLC8/U3APdzky72g2EFOrPvpHlQqUtiHFmLKq3HO4psiMDwAdp
OlyyrmpWYfogjs10oAUYadzF5qRnpETCrg9Tfu9fy+kp5RRZepyh6RZgv4YcH0oZ6Udn5MbvbDdQ
eQYiOD9BgTUvqkxPfIZrtGIPEo6UpL/Y/ra+nyPyOGglNI4SV5/Gs9qlJV8aCy7FxzJvNiuTXn/t
UETWqQ2JfQUaw10GK62qzc1XskvcnF8J/u9G67Lomd/C5pB8hHNhQO3eG1Bf9dlgoPPAhxrhgga2
1AuYb4CQ+KCbMeyL8TklmcMiDc0dge9HpumIH7RdKPzvHYoB6QQ2NFhPSJojZPhtJpg7RM01xA3w
wNpYPr1uuA7gJ1WMtju3jJrhocdVrQPrSqGqIS760sQvUGmCRWmx+VS9JhEVtWVdaUN5upknS/B8
YWqF9sOvjY/qXBAhCNPONLBgaJ1a56hF9p61WgDaw8ZqvC6dwJcqQym/Id2XAk02TWBHpOG7u//U
rNrSa5XUgKxz+KrWL4TDt6ekKwQV8mGJjZ06OTwE2NeDzVvQHBvTZOhk7lRxuB9ZiSy8MpeY7fAq
MP1RTkWe5gx/+WsvvFYPRgTL+JYgNOjte1yux0lyftgjw2ugQr70ieSZfYDAZgBgGnrgxOXW9TXl
mBQXcBj0doSf4hAkOPSeTG2W2u+eQ/QVJrecKMVejKGG6Tud3mw85HIFzdX71cvW2ZpeaVWyEc36
CSkyhzNRPDRiUBQ+zf0HizSjsyPsNVq6hSFETWjO0q03j+ah715T3QamVVQKq2rsshh+i64Klu8+
drbGqPvX/tEhOcj2X4wlIk4JF7YzrE4l5Ty2OYluCeG7qyp2SyuQt2vVIQdqhK2zojU2MqHCT3jR
q06vWvwbxGDmx0PpgmbXxxZSvA84dpEe8P6Ozq+J9O+FjH/VTr9sUoxJpy5bjxx2ESxCDKb6oKMp
+esPTn6Z6Bb+55wLPPjymHQVzUUZeHOL4xqbYusXBipPnV/WLe2lbQBPoYYS/AVsmYN9OMpxksfp
BwiWYVNin064OPcgHWwcdjzqvj0Tz2QTyYb4ybu1PqMwV4k8OCpTXz49pJ8IOpeNFNBOwxVbzurm
oCu4qIQ1L9gKXansgZZaEFkN8orHh8J8MZeuahxw7kuKfl46pfHDyl2+rSsxjldQj1kvF+EEGLyH
4YYmWkybu27D5m7vC4+EW3zrYXQqrCgg3Vo+CWZB8q41qgCuTN1EOCtRpuVXztRIvrzLtEcZokCf
WXHWNSf5FLw+IUskuW6zB6hxTabFQfhBGp27QDFauWXyQqNVlROYs+4EPLLENw9Qmoz732TLpq4N
h3ovowo0qsAZxCvD7dJpWq/2dy350txn2sZJLAzZYv8wlYXeN2Tbc3ikTyn4+LHwRQ/YyoVomUzA
VDlRkH9wlWlKyqdxqvKWgX35sJbUyzaHZHKPKLJBXMfqeX4EgJ2SgDMG2ddElF+c7t8DB6/VjgcK
FvCvympi2G0iLb/4HdgQSV9WcglRacqEFGhDyQzLQMEQZmRR7/Qs4rSjPV7qCsP7crW5yB5wAFrb
fK+uwUaO6aKvBs8M6KjnRcPC8Ok26khK/R8Vy9Exud45PY/u4SkJdLJyXpDUOwehFvtovcx6pJvt
tEuZBp44OF+KfZJHfQsOpnIG3WEASF5Y8W0nCQt+w1vUfdRZPMrjSJMYG06Kgqx9Fzz8SLxKfGHT
h4OKbt9UkG2JBHa0Y0Lf5JW2W5FVXljLKdOeDZTn8T0ZrHkTxtqex0kwp8/pSxllr/NlKgm24k9l
ymygM+CWQuPCfx5xhoe8CB1U5Mgs9w1StTbQFu2PQEZ0UflSWvTJRNUwcwbiMT/IU61EXXym23Oq
DcNT6KP6SzeLhu+ppiw4hbywX+lEUtcu89V7QNFdBiQFwpxakvtGq/ak1w+8f3TmriQWXOQPui0H
k1AVwjiUeXDSgJFuR5m8ZgmehP6uKnrP6rVS97OVDLvm8uL7Lx/Sjz1jaaXqbjgdFzYeKg9iIhub
qt2Uu6AvP/iVFknKiy176cizYcxCrYGgilbUV4h/vN3MQ1yk0aXX2s3VZMeEGgqI4J1FVdjczHYv
lGU2leAszbDnA6E+KUqkA9oyr0rSRaU9ZCfPOewK56rUrYr6CTirPPmGCMjbLr0Sr4ld7pCRGNnx
U9j9S1LPPvGOKO6FgOujQoPvHhGs4XxArkszxEsINLArQUed776pNrZkfL77r0BLa7WpYj5RibmP
0Fe+cGCVdiXYpCA/F5Ji6CaqD+TxbEPLHO4jgcjVtZYxM8Z8OEJMnEyFHjAyAVqEhDEkPqOXVipD
4/3uOyML8ijzPW22r4uraWxxivhBoEePGjQoEQabCicyDckKdTA9Nuu3ZS8RkaB8/uDcsz9qVSWR
5W/ff7aTzE7FnkGFkrIM1U/fwnCRB28aU4xX3CApqEm+pbUzNV6by59deR0IMv8eIS7k7fMa5psj
vN4g4I+YFNvfb722I4fI3sYVIfz02y3+pl5TKnm6dM7dChwHNleazS2NBOSeent061VKNnqQhTNO
2Pf+jkl7APNUPwLfYy6gvics+N0C35pkCnaqaP8MvW5uxBZVQt3rLz3M2x3c9cEwXkaMR94GN3ji
67lPeYMOKokma9IW+u7Igrqy2XlKwYudQIG9gaYLv+GDAnroOzkhnWCCEzBrim6h1XxyXfVSFh8O
THXFUS8MpcehMLdXUJ3AP4/cbPQ9VbchReRUrkedLqNdAmF19ZEXMmICah7OnJpXAdw1lwH74eSd
RyQPAQMTAX+RTcVHJ5lkQm8V60EuR0luFQJ7s+7oLN/Qo61P4ZWDllYuG3yqYVdXZqM55Ydp2oY+
7QlvlhN8G9cpiy0bVfU5d1XGlxFuU693ulw8P9UERD1NGr2uxJ8IDIsufmvIAEknS7sILUQAVFFm
OjABWVbt71BA8uil0JwechU259Pbumpi+AsIq38ppE7P/GEg7tgaKxsozE7m8b0+RVS3jnXkEhVx
NFdIip4aXklN243mcmQYfj7iK7z3smFwEGo6SnvhlBBfemxuVA1Z0VF10WTNhK5C5B7rNw3jcBW9
BzahI0RuEgTbzAj0IBDRN1ZMOtzxHAfrdnbqOg04zjIykzp356JKpp7LzUSWOZx3UnOxGzye79zk
xAhcsYOoJ7zXbDt0cVMHDHQWo/e++c2oV09Mu75kPkW0xCZ6Y7X+Rc8wOoBND5C15yTKJX7zvzwL
bGlEteS+u3m4HjEPPaxugyZUjtlhkm8IfAZzR1TuFkJy1jydaKkknHqxaRJRFWu8JYAEw1x06vb1
cimdAplyyJEEJm0g07O4lu9VfbMxKuU5dkRUdI9FxYvukyG9DnEQd2c/1+p2gpMAeQvvwJT3CMvn
MTWZf8XpWpm+DbQdU1QFDT0AldsiPzd2BFLuzzl6oZaavbBS1mBsFBMHe98ehRgs6gjHPJLJ3XQU
ttcV1CGGS6X8T8760/I5EfklsP87xPJ9ZxPRjDsD8DELRckiA2AVrBSe07O7tiVVirBO4DELcAgh
RGuKZiVPvbDGQJgqN5X14HMEKyjJlQbOokB+mX9ySTpAeD5C3hTQgcbh9+9FhsfkJT5/q5cuO8qb
L3fOQXwezJYEC8Ppiblc94p+PyguwKX0VpPr98wmoGY8Q44vO+epPgKuzu427+TyK2w/cDe60MCW
w7Kj2+OOwB8WqPTbdtmgCkzIgeHYX+gffvRZRUHib/iMfCMKeSO+JRw0xSbQRXwBmopS3VfUtCZT
YWz9r+xiehOeDLBzxP7PAKwJwQfrddMB8pD+NbRToC2BvDoxkR64FXCT9kOF4yoTIBERGNYaKLih
WDZKOWX1sKGI9c96+J/wGN36GZGln771bL93IaqVDcW5oVKyPyxUdNb6jQMc6b7nKzC0DFNCZMdd
ahU5uKzCl+Wqm1Sf4f1k4Fy9bx4UZn1mvuSXiqxdzll51lIiO5N2Iz1hrDijuaQnk/kfxCpJAB1g
1URigrPP/NAbPHiVWH15kBF6HSBFbLFTW/DlhFEhKAOIBXtaN9OWII/p+NfelFd/0fKFpS3rjcoa
Awi61rnVVw2c/FL+nrfT5yuM+nDIJ3XpjiwvB4dgn6aVc5U7nbJtWddBiNC5ByVL02eVebYRNDsK
otEDMMMdre4WfLjMewn/fIn8cpvyjX2hZCMRzx9hjLujsofvpeoMPxfPoQMchnZB8Lv641oU6vF7
uTvQYE0bTp6NiMLbIJhtPzC2h7ZMx74vfa2EEnVbULNpbnN/X8usqIcHoies3zBlaEBLkwRD38QK
gft3oZjdEnt3tG46J+3ZKwY7U5BIOYs1t9fO43ZCX0GUxlmDjiBtqwlDjkyawHJiHfRELwNXqSZ7
xEVCJjMS38Ziak6M5CueHjXYBg9xVOphjP9T51Q/e9rZucim1AkSRUfVfRy+22jvI2Qb3dkwkjvf
JKsvSGzsi+cV9ER65RH/2e+iHpgd8+EV6yWErgHOwPJUu0upT1ECXMFnDevDEVOi4PlALQIGjccG
V3R8Nl52vecB0R34XI8fR1A/IlWTFGzMvKzT2hOA+5bbHD+FXGS53DNfokA/XAw6Bhx5NJmwfN3W
iKzzrx/5Ik9WXNIu0g1ZtqBjaubKTbulp09+ljx3zzTH7kRnUEkP1o9mAU5SlrJN5NlrAnvrrDNP
JMpp6+vqgdkswJalDbsS06yIW55gyYDlqL/dSOmJ7uymMeHWpwb5V4OWK+3TQxubBBvK1j1uBJn2
xEzcfzSPNM5YNQ9C6cgt1IDzoH3KXe/h8gzn1RMtFnPOVfgV4ujLaoCqs2/Bsywv5MyLGSWE8KnW
bqRd2+gzxlBGijXhlK6T4AM8OF9ka07nBMMxyUkUh9KvZjzKL/z8g7nTBLjrNTfDEcbKI7cSgATo
a9T0lt2Rmk3agBAJIrYm/1cSe9tMnnX4TUOLvrrS9Tk0yJ85MDtm4dJ4C6V7lU/BAzqReOlHlqXB
foQerXL6DHvpkZMEbEZuYSp7qYyxy8v+wZb6FV+rDNbHBd0kfWmFA3AWhgzpxUYIgHkjwOcoZpfi
d7E+mraG3Tlg/T0IySpNOFDcUyF2rG0IQUz4pB9SZzACRgGASSveh60BERt4j/0G6Sbabi0hQT56
n42S3piR68qje+dsgyDvxHnY8u7xQojiYXj1PhwfzGGVyuJ+cdP1CdzpsnOD2q6pvxdAwP10XYcm
9rsH9YD/Q6fZOYTzR8hvb1B/1zM1D/iaP7CwP9B9iRPqMQvaIyc0lsUw89pdFPtZBHumpTbYIXGW
6yxvSJv3xC1knr3obJ/fCU7ncILUUKchYXwKnpJPpBlIylyS45J21Y9TggzK5+jtdznYnLR53Txh
PtgHjAe9FPenic/VBP2yTk8jAvL9I/2ig1GWdHLq/UVxQ2fzYo7vb+aff3fs65AZuqttXzJQDpHh
HU5HSfddowz53IllcSCwEur6+XVFobnOpb5e6w10Z4Mu3iKLECRVI89X3AAnQFGImKOb7fP6RSlt
SJje2k9erqI/WXs5TQxGQqw2KGIUwCtM7jDB91cSuFbGOKAsiyWIVbgXFPZNc5UkhS0mWFWbXHDp
6cZgEO2er9XneIIOhCx9HIXP7uZNVO3ZQCLEc0pwNhbqWVNYk0GYXJmKpRuDFv3G2OfETqJi+9mN
HMxjs7BpwrZygK5o/eHs9ODpJ2pjru2KYYU3Oc98MdVNfA+O78uI3a8kNqeLdvf7jGmci45TCxON
wjEFRnJS/LYyGgEfwogBvsMw21FLzWzznUOkG/3SBXgxrREyZl2oHxJee9FI63g0fIjIi3nX30LX
cOTLD+K9isDzR4Ep0I5rw+HyruksONkgKRNun97pm+LFWiqCReXGHLwpGbOflC5VyInj4iCQtWdH
qgfU/9lxcUYbXLoMHuL0jN6rKMMToikZ1YTCoAGp1CbKsxNp+nLxZMbXvM68EduUItbB1YI08KB+
cF8QzCEdcqegXWi8iMrn3xKuRdCs9FaQOT6hYRrdnBOUiHN36xxS4Q6Blyn7KlHLA/2uVAyVKJ2C
9PpINzE8gVmnfRx5buUTkXFDgcCD4MxsOXfiAbVxuikK23HDsinXSnFvF2dRMFHuGwqs7zzXU9tP
QzcUZnYLgHNJNaGe9+vJRRiKku/oOzCRzGytFZXpClV4LSF0e/6kN3zxi96R7gU+5KVYVJR3mTG7
z3sR9omRe8vbyAiZ81tfBbBcaeQHOXQo5B4ic7cVpg1mKk+8BqZLUyem/e4uD9HuA72fbJQJqr5c
SWDJofpt8BDUcEZTWD4uyDPNknmthTUQiWFEGP6nHQYxbk6TQxvL9helnos8QdCR2p3ywwEg3zap
pueJq88PCqAy1GWb+ueX2fbg/VizsuQ7A9BRhO+Y4zmXZVcqqeM6zZK3lyeExfIJZ41vXgtKRylL
BW1gscpGBWFB6n/bO/6jdOZ4+7OHcq/eyTACKzJzXI6zaIolTOvgIEP6ajF7klaBruwLo1pR9sE5
pleGe8rY88eqQAS/AlJzWWMFaXeSw0WjGRIH4OXN+Y7D7TV6oxVYQ691YG1sEKtZNiH2YhrZvQ8n
qHg5H+Lm+Y4wZS7KB/EcVWKwYkeOgKCLqSHEI/dnonti6POxJ1vQjjN+Y4TPVxNg7ifPJjk2ZHoI
Tfk3xJkxhkfoMsLfC78dlzteW866CT8zoJHtBBAngQMmWumn3Ik1ugozQLru1I8+1Q3PhUuTFWnT
Sd5Djl4bMkxU2PgseaKlzRtriU279LyvAMtS1YYw+xoEOZ0z6vCKbxC92pi7XQi6ohI+tOKwMebf
eMam21vGO9mNAd/9kHg+ghQ3qUNmMQAjQmXdCyVCxquH3VkZgpcvczjj7lHklkSNBHxZSaTdfUye
1aVOzMv6xVOEhnR2sKEIvVBiEKrNMa8NscArTK8e760Z4NALSjFB65qCa0813HtajFD8M1EjG7K2
IZNzmxp1kWMyADCbOJsKYIvpEeDaj9bjecAzO/yzDNyyFb4dPxJMC+xf0XghxigegDtnniOivysm
Huen5npOO5lKlZODwAAxP8dn8Gso1+UuqdSuCLeg6aL/oGJfoRHJgunryG4vNLfGxhfK7yfi3FHM
d1YUwRLcnYsrWHZ71Dca5ZJOlb66PzwG1U4aYGBo4JsfWqaXIx5aqM2pIyFa2zMUUGiZCyqi06F9
CE2YCvq1LeEjnYyDr9kUNxyCgGix+gB3PIs2vobv0xXWeRybXnS15JNhqOaU1vQMu2fq+Mou/3Pp
fQ51uYdv0mMdgFL+UXiDrsTSPPXjlHqu4mD7Rd7IVBdXCh0Pmvxg9jjAVkkS7lDV8DGg2r0pbuYN
ZeioEHSG58WjR2wIldBIe/W+f0nwFWjcTwPyCaqhJC3QeDQQXN9gcKzzGvSb6R7VxnIStuThvMar
ZInt66SAZSH1dntRq91eXdeEd00fPJYjSKG/bwDsDEUQuw8ayQnJ7y1U2Rm9F/eYG6BRX1m0rFiH
VY5cY7fsaB/V6L6teQLErsHDt1pKMpZaWJM0e6pjOH9B8PD4G2xEot5nWVA+6RpR0crf6bI7HDbc
sr9j1sHX34DbuvTtdNBxU2CNa1iiE2qT8E9J5WAZoo0YSn+4m3HnvYl8c7QHbzBlAZgEM1irZfkB
sO1vZzVn5LsVY4RzvzLaiQxHSsDCpCYJWq2v1evLEfq1doFDKIyc4RiOJN1s1bKymSBY8f/8FuKD
5CELo6K4f/1ayDirAlZA47xGiI1pG8GB7k8rynt3fMUnrugVZsu52q1HGwQBvj3tqwE+HsreerYQ
NY9VMJGk/nmFbuEb8N0KiFLKXrGnI7oJfqHSVSTQX4BxLSdHePXxY6Pj9KObiDu9yM8L+BNIaWQf
U9ThoiTgKwteqFkF4pH05fEjuDnRAllx50PcUP/YXTTkTmptlLRYs0KmJghxOct2BLzAu+EOhd5I
9ewqGPXP0oB2jee2AahplMF0YEwJu0qFIqpnOfcwZxnk1phZ0vxt8YQARyvfkGpnmdr9pqotxmLk
zzPwbTNVkvl58AGgN4yp8l6Dk2qjUYdeZseKYJM6gaNVUMImzOc+fLH+RRvbcoaY8liSK5DkW0Mn
opyWqJX4h24uWxGlzCodgEKbwMXpSsy1mAflGT163m61I81/SC/lWNb6Ymf/uoH6RtzVnA6eJ90L
8lFORGgsQg3jrpKFYOWrCvnwlpJZb7xCUctf6d16PUoyRSVrMPVPxwbQkRGyK9xZ6XC0eqxODUct
pNy7LeKBpaF41Zjhhy7tkoi6ko7Gcg40kg7mKrnVnxS8jREhcpDQW1B/sTnfe/tM6HOmReTHFP4h
4FHh1Y1ORc1FBTChoqULtymt/bN4dZZAi79IOkWcE4p16bdGf9M3DEbOrkzKEvC0tnpnHFU2JepW
LbzsWZ6mepZcpgzcmETIy/8IEr3WuHlVTXA1CTdPzaVnWTmy5ClfrodJAQapRfgADSwdWl9fjEUD
BPpXHD31xbtNZN/Gr5BcbGBTrmRb1Q5hJQVOrc2+eJgaSQ2bdIQvR8RSa3tbtmjJj7Hei8gjPfXe
Wk7mEJYsj0BLfLszVRS8sXdEgrM5tcGpBJcZaDmLT8H+NzpldqSRjBKnTUuxnYA/lgapfeUVXZUw
/9ZUmZqmDRBAktMCA4zb69ebBhXHzBx4BW3nEJ6Oa6kC/eYhHl18VoZesGAfHuJtj3GWeCth2Jg0
inxJgvKF1NfjhTyO0lUW+QvQeOeKQmN1eRkRsuSBE+Abd/qrYMHkQMyzRWDjj5EizNe/MJl6SR85
JY0uD+o29v8HY7i3In2oaGF+DxZoi8hCIVSALHuzh9LzjFudcsj7rjaF8VfkfnVYA2FIYZJ4sX49
SoC7Y0jrZ11WHSbXK9Kfe8tRSScLxXqrveUIHaxkU4aaY2dbP1k9hb7EfiR5a6MZhdJ1Ejn1k/iz
90/8YlxZ7oMfCP97CUknklnn7T35FuKM3nXEwuLtz9OCmgMLV6S2BsSr1n9R1epwPJN7J5o/ws6F
C9vpOzQ+wzSP17lyYsUQPBGCbNPtBtRN8PfdequkOnOTJOQy+DH6Pjfe1qGzBruMLoprDVX42UuN
EC2kP9yMZCu83O9FaJVU9NSZIhnpRer3r84QwxnMUTtLiP3ADG0mUZkamI7l3TJl0SolP3jgM1o3
4otFxR4+YKJVecZqB94V64C3hcjZqSiLoNxE3cYn3lkh0+Sc5VemyhMAkim7YeJw3s/sgiiAgBiA
teFb+EkhrKvpm9LCp6sVaQ26tyZJSL3crz/CMGU10j/0pQAmRZrevH49LwGpv6G1Gm93VcC3/0jb
mSP7+7ja5p7c/AV1bpsasbpQEDdKPkzBYoSUEcEQdxKPvIXGaE54zv5nmAgMSXld6z7tJ1PMyC0W
kBgie1JR4JZqTDsGbz9I0cjxZvYwgNP8SuTqgpKyGIURRYvhZuZQLgASYaxu183kQdiocGz7FIjx
nR3yeDGQDvlE2mIBZeC/ijCTKyqdll+/Tn7NurxAFthhjlhBXpKsLXaAnd+UYuz4j5yxfXzb9Bn/
XdJ1t8qR0vXPU3GHSmsR9JZ6noIv6bXWWf9oOzCU9SgdeX4OU1bMlvgtauYVQrsS0iT05C8Oyl83
pFUkyUpiiVW/tDoPAGuiDvrHAorHhuhJpUcELI9ekhSG1L5tUAWnD4Gs48bXKwnFg8gh+GaEZ+r8
OrempqBV7DKhdQ1bK6yR9jKCli0sqL3tqj2U0BwcQt4UMQN+x3bkPcqxrO4crfiZeK7PDCvBqWtV
BnX+g+EsEh20IhuXdOTvXojQq8OmX7Ao5xHFxhJb8+JijFMHpiD99C7kjCeUaR/2Tuu+r3R9hlnE
P/Lo1QC0Nr/O6AOXKeTx9biO9S1UI5MR3lB3xVDLUOxhQlyhhOrA2J/TFy/jZ+tRhyUGLKgIovi3
0xq36saAaznyH0ytHG8yVASZNVCKXRc4Lae9IzYbpXw7iOzaR+pafCziZ89OJqmO8FbZDxmIGKVZ
U9LHiycr3lrU5eAdNN2ZpIZd3uQykbl+uJOfDE611jV4jtTbJolgjHDa//OCIRaMkU9KaMuWfMEU
2zcvW6+yg4QBrnANybG9X5UgEI/flXDudIj0443Y/7BEYwGc8oX3cEei6pcEfENFwTc8q6hnidzT
fkBIpdGZ8XZUMr5qP1Nlm3aghirS7Ycg+LOBLMGPi/v7G3Dsw++rvN5qTfv8TBD2C8TZyyzK4ecn
6mGIv/PdhuouayWnkT+EylmrO74bSFeHxkhizSc8kYvD0ZGajy1dMdqg+bIX/4X+EcmlFriUDXAI
+pDRUaPJSLNxk3w0aQKRouxLnu2aR/h+esGHUWNF6mrTSLLSK9nOMY7o7pSiIs+HHubZavNu1gwu
FQ50Dz4uILBrN+ZODw2N5a5uYGaYBAnU+kZhFRD45+F1HXuvaWFtdW3WEOWvQBvjUb+Tw4YGBojg
zOKkld/1dZ4Byt8wycKqpuRzWbuHhevMf+gDMhw7vDTA12WTJQfneeP3VfBX/+aP+8QNJQ+PEnA1
qWVjDl92Bcm8YK7cmUqEhQH+E57cTAg3WOnzjUegKFIEf7wLkLb3/2w7i+6LAsVp6aeSkkYjY+h+
Nyk2NVlwVHxmqdhnmAc483RsvCiAEQJtmGXUcYCWiDZRecx09XMotwtNO4oRBRxRtumd9GkPVCzM
T2PAY272bleRV4DS0RIxI3U3rzABEiX4SwrrGLzaR4S6/MxUpLphN7tfKgJ+vBLYSCMdQ2JrUqNl
8ZD5aQVIQ3E4ZMzWL7avdgmOcBkLrVWnulVaLxXO4myRB9RQkrpNrMM8gniRiVrDJ5oLwfh0+G1S
XSlOV4YjLzYBj1KRubrTG7WXAnGy9K9AyGbzDVU/um0vnqPyu2ahkbnW2GO1X57fOgqufqdP2yl7
OKrLoHCaiZDKVyS/hLX6HMW5XB42GlJUqLTATzPzS+NWuV7+Alo2pA12h1EuF7L/7Z1qw9MxHHuz
M60SOg47pxrjo/S7wkPD5yM3Ff5rHNZeJSm5JF6N+j0SHNOsKKuPiDCCqay5wS+grhpHuivVTvG3
pGRKkzOpeXBl29ELJiH4S9FmWoZ14ZVgOt8Kcq2JkmD4AMkNMzNYNZn02yTPuq3AMz6TySyjgbOc
dUwI6231rXRJgGftj6wkkDy5YdTo6OaGfpfFJOKV3GHwhtmu4pg9VuDfThGYJVnAWnRIz+SU/AeG
bzq2uR25YvPZXVYEXGgF5/A+gUHk2s6lHt5MyWLFq2YZQMvQ+EhkYMGBpEuLmoHM8LFBs2up6T+h
bwoedT1uVKM67truYYT9QNEX02FSudNij3aT7YkGjLe3VZT6LUR6rByxmvNNiRUKFaayrJTdHccB
HlfvYGr/v41H8Hq0KcI4a+xGim+MU3dfHK1Ul0FWFmfvQ9iTB3pkMlWp2/znoOBsucMELQwNoZUq
9PRyFbRF7Sh76saJfmWDXOW7XFnajz3WIGyaeCeo457Y1mBY93YNILmNXeMGWAs1Fa9lD3OUZTzL
Yzdrh4TRKCRcfNLJaaHzpxZlsEMI3779xJmkelmLlFZXGg5RCqb/ItWCMf2Ls5ZAR1GUEPMudoIS
dIM1nkQjTb6HVFpdqojqWIJNsi47sI+F3EOuE+nNo8McpUPrrrV6PFjoKGA05kX1fzFOGm4//+YG
dWiJXFIVvg791WOyZsI1+ubjmBk1zDJWZ28IczewG7ihauCGiu0LxXWDPWNuUIfNTYV2wPoKxPqo
jNia9bL9dtkUYRPtDBTN83M4h5PAKYyeT8GM7N7GpPU9a6wUdg18cN5E0L6RJPJ1MK82SebatpRx
zemIfEG9/J+SlA6wbShCq0c+XWXsJDE++sX0JHrCGcMWWmteFupdI0Eh3/1vie5a9TUb5fbk7d7j
3Dl0KIR3X9ALuTjD1mJD364aGj9674sVaGy10IjFCiaHLpen/X36ka9wpW1BUr7quU+bu1AWL03t
PRdoP6By8QWhcr7n991yi/dllbIR+JqmCt0Lt877P5631dxz3IvNzPZZCfyMvyr1lYGJvH1vTw3o
bFekCElpcSWyonYZEkC2Luux9+7zyGmdmYd99U2QXI960mlOtb/qrPJqBT+l3gdv7/evB69uC18T
vafLqV7Unkj/wuo+gMCwpKjnY+jFBGmL8mmAi4pa+XGRnJnPvRP/1DzMuddZnZHRHylCiuYTNlFP
QZuyVCx/wT6rObb9BEXuFVCWwIiPOlhgrPAEkZvhvn6K4/W4Q1pOv4GdfL639b/urjIybd1IyGvi
KX5mbz03hfFTpPV2uQATB5pb3pYnKhDUFKOIr3cagrx+YzsWrNaE/gdzBlHyN5ivZNxG3/nyiL+z
34YiHDYCAL2496Od9Zl01Sycw2VTpnrukcUMFZggzTlbQ5dfrriPEQv3gCeA1THhPN4gAa5Oenkh
3yjXU7c/87+LgYCxEvPtMJh2uihiThXBPec1emtivBeE/utrsVol+mCmlby+qVkFQG1ifHowX0A3
OzbOlO5XZJmlStGkqFFCSbnGSu9/rtEasvkg9tG+xFpx397mCgd3BhpFwhPgUok6LVhxkOUhoPUy
zLSKR3Cb85lbvyOHCdsz6qBZlj8tXsAwpc0iavLxohWhEbVkUKKunUjdQwlQDGaMuuknfeKw7Dhz
zp6qLdzxVel6ftTVMH0ESPcXtZisnWJ/falavq6t19uOgslQ2ov9m+fdyKy/RDgmcYrH2lyf6NGk
SLznHnO63Kza2Nx9s0VA9qET3V97EuLXf1QnKkiBoO+eV1PoT7FRf+dU6CpB4gj+K1ASvpgouutG
5jErbKYMrdRxuiOaNSdww8AgMCQJBzehmYQyMCjtj3lcDaIKcQ7Hj10R9tmEq0Yj73usBAFbmnd5
hUfRGqBuZZL0Y+m6/zEHzwSKm13zLxFmG8HdxZLfa+/ItX6ak9BhDmulHuCSLIEhmeL5tusmYRBo
uTGCb6lEkdd2C9vuW0xCX8/bF3VOlDWyi4MBKdlYOOGpCJp2aodD6ZHv3lYAldJeeZsyZh2Rkz5h
NvWIqWYfncgvSh4REJFlVyEWw+q+BiYBKw1KJHEnOwiZFiZL4j6GncZoOYp40VNWOC2viYkqQYAX
iWMnWWqfReyFe54ft8vhmkw/y0E2JayUyKRBkBwW2v/0MhaU9GkNG+OCwBU6azFdKdkfs5+DzDDE
BMsLNota1AtgEIKCYN07qmAkd2HdCqXIW5kwyNdLk6su+UvclqlWQYVaDp7B6wRI694H0zvxL1LZ
heaLprsgwvfQTjZz7uq15gz7p1iMgX714Jffj0beiAD9bHyp95VeOxO77amTPJvS7VSstZN3Bv7n
po1cqAz0nK+r0io9xVGi89KZ5vRSmgo5/djWXYM33IHZqgl//sJ6oQHyEUvgDVUHjHN+TBs9YGWd
OknoydZdDY7Cx+EZ4yW1fbjKvdDGUkQRABeIsrrVm2sqskz8pLHyjOwJ2xnCACkZi8HDBAau25SZ
xCWdw//DcHyx8IreMGVxJQsgwb2Kv0jU08ibxR217CRCr9djBn2vdRoKZpFL8VB97fsA37BBxU5I
NkeI35IG5bcXfmFJpHy+/CPWO4BRvjkZJQhJ2QvjS12SAIWM4nuFFJx2lK1sarDG0MWJGqcZ2H8X
ZK700slarkoG+aMrbu9Kn/AK/v6BtLGTPkufNSfT/z+bRi9eqo+eLbtksKl4Cb4lKlUiVpYFheF2
aBSy/miB35aVEQJHSm8tjRlIRkJU+CgZ28ODfSYlU5nx5cmhqjeNm1lD44nvYnTC8L81XcGE+4cC
XBPcgpXBalMqe97V3/EO1aKavjOpPaskhUA31Iitg0lG0PpWii5lrG/yqqn4p8Cti7E019OqMwzt
hXo7PQDzZ3oYor4H0fvrnIHJs2H86NiFDgcG4IDGivJrbOq1vp/C7dX3uf9NBYQtt3u6v4CCvdE/
PD/7wIN+yl389hZ/Ocdid3cNiZJxlCgmRoS1vxnX0qsAPUdGHibs0aZ6HtmTU642i9+i2ge0pPBZ
OCJwnGTcRlQ7Bi/i0LW2U5PoIN10qaC5G94xFNDi9xXCu7RtxRn5BLjsTTDN9cVst6vG3Hl1BTJ/
rAXT3wRLktzHeVMQ1tbEoxvDGFQOX99dVmqzRc9KpaDYQj9T28M11WJemEXxIe3gDcD99PZNSd1r
36jKhoBhhC0ORKl7JyTeK2ot17HY9JBxkx8x1/uknxud9npWqs3XO07Z3LLyuMqvzLShfIQ/oEjZ
ufBOengxH+XeLY5Tw4yabZBS49Soa/1lTeXb8zJViIbrWfJrwVy+Vt8KcnqMsGpPUPMoiPcCJyCn
MddAObz56TW8ALmpn9SydA99lNbCJbHlqDKiBjS6/zd9Rb5zpvN5w+LAtVD9OscfskFmFZDsPm6n
WgLA6f0yDAirm4BxSNBfxaY4ofl3DzdLEHl0y5FVar7Y8SmgXmXFYDi1E0QrsJ6Od1zmSovUUCVH
ZiiQ8Pj7QwFDF9WTWVHT6Z1GQ7SxTlOfbpznJbZ7s1ShHqBojX0yqI5fWlfU+xwSY5hcgXFxGTJt
luqUWle8mdRXN2L1AlafT7Ng4OLmG+2eHKOpq1hlW3vmcHCtln/ttrEu/af0HH9vynfP+y7TFzZg
THxEv0jkQgHESDaiqRF+wY8agCxvez0lYMT1IjugxwPzV3qbBk3ZF2nfBBm8mhPxrCSaAFBcuS/3
KXWRj6C2tUJcaAWWyUeSKH0XDf5Fm4cOqw1fmt7C0IeR81WjTzCJgmQt8g5JMCeh2T24Xs+wTSyf
+3KDc+ECFxFBdH/P5sUMx1xdQHjq6NKV5zoucNCoYp6HTVoAboI0HHRHGRDVIgUK1k09vat/YGM4
2CBgPt8/G7W1dgGcm1b6YHhwyR5H5yZ8jVS2hXrAJ/vTLvQP+U+yB8zelpv0R8ug9DoaYlyNnHU/
t7ry1FktxZGG+BkFwakbMXeHrPjNLmKA/cn+onBfPlr8sWk2FBshWhrqVCL4GhXcP3TalobxIaNX
Lvmixe97W3aNE36fzdWMHoKl/1rrkBpfrq9vwojBWzBaFs+VJy1/cXy75EnKQD5JypxwXaROGATE
0wdmn92KslZYAoF8dTzJkPSiB1R+0z5f43IGyDXc18bLLp2rtsmESgMJrfJgpJifOFymEnGR+bEp
6o1V3ZA8TWGZeyi4FpLeyUc02RwQiMCpOZNa3GFfIZBbxPgi63fosh1dQEWbDdILrwPQ893iW6Vk
AthA5Z4d1ni0lkos9LDEi/skgGpmHTOZ8DeD2jVoRvUCXMs2sxvymKvXR/BtJZlwBAaOcCdoqlec
71eUffXf6yJHzarf+FnXrrruLP6AJyHYDQR+I1JemC0RZOaYo0v1t02vgd8Qbv70cJlB8VzolWvz
ou/wYmJMwHhHWYeChDKyZ7WGNUalipNvzxCNitiRdqmk76riZlr6QGcfoPKNoDcudC9QBXCB+N88
XDypOEPc/+3zsNqJB04/x7hiuEnclJi/dfo5WTYaCs+8RNablsV6owUeWC9eWZ7r5w0ueZFS3TZM
jmz5H+VFHbbPvABC+Kw5+nhDyrwcDApAqn4hnsMCm3vVtArQduGyvNpsX6U8k+jIJf2mGhoOimP1
u2mFZFTasJxznPx7rZIZ+ZKOewKcpr0M6zwMiSJcuLfpfLEButEj3/+15qsVXKVjel/ugg24zLKG
G5jh/Ovk1wj+3D0ps6AW5r1wKLtwCTXPhjmhPfplJ29vCX0Az3YIDvYLElq44pZyrg8Au30hXDJz
MutRyaAp2NGhjaut4P7ULvvQTJ1sdjw8OIbVkDC8HoSSZoQmM2x5llCIcVcqBwn4Ciy2NJpmI8o/
WTQM1d0e7Uv1OEu+Ux4fzX25RX6Rk2ObnfNNQW9Dgoa/f3Y1OLb6I4nNyXE+efO1eOPP0+alQMxp
6L6Qmmp6dw1Rr/pBVH8cOahX0I/vNpv13wPbU79Nvdt1qo7oc/BhU1BxrXAxC9/rp24FMCtFRC29
0k+1J5DEw1+z1EixzpyczH5+O8sLmsAtil3rD9Sd8F/+VoVhgKSTsOnv6hR9DFp2VG3Ubpg7oA9P
IhHCxZm6NGKsB/PuRWdAqnZImqCRGyKErWJ37TsStu5VcFAj3zbUidwX4FzdoMs7DakSfRHs3s4a
d00dSTHKolTggAJnVmmTkfeUxBgQRvhjJD7V3SVaMWma3CxQiVgCF3gR4B3xgTHWAITYIyGYf3BG
VSkMaovecfH4OWB7R1gI4lBC2ih9+2WqPHjAHXiInfuqli3WsmUMdNB9yc4r0PDlacjwnUuiiwEo
ZQGSS+9S67QNUWGXvLcP42tj2rY1FOEW7tUxVqbGeZbSAnDuKBNXMj9c3N4MQj05Ov24V1DbcKcv
tozFbdYUgN0jOGIXppdtDTznKeuWon6hCLL5Gy/YvGkXI03hkLTitsfR8UH6ybWORS76tR1wL2UN
ZYMklVCFj7ZAZFTXBCIsBQOS3Jc1lqo4yyGSMMqpEwNXHzsk+KTDgf/ejMhHyZHxnH3DwNqg+oRZ
18rQwsKzPwrI9be2+2cxKUpMezrgiKBXQyFEOwNsc9VBSMPqRw8iolBs7YHxfqZgrXx13/xXFfB9
G0dW4g1heBgaq+IkK7g1Bz7HwBV8Hsalipmw3TG1SNCktgrseygsEb7KBC3Lm7u4Z0SCJ2eOst0r
cgIP9y8FzxF60lgQM0NP+CIRfoNlA+SggftY/bpIgh8gHl+MWjfFdJze/5B9ocbuH4ALtF2AToTp
Oyt/jD2K+rns8pn6C50zF0WzNrVCdGD1MYpnTGmLsaDUaPhUjJZq3eq5Wl5XT7hTfXq1KD3bORxQ
oFgPVQ1o15YFY5dr+3zMvO7oOLalA5FH2+b+QgqpANRM16KBhGhH51AmUrQfSTeamoDIVMr8k1iu
bImuBYrtJvT7bdsEUG9IBYBQ4NvB9nXCUtaXhUIGMTkW6RSSDN0SSuiOMx5PD3TjsuinBWqY/H1D
+jb79OdnbsvcFd8KNoqgZ7boDZcRr84IL24VgLjQSrxAiDkGvUdciT7fGONqmfx1uhBeRv1KLJ9n
cJqnHq5ZnMVSXjIBdSb7Y6BkmX6mraYbcqFafOQhCuKh7nI9gs0Y7zlnDHx2JcdTp1qBO3UUkj8+
FjeKS+ZDekoJuUVr+0qfTh3v2b9WjUn4hUBLbbDFGLqPytWj0/KGgzhHH0a9yrMtG6yEA63/BGei
+o38G5ZqASZLE4JqIWGxD8SlWvuclzgeEsPJZC8lostin3rKmGU14s1xQS0tPbrVc6TbE3rpKYzl
G/qE9XES29Lv32ImfF1QfZCVzTL5oiKD31NV6B2GugMFkHKZZ3uSP8nBkWRLoO5jyzgk4Yv7ohgk
B9HlKtiXLHLBoG+vUDsQMAgU03X+IYX8/8pyXTlb7no6cH1FHAUjnsVYQxyBQED07MIWHrNxPkQr
k0XrMoohQb1CMzuEKAnzXkLC3jnaF3QmHo9QisJgATxcwrh/vGPVkzmepucD5LdClb9NQv3vIbpa
lwQiwyJcyH7rI4e0hiyzJAK7oNFCsRwG9CSV13aQfdeetGN15SCFT2GjceRI87J0zdEF4jLBI6xO
AAAyozui42JGsWJl4gIqkGpsQAFUY0AgGP3JNWPojKT3ugRR9+wuwKkLC3VIhopleeqaV6wxRL3h
D16a0E+IgQggyiV6NaXbxmbkJxMtIGIT7PbTFt/MzP4PbEzFvOgA0B/9Gut8Rb2DosJzUaGz+K9f
E2I6/17fbmjeIFAHXleGXxfpeqD+FO5w3HHDzrjYzb+/YQimYQfcwwtNfoomo9DCROMdEJcMUbwF
bnTufTRW37r3lcl1v8zbG8/9sMUOOu+A1+DCeKtp6GqTDGvgrUk7QdsC8InDhFTiLiyZWt5U3Lc/
5aD0IR7ksnu+cbt2sRrJ/4k3M2ATrTp/Y5Jzd57vvS5G/n9ddD7w3HR64F9MzyJoqzS1dsN7vKD9
lm35sjkAu7E9OaLk5HeieRcvtDVcjaSiPTzNd7fN2LkTtwaoSwFDH6f0yLEItVCrutrvYiJVDV+U
M23+AO1380h0WgKJbg4HTZ2B+U3uvrN/iptsnd0w5TNUlRqwjhS79Ocgv154Sp9YAMLDNnzEpgey
HWiRgoJp9GzF16YZbn8C7cApaeb8zGwwijwwfJg6eMa7p5139V58d3p8GpC8roc+EUaJiAgNfl0b
qiQvJIsjLwAGXfkU+huIs9gjqCc3ceQpGHbgxp7bJ3NDcqEH50v6+3IQdQpeyPQtFNKMS+wWYsFa
5dFHRGSUauhsnaphuyYqYkUMmZB4+wTUGgWuPf/2BI1Nx5EJhY29ATmEi9WPzMpAf7Uzgt1JXMb+
okxJGXlXFItYRZSHgVPEtv09YdD76MtFn3lQooCnNG4VPFPdzKhuaqZOKHe4PFS0Yg1QY5x9ckuF
SVfPAeU+9dL/y5+CtpdZzF3V/vuIjbLZ15L32iJnkhZDD6Stu44BzJf4Nx+f52QoGZtV75XYT+qZ
uUyrj1S5z6zTlp7oCQzglIH2a4BgbnlaGaC5wP/re0bWurcpjxkiYEgVu09VMydXr0xZ9iWubg2d
mz+HTkwMNFfMncHuC468zu/Dt4xNz16e4ODXwrBZa0c/yWPB8WF+fhNpHJmFt5w8uf8cXd5n9un4
8fGJheEjxiOXhX6rKJ0jJXpRQg9OAze1RUdsDjUwuuM/Oc64rV8JnQM0E3f4umuVW2U3Jv0hdqo1
pk3U71eAcEBcokIY9xTdqLWttVZ/XIR6PaeNvoxz4DmsuvjbCRQf/QgQSsF8iTwWAJkMvH+mrK20
TT1C+h/yga12qMv1HoGtDQFVkZ3AOE9BgUEfCG66w6YVLRm8yNefao9QNfJxFGaXYBm7mFjg81Hd
UfqLwPrcMmt6Jqw9/pk6O5R7GIeECWfJnuPufzzICPFlmQ0IcUeAtr/qybkcQ9asuqzH5B2l6Xbk
jNeX/PGnl4mFojLlW0QVB7TGpiWAmA3m9jVOiCaNi8fw7rlqVkpMxXN9OVkllrx3VwWvgllcGWEv
aG+pw+JWX8sunlqBqoeQLDtkgQLc7f9kPqT2uqF/eD1IObWyw4KRArkjxkzXaQGnq26o/D13mdLx
8ry0aVQR+5Z7onQ2cdmxtjbzMq/q4m6qXebisfxZqbMxkdCCfJ0pxWCZf9FfvV3gcf2Po7E8Byab
FAe+YZRoW1wOuWoVmjXBMfswGWm6PaKlDe9hkXxdkf53iMnyqvIVgAOY2LwqW9T9WUcpTeu054ui
TTlHjzwTr12nKiVKssjbGMJqCqynK125omLlLHl9YxlB5USWkdXFNdexi08c4CfkVtcSQiOkrJRp
fE9QwyZfA9UzxyMNL5WLGJDiHZUMsE0oEb8ZrAofKq+1gR0Bhd6u8iCEWe6SvUNyP9OUGaGKnpy9
StquFLR3Lm/WUbNELzx0zvwxyptX6lNukRpaMidgL5D73UD+YeJRrK41dkxAsLALqVxT25wnE9zc
fuuQZva08R9mtxzu1+Xg3wf4sv9CPOexK7ImTOjjZDpEp6SifObki6DFPxNB4ulZh+un25irM1t2
tBw6ECGho1dxUyIWc94eYtv1WZofqHnBH1EQ0N797AS50kvi0AFifphn04olG59Es6UnR8r6kVWt
5W6CmwI3wzdg2my7VzwWxmJDWJlld0LKZDnJSo673rHi/trZR/Y3Bfth2yFqhOoBc3eDeuks/A6p
LwgLzAMAtn3hNG9oYghcFzJ8zl81QvtNsdmN59L32XEIOE84MDiVHJN5lQl55FWfKVwxn9xldqOf
LqA54yKY5zCTYAzIQlVKlQyGppzAoiX10IBAtmRzyxMViqWtpJ6QzQ8IzllvMn3kWh2/Y79mRL9f
B6xQcr5od8hUk+kQMGdqiRxEwRWndv+573D6JAAMXerMlaQRacJ8mGbgqQkyYSiGR/LEPbAvg/zU
eu1LDQeYU4h8LdiWlyv4uu4olyu60nuLIEhK8whWvcLqhChS3QrUR2TetzdsuomKeZ9DVRXDn1Xx
6NCou8uRo2weOLxWhxJ6cz957YI+/+YMxyFB9t+xnqnXYb7bMRaMOttDxzaf58GtpZcEo8v6cCYc
NNGsC7Ewrs47CX5IYwcZI8mfaQHHEaKrFFyfuNHC96yqe1/liCfPyLyhXoOeyJjGZNL6D0SwQ7Qu
5pTsdyDfupqcc3cDBL5UCK4xT2rDQQXhEax9yup1iKjxBCUPuNIDidDQIiTIvBnITXOlk6WoA3Hc
ESMvS5c/JCM4L6t5rsCHiqmExuJ0HkNAIq/u7K3/H9dLDbpj9y94gFfIllM3w7pIRyTEz7Gyluei
1SdEBtQLYGlmo+utBgKMAoy6z3e442rI4Pyj/NwrDZqzZ8rkzm3/ilgY/VJVPhkhQV9J9vwOnh2U
wGgZJ9KlPOZISHld8LwnEu/e44aXcuqfsdQ26Nk3ygC57gMxh1glJcXAo5wkF1zpExxSgRuLbg2n
uGaSSvQCMBDfUoe5n9S9ULWvIXVyqFNkgytbbFcPyURDk57aO/j2WOl+dxCm/Ka2947YL8Su21Wf
CVibrQEqCmGQS/zMzebMoRs3P4X1/A0hHR1giEMynoNTsUB+WTrioWTXToo0N+x1MsEe0XyhtKoj
v5Y4MUZTpMn7GHpagbGrqMbRy2FWg3Ia7PtzweglPAiwlr3PtyO2K9f1AoGpXxli09sSwin89ibN
s4W7TG8LWISJTMbZ/A9I10kG/1ajQkgL0s4P0zTDG5iZNYg5iI5NvHXGzYPa9UTuneL5mguJnniN
8UU0kpXT7ZZPjRwZwEs3ZEBYjf+3AKXuqSheHctUXKE6rXOHqF5DrGGRr8KeUKLYh91fqfWC+vH7
HX1usotcUZN5R9/RwNC5TSJ/GazGBs5ygHwD1+u8V/RiSlqbANSXcRrWJjFQV3IlPyfD4JPYuGBa
lkZeTvnEb5TpuNfQj4/6QxS/Z3EYBcR97S28P0zgPRiqfiSoJFrnuCb0U2tTkpw6Av8f0wck07p6
qNCchREbAuAC6O0t9CHOJhciKCh9O1EhskxlV0NqPbAgwjm06XTD1sBJWZsknmOmhsL9/NUWJRua
ak/zadyoOrXOUU87vq2etWmOiuuh7uc1R8xfTJW9pF5aOC1FQ9p/5BXKbJE8j+hjYs6cukNwylZz
tMVvRw+BSVf6dcCfqTRqUUzq00rjEYjgKKlQg0M43RyZ+H9PzSUWt+jmLwOER39/+fcnTNOmOK/H
GrjizXjSOMkpBRe81i0OyFkM5N2Wx+YgwCS8OM8S7Rr1HQ35DXpDvKQOV1j7ArcCbDi4jMW3PJQ9
DMZ5jThfruKP+PnRjECcjmXXUglZ71k3Kknvry7N04GtdoF9szhh8d7G/HYFnoRnvHl1CqZO5lad
9S6OAx/YRaz8VurJQL+Xjwwc8+JI+PxDhx0781IM/Wwq+q7awWlpYodiLzGRS9t6YLr+mDXu/DyH
e24W8Sfudfom1s0iHuOThPKaV0LeimKIyhmAiNtBXnHTv/6cOevEp1Ev2Rc33ozQaQGqrOq6pDyR
2exIAuSDH/BotafzMk1p3V85ssHNt8B4yBNWeGjnkRTYvKr2l0Wi4HHQKF1jtSsbarJxFctHx55l
gyVJ2JGON92jlOPH+DotRSK0bRNmFHWPv75ILR4jifRgV1pAnQQQaApHK4+7PD9QQ6RycuvpQtYh
tTTtqs6WQxGKuyT22bXH1MEJeay4SH8iqP2Oybv9p8QT3Q/ZcxfbI6R3qrb72u8hMq7Z5P6i0+/X
Tp561n/k2xEohyo36JSMmn7Q9OnDm0+2erO6XHpSW6cjC8GxVnuRE4r77zqe5k94S5WJho2jHJ3u
ZzAQ0Only3KV+MZ6jZYDT3cd9fJK8S3vm7rP//kzo997QMURR8oW3wrhXAMIj4LfkTR5NvZpqBBz
ShFTOdyivG+ka1bBkd8VF0xgzD76IFz4ABXtLwk7IZbd5zrHugCS/e450obcKFHJN0MEhrFdKV7f
fsbJ2/we/KXK5vox503HDOMSS5WemrgRqGFnbZ08BH+HFlea8ByCwVxQxsEx/wBf2gE3QnqYOwU1
SG4GtAJ1L3oUGjpxWcOrJSvxMCofgXTqBluoJdUe3Q1ULH4tMrcBJXnBKV48jHxWk1HpR51SOKjL
nSuVP4nDGt60CpxkCmWyuJz91pFBekjksGzPebADv8KmJceZKww2cQOdoz1J7uh1SQ6zEeFN+Hoj
BgE7nUrWcc4FhYOslW+5bf4k0DH/IMIL5Jh6u1SeA6HTlUVZN+btIszQGHwZkA/B8bpemMHEO2mO
dgCyGgiJALQFJQacJXSJRVPQQ0++6wDEahtkpu/hrsltT15b3BusaOiyCGz38A5GfUALraBDdqbZ
95+HI4EueuCVBiZpg+irwccxaZKfG5gwHiERZvN8XYoswlT5+DlR9YI7fcaLkJBXff8v4qoz0Z9/
YseAMJ+i2sb1f43oXy2ktEXxMp+t8pQVkOwNxhYs6QqH9Tq2hS17TaejwB5UMU+C+1aQidp1KtEN
PKJlED/823ToaTxNFnGHEq02Io922f1lQltrh2ylxAmwPFAjm1rQfSZVtysy+pt+ErMuAIafzQ3O
PH7D9vV8HwHQjwbXOSMnwRVGHlSUZahjJkSOva0jr0gJSaIjpZuRf3iHDQUbs7b6VGmT0M7BHvJ1
kQsuLvYx2LlaxCpazlkxzZx4j495w2aoCx6SxkC8DMwNmEI9B7Ob5mWIAhPU01dRnMhqM6Xm+AP1
xQtQa0z6jGib5lpTLM1Wp71JOUA7QvqRLdYlWc8I9utzRBJErEjR21wVVQ1j0eFNSwfG68nHtQvn
FysGpBsSD2dhGDa5IS17r4T9UL6MGrMs1k1KJ0qIH6NVMUJ7wsBeaW0PrY2EKjgswv4LfusvTcxY
ra9s6QudzU8sjTlxvB1oGgOhEzHASVG+YKVXlxQPdUefBAZJvGnYTZxsPCrmKTJwhvUK6Dv/2Lkt
3mkDekVeUzGPiSxwt+8zkeC05RxXHBRANbOgtkmKtLshB1XsoLDUDQykgT5CKmBkoJlM4WrWkIqG
QNRXEzcTJsA4Lpls/tghRwoEmfC0C9KtIi70IAFp/lpk7T2PS8ClHN2LK/A4xv+/I+nn0MCwev/M
OtMQfgYM0279KAAVLD9AmNi5mzNnxaPGb5NxXk2hlJTu2hPnpCueZtmyIN4Xwd1JdJHbWpUYr02/
YUUUUp3EKVmLnMNWn40Q8I0svoO4RjHXYWGYl4bAjLG/5pPxX4xRY2xF6xLX1rzsKoKXOTcTzDc8
lrbfZMVIdC766CHt2r4UYsw9SBQAO1Ip4eTNeTyYOrRbYsk3tsmt4oREjaQqxzNVu51BIkqNnz6b
YXfZqqBlDQjt5BOXGv6rWRdoLlkT9Vi8UtB4q4AAp56mz0mJh64aJ8ECsNfqcAP+NP9vlHbAOWdf
kFZF4Ho8fA0pt3rrks9tjAqCOeBDNQJNlceKMO66ztYrYVxw+q05fhzOEUe/eFJR3k2Oh+rgkHVD
t3ioERiHvvF2x1uGdTmyDod5AuIDZsIdcY9R6A+9DD5R4O9TtzRhcVhT6Fj6w2f3eJMbJ7hgGFSu
gJVyE0k/oBUtaZDFIgQvUfO8h80pygmUQjv3rBsjXa4FBFYSeKjpEdfgGjoZR/Xvhk0oBnwT4/i3
JiyHblZMTxMFUAVriLCAarfy9G6bG5NSfMnen7K+gVFS71ySG+dh82RMew52NPlzyymRaUupxZKG
OZhy8iW1CeJrg7VWNhmut0VB8EzxcOWLx9QWbipX+64PhRnRb0lEUzrLtS65e07CEPpiSbNT/pw9
UIYiCgdqqgF4NLXdTYDO+c5UDySNDBtxMp5a3Pvo1F6CweuYgR/oM7++4/9GS1NExtHdbom394Lf
m9jyzQ4XMGzw3HZaW887zcxY8rDMqmoS0o0dIdipFJjM4j2HJkhaaNMPsa5US9gfpDwiP59eNQuJ
8vUfTgXgqOriIywV2arlxpo85Eat3pggf+jmXq8wZYVEOvZA9ncZvSc2yf8Lrj0VZAAj2sHVIQAz
dcTDdUtaPeVpZ4roz/xHi1Gx43LBcoyIXsZnYcFYx/l+s67CMaLKimPV2j9KlFx8corVE5aF6vUm
KlQiAvlRwg7lTn0B6RpCX52cnmnRSTh/2xN4WEpH9IrQQk8qYmzFq8ydNeGnvMu6hVEYAptyZOW7
06jATkUD/1VixgZTsCmmXrX19NYpv6Dlrk+fJdcax/eDbv9usQ8xsqRlDKMVuHrVZRFSsd+3xuFF
spZ5r/OISzyjCp8bi0o9ucgkbWxh8ZcQo9GYsvaaI7lFvXzPVN8yFIH5lS0vwfK+9Wxvn16mL6QV
lF8oVcr+kryxL6JZ2LNFM3WL0N8U5amk/AwudNKzfi0kRX4ztvIANx400kj+PzbaOqzg3/M5hOwv
7Ox6P7ISNogB6pOsWVvjR6lFNha1HD9X2/XpCcaitbN62HG8oR+qmSrY2OKb+USkVp7oNEyZVQGF
/krD6zWNiKib2Rr5vQsngewhPQtP/73RDCqHlilA7kHyxvUnJOhR0AoMGRKzO0pJOrTPu8b0enYC
Q6Cm+744wYJ2pHOwPsQxmRYVNw/Z2tpWluIJb+imSRM8OfvZo9L2oytDDWbtgbz2nmUeKu9Wt/xt
1i21pdRZOTgoRhv8hV5l7EF3XCF2itkyMFjD3ED+tQeNPpFWxeAixHdU24aTLlCJu1KRdeRvH/5c
hoCaKCj58gg/LhfUBS603MYskYGtEJNPk7fnr52TkzPH97I5iR4Nui+BVSu2IkfW/sSfczmudFDj
NGzsytFG8KnEQxdYdleV3bBx02L1qD2BpEXVIr6EnJiBnhaYvVLlnTm8Hsq51ZhnhOm47TOgKwZP
aVni5AvORIJdeBHeqEZxdwCIB6GKQTpN34AczLw9y6usycOnTlVDWSPPNA/fKz12ZU99XarJB/Dp
sXhkupeyv3ai+nAb7FjnXrZdAZUUHnAQz3gS+UEd8EOlf18WQMszgtqkomQNMncsCyv3WOAS4uA4
Gu0VYgaWfWPeR1d+w5SZgoyHv5iOB5TZ3XuWdJIphS2BqBnDU6GeBHEBZCp6DmILGQYxezcYxPIY
BGpjSTrvRLiCPav8ek4QyXL3TAcQieqG7j8HJcP3oZBAU/MWv0A2YKysAHer/t8OXREReWHPLXql
2XA5LUeT8l8a3iLJl7ssJZoVBWbXoTdnKJaM7fVD6KuCeqg68xlfeXzGXDl+zNMTsg0ht0zbmzIs
fbNTfQiyL881qY53PtclKWZx0cGaNNIL523vqUfVnElXq9IW2mZK+Dds4v9s9CMfqF6T4VsgrcEu
peCDMGEHxVETPTbFAyxtACKPHlhB4Oe2tpTdwRk4ximlZsKTWmfRAhRQEGtgWQptdEvXDoaYd0Hi
rHzKx5+V5D8d9O+CVGGJIQFhyNe3apUww0C049VvVzifgR/i9+agtSGPtDGN1wqqv+IDL+AhmC79
j//zHChW/JVB4Jb/5rhMs/rQWtgDqMKXO1HYCegbwTv/CMb7Ft3gQnOdw/KtOAbFPK5cBwPN1/hL
qN+eO4w9mf0m+lfBLcu4LG20Y5RjkXW0FFGUwVzgQq0llBh7QIAzBZs1dbieHGna/kzNrW+wV9IM
flHrAd51uVtk7J+faL/1SQDu7qp1RnZW2F4A+Q9T5BRjGJUI7IuEWew2Fz5swmAgeRGIey4sJtC0
DmLIVrbu5y8gz3iPgNJbj3S3ihqmzzMOKieV7iT6vEzeZ4Dm7d+txp/fZn8VsFwoKo1MkoeW4jdL
+6T5/XHlEIEKyaRucfSZh4UkEKFmlpDQ635ByQP+hkoXrUd8LAaMp8dKhHtXHt3VcAHwpwmmZKGi
d9ijYP3fBxWHeHXuW9nkpIcah752fVXljURHFqGuAL4rNXBwwHFAGV4enzSRzph/0UhmjcjtWUS2
7j6nJIEwc+ef7umJUYxBrZWuhx0TaZE84jizUN/o7MfvbSSR4o8rRZhBjc2CmnRsZus5bk2Aj91h
oQSSY3dpaoS8uUPbpMR22QN0YkGQrq+70f9xD89wxSnVQ4xxakSD03CN7sn/ry5xXamMPSlUrTBF
QPQBa+W7r6VX7jZMHzApfwdqmhFatFOVmNyILrI+bCn08wtpUqX6RALIx4q7qGPbbpaDX32AARHM
Z/QCFvjlrmzPD51jE3o2UgZYhiEfkHyae2og3HtUKv0q03u/4btFFPJ0Gv1FXOcFMxwdvGe3c2Uk
4OjBIiBVeZMc//4EMSlhqSN8y5jJTLdSypEq37gOP+HiL9u2hIlayX18ZDiIgTlm1hgeAxqH7i1W
5Fycg+kSynjz1d49EDRJ8DitZBRhTnXyzM3M2nHsRlqcz5wYAz4O1sCNwZ04YNFu9tIMg5RG4GhI
I7lMVdEFY0xFVfbXwQtCLrFUBIP/nZn4GdM4St0AEHT9Faz1FcS3fQ5Ff/rOfiZUZl/ypeUNu9od
6izlBtdB9oE++zY991a+UOdqVzpOBktbWUMXK4SvZz/MIzO8n2g9ANEbMhqi/V2iJZCZ1AvW23al
/uoX7oAHzkGDp+0B2r19iA0LcWXZI9/7LTPGQuofV5eAcgL2zR1Fahrri/MP7gsQSMipn77brOOc
Q0REM5bQJvmgUs9PcPZO7PW639JWaNsGtSIyh1UvPPM2VAgJV4pWcRPkDye8s9I5vr/jUTXRPqXS
tjlJuNIUa07Lifi+s3r2kJU/hFAcLO2NVrB9GR4jVHA7SdZBZoU96GDacvwFEVfmtirgdt0rjWgS
Zss+5vqcBqaAPZyBRY5xOOencBbFrWPLFvnAYoxBDiyfq6Q7Pq4lfLHaWm0Qtsvld4EppCRUcM7q
MyEYaBGcqZtRaRK3sRwFgVfjE+Z7F+QFDmu3zR+aMkthPTbZWeI4RLrvP9qPYBbQTJnJXU1CkegO
LuQY4VBtBrdETZRm/1Ek0GHqojDifHh14k5m2EPLRhSar0ZvuF7r+Z5/akDafek7NVyjFwV1uRy+
L1TWPxo2+AzkDtX4g9ak2wCDRXk5uG0AmMjQVeXPaozpGc/xg5mAhrAib9Q5ZAo6Ul4FKjTriFB2
2UbrlJbreH2NLHH15gcZhnEJ/GsJtRrZVOqtugduMXoR53CenFsO+Wu51jX1Oe+N0Soo3lMBBYhB
np0fI9RY28ItLcZm/ov/udVK8q9o9qsf+w9vCLGhpdWdb9ic5Gxo+11zyGC+OM5FQnK3nKetmZh7
R/b4HTeLZaCi2I1lCzIjoF/JEFX96u/471YMRiCYmqpooA8E7oo1Usc1v7owQRfjxvtxsvKBVKRD
dfWb3rNuuovLknCUwdk8Ogt5i225lFTvlTZ32uE0gVcPnD4MigsvF56pZr88enfmkHlAmq7VPxFc
X23rHHLQbPTdcgPlOE5EbhECSysY70LI+zFgS85ws2CRrKOqUMIvsAE1LvXGgRRfiJL4BVElF8ks
5GIndze/+HTdbVBhQox5IiTJc+XIgdrTuv/LCvdTcl545JiggOVB13GWHT8/HOPyZUpdFa40ZqyI
oEHuQkBMbmoC1IL3hTH77gCpKBG4f7PW7GEqLWHYGSgUPB7ctDfz351ePjOwjRKTtErMoEuz1rEp
TRHwPk74zdcCd/+N3CQW4/Lt1YOzrmy1t595kV0QKi3IQEf16cDYWKn0J7271gSmFABftufmO39u
DTgMLXvCekJxp2gyix0oaip8igq1EzAr+0hUw1ooexxgZk4lvYsgchHrEOGDMpX+IUKBXijvdAcI
anZHENgAJko80t0vcZCcS7NJF0JspX2NPQge8V1KJ2ubUY9i8Ai1XNSyyDeEoE7FtnqimNyoo4Md
oYHsmkoCUmQvUt8h9p0KFOAVA/XY2MqsvWFSEVKBztbkTE2rVH/zFE8+JDieRrZ7ZDy8otngYJOY
2tGhzFUkNTmG6XcM02zsm5Sk6EAGfKvRaGqvgMWjxhXF2wBnukGbHySFlGavR2gEQYVwRwceDgQA
Gytv0sAfsIMgdIV+4WK3y+Aoa/GdvhfP59Wqn88goN0iRCXCk2AQLy2KDvDNV2BA/25S0DWt22lr
xQ7D4AY1DKcb6zJciAftzSSEdQHA2nwEDA2BduNrl15HtgLqNclIBF+55B3SCHU+mEGprs49grR5
AtLCAKyVJA555hXI2YD47DOhRBppQ1I1rVhI9bdsvG9yYGDlmB6v8fmj5zLZHbPNOmWQPYkAsa8h
k4XlccD39YYGKGdtqCnKQzILtfRRtjLbenrwq5HxfDLg0MLONynKmMQm1/EXLNw2ya20WddztpNv
f4Biyi8A5gxijvwDRYLwlK2zDxf3MH3wFRa8/xD9ebDjWR1JxdPzLK2MZEU/pg96ax9rSSEBPqNU
IQuboY0hcz5VLHAF7eEMoY5Zh9Qrym2qk1lG9JN8gcOm36IgxE2kPMgrfDKbifNhDBVmHI8Y+XJU
FE1WRuBofkNewNLYcbYSWxG6gYtIpwZwnu6eGo5wRMUNcxFbiWfbH8hvU/KmQPp4dsLF+hsYUH+V
WZ7nTep6obBC1PvqWdlovx8n9C4F4gSS3Aih9ic8Lcbf5F09KjWPvRk2VIO58GIlmi2i3uBAk3Qa
uS3T253b0vHaOrgboPtYbjubwfV0TfTa6W5rw5haEzuh1BrBCu11JeWQ60OO54g2M87YfePk3RZG
jqIQtaOjG64nHlUuGRnva+uaYz7qZJrp1HM8VSrfU6mD/98JSnOkQce6oBURvqxywBxeLcbYYJXA
hrlaXFa+w1YhJ7nK5vqqiJuk2bJuMtewmWVnyQXv2/92NYLfpIzmYfWFoJKPfDke1wHP5pu532O2
LP/5+ptRI1UZlKRjJelurI3+PgZEMqfwMEHdjBtb+yq+NNt20l5ozb6BJoyiTS82XAfbdyD/X+Ka
T0sbsqkgL/E+QZvV76cnLA46B5wViugs9tjKteX1Oj3U9eSZEdaKOa+W/NvtsqBhE2cqMEPQJ1vO
98UfQnZm70yDMwxvhgEw3CMgGsrvl+AMUzUVomltvMA/kxcF1tWCndK7WT/UZtBD/kr5dzZ7QRmq
27tSOQWRKmE1b8xMQcC2o8xn7ybjX1cI5Qx9JxxmQjII21DlTbbGnie8Yf0TyrcgY7lzp5kHBT0J
UPiz6ZldaOYkjSNwdrxq+7tC0FRXtdLXzX/+YrTDlTdVyR+U7SVmAZGwFnjp2dvZ45FWcX1Y6OmA
fa5va6Q6tVU1OXAkqDIKMBZeC55w7c1tOUcIWDGe+lt7EBd9rtPwiu5TorPY/FJyDDpC1p1puEIR
X1Kx00seMVHwVuriPRRdsfgLKqMHq0s4YNOx1F4qp9Gk5Y8fCWZb+LZLTu9BOCV8d4yZIHzX5/Ot
/4m8J4ksIwA/IAmAwbKg7Q/3R7i5VO5G09nBWeGDd1G7etOmaMEjUet6Zftd0D2boeGMYXuZ+GND
eRTsiR3YkUo6eVKOUi9FhVy1zY6dIBXvXRNe+wPAzRXz9xQB38L2JI9iu0yHFVw/jXbYgmarzwRq
/MZ/NEivyD9zCKFR8kk0qP0uK0zeBKm1SRg+PknsnjNn2QO9sFn/Wm4cRwWtti+N+2Ktku7FxSil
GwfJmghF+bp6NrfFY2nkgmSpPbIo0CfzZfv/eXuDKbmqWmEolBrQDbQoV96mrYFJnbymJlMH7QbJ
vs9rK4A9JeIUrvsP4gjagKyxhX7cDR6STF6H2BmfE6vefoSFiI6FecmVciPCIePFkTBKe2CtuXw3
Mp0RFoIkWUqpfS5vno4OT5XI+WeP9yKbWAOU6n35g5XUkFdFcCmvpgWGa7XJjy+Ydrxk/9++IhEa
z+DwOdAU1qWQybdwQ+kAX17LqMZJ63Sd3Eb5VXRemscQs+2IsaRV6EXE6vDDHFDE0We0GH8Jw+6X
MwHJHCyZAIBKLf14RfOzxBPBAoF+REdJEmDJpdb6eSiqQtMp/uGLw4h49aojkso3ekvFM0Tahx49
2CTSDBrnN5EsnjyuzfBOrGwhBP5YTKy4x1fqPi9qwWzoQauPzvcDnxd2ZE1SnPEG9hHNgLBzLLXd
xp3J7EiaWN0+MVzUF9II9h32Ly/gJ4LN9M/5Gz7mTKqmDoar1w+LYB7x8tzKxU/ZAV5Rbcfnvl+i
Wu6iRvHY8T41vYDWVfJBlUpMdFoafpozL1QWoCeuEAqETLdxk9mvxocEnsWPQs8o/Lyz0saOx/Vn
sHSOIXc3HuW5RYkiz9887EjquAgwv3go1pT9krBFHkRi3KKPcCQllYtMhG7xPV1/2gD7Mc+/qMyX
qoSMj/w2HLe3TSHaBoDeoya8Qki0UV9VzwjqKddlN1tOPgLmL/+qLMY1DOIPFjcswWce7nDGIduO
d3SZOSZF9wC82xU7MgB24hOUFQm2j5wTyoLL+MX4KJS8vQQCoCreD5GJOXaOdRneQrHEe9cyoqQx
CJS2fkL39Pg7/6ArbAhQwh/bOWTsuEb0ujbMDEODtUnjWgPhGvRQe2bPnbuaauFUBpTwmqmGsqll
giWkAKUEwjq4EqCjtEYmCODBhYeGxvvU4aHChaMkKSVvdfo76TJM0otCgFiFo2f8mmEyRa2616be
PPg9bj0jYvHhBRsJFgZZfjwUo4DxZxJd4fazb9ptWjgPDsZ7KjBUjA1WohLxbNlu2AbtgtGGri7o
DXV12Q2rez83/+44WwOWM+95GS1qbQNffP09laJLBxhfw5RA7oI2vZq1uzfjxvwfXaU+V9aQm5Aj
JEa5mv6wAtA7PqpxX8i8NbXfKXPQFVcNv6lBreaZ5+qm2427PRn+HKTASOgyIh0DQ6sNa0P6Wlgl
o4t0nZ6Yj1qkBA3PaqZqC0sJs6HSXZmNNMCwPp2Z4I5bxd74xW0sYhcDffAabLxCvybTq/kJDXsz
CVeonZmKuF9p8SoL5otCarA0zY1DsIMo6l28Gu9exIJkHv9CapSanjip+dlKa10Ub3YAJKI3NEQV
DU3lFxfWsRKC3ZDIEpjbv8DZucT8IH0wwjDVSmm62RS9ekCrgSD7DTan1DH12AS/wm25NKqpYbry
tJgOkiXuM/C39gzoJjRgdGu03vKeYqY2RrQcya0Nhzf0l7/Ae4iwY9eGDA082fDp8qJrVsbU5rSd
gzaDNdx6AMB2xhJoNWzN1tQ01VYDCW8yduY+oToIhrQiXH7ExtSeqJO8iykpuIGnN98LE/yglPJd
sGRtIGv7kCpSZU0Jy0S9serFsI8BLTCWQ10DEPc7xiQWMziG7OmZpi6tfcY0s/JOKTNZBMzGEUqZ
7SccptXqJvIHyOrH8hfg3aLp8XIFtPYNhHv09alxLjmpwJkV7MP7D9o+EKf4ptxXFZ+BszckHnts
skhGqyJ8lPhcLi6oObjNvMu2HuAOwZzBruSRlX/22zxezfynsiCWt1IMeoAfMSn8lO+8Ge1k5d7H
OUfXULL7zMDN1/l9h/55qbBiv3oK1KliPvjKb8ol8boNdNxiClfjLhS3D0wLau9I458tM+Q4bQ4a
fznMNyGgUs/K37+0tqXk10xSRvRN23gEP/DaQOZBSoGT9kCnBuKhV2vyxVO+BI+knZcJ7+MM1oyZ
ylK0lYjPsYQTOI42vRM0sC4xJss2V0ZImKRo/fjp24YHrR8fPf3F3PCcms5CoOWOR2nDbpHV8ypp
mwfNrnUVemHANEbKb+c4vBmCeRkwE3cm+fGLu+1Rh8Jtia52o5iqGbK5c5AlrWPlPymM40Mk5bQq
NZuKW7evu+taSONFlWFbxsgq+xPOQF2S5xzSUnkjwqBrUOMErlBqqMO3z6taLy8Xd7e6ELvhgrGI
112xFLl52q6++WXWXQYHc9O/fRzpuqcasNZjry9CyLQVhwK/G/McQu+Yki8Fc0oKeKqk2xhRmpCT
gbLhNZ/M6K8YkKXwa2ailG1UmHgo23uUbUFp4v7w6MMgSeVcPglsik5+ESRm1aCcu8FpClOT3r5T
xGfJHt5OmQoUoyVgLA0noVg+Yo7u7aNzKeaCpzLMSwZsoovAckvJ78afcUEUrgfFoVzXFo/NUekf
exda1bpKZb2fkJwVzevN+cNL/dsKwlLcqK7bsQADzahDwQQBjLKWyESH5VVGD+uUwARk+zCE//7V
dxKVKWmVVTQxtnDdMYpyTxTzzKJgoOBFrWCWTriJJH+jvKfjMZqDAEg02eVusSHseXUamfW+MQrx
S+J8YFMpM3jcPCW5vy9+INQt/s6fQtrn86n9cRuS0sU9bCPKGPbvxLbM/Qd+O9xAM9vpXekOibYF
oBAJbNbpEdea9uIzHRM/bouMafpOnUBcp+l4pDCIjjt0pZaFoRAJCybftNYheRANtOwY7wyULooW
ILzmDh9vIgV7YhoorQl7qVtObm6alhnijTIPlYd2MjzEu8QV//E1gz8wN0taWGNsmu1Y/GurpVWW
ycolsUiiaaKu9opTx/nomULJUOWj6Zqdxmbwo7KM/qmw3+zd5HsLSMGDRDmIp30AVHvMWFkMVP0p
AwyyytaIzUmnhJkhsn94rEQipYE8weOwYCbRCddx6d6KDT+FZVHIKhpUjbILMVFgQ5zf+zdEo71/
wlPY9i4/UKhkrK96CWHAGl/KurOdklsJu4rKzYLkYfNXvPqH+//l2fnp42M7ebJjjhdqib6mdp/s
1WjAAlH7D4jHM75IheLPNnh71qq8TtlilUoR5wUP2EHgFYQBDqgMxs5LXkfQdVf5CEBj9bQb9Rve
SLR0V1QdVg7KlpWfV50aNKI06PDjn6ivoHC9bAbpucLqn/BXhfxxDJUy9MqaAUdbwSeBFfdSuLrG
bl+uD/JmAnYDG+2P7iBri7AebjBsaAbghAEcELpiWxQBuM9/ScTrO5oHAMKFuI+HWUBheGhtVM92
2odQzY5BkbCxJcGeAdXeVwm3G2ZJijVkdI3Ba+MvjUnDBXMFHZ/ymyGHUihzu90VWq4lGlFr9+JZ
SgizlHhFEKFMdG/GdWgjp9WsnzXulIgJMWMfo46mzJ0x9B3n59SzsdOUWKfQG3oqOgMJpWa/Ug9f
MOMQMY6oFocG5ZDzcikzrnIy7RkeeQWXLYVhaamAsHcX72JK8FADp7rkE07ON8JILiWOHntDdWGm
CSG5nAy8wb4e1iB7AmAv3fDuU9mUBeoIz5Y8/07+F9K0tPRvgC8TnV/GhOHNu4uJ4P81HvnvCzIA
M1hzH4OLWGx5KyCFQCfhaAGUdCej+/bSIGYD9Xoh2zERfk/UNNpH3lQRbtWWblDpAEfmCNGTxc6b
SdM6+edqdY4H2LHjRTdbrrhJoNQmAF3B6LmdF6PDwD27OxahGk5Km7MqZhiJn5J9QBWgZj+hnZWG
9DryoFHn88zfGMOr8rJlKwMjpjapLmuE75EgyoHKr9aA+AFfBegMsaU4HhTbD7fx7WMT/ysLqPE1
KuLokXIuqFzsX0YMzOJ0aiJ+8TS7iOCWn871cZmL+NXKwnlnq+H0mkibetKW1kjL7W4KDdXkQhRp
7UV4+z31U06d6E8NRZOR8i3LGLWP+p6joZ4Mo5bsKx2E6YOImbq+xYzdt480tGgumBXlWr0IYMGf
wreDb/PajQY86+MlK+wtRtpXPYcmKCyLvEei8KeYfa0WYrxxHL//pn0lvz8lUOJ6GM6iL7EbDc4z
MHANk7NUPS3IVoDUP/uLnWsjn0xJf3tCjh06js+3XTzkpnDGga7msbSV2gjZY2YK8pcvidtk5mlu
5UM6KL3dXJmHLQKZXkvE34st+A4ABtx3S8KCXuy8vAhP/L535ZgA3xjyyMQOE6+lG3yEFSAIGNQr
/hZJ1FE3wG/np602iyc+VuVwP/UaMUSdJjRrOuggVdgovPG0jJnOD7C18MU6UcswS4xw5Dk/n/5c
NlUpZ8oDJmXtjIbO9rnj0mbT7clPDRYSymHLA+Up0DbmJ8agPzSrXFgPQTzIGeUYWus2gPgpIp50
0hq/BC7Vp1b3TwJ8DaQyWZOU1MPCfuBghevo7QqoPbn5UTmsj+4MOEWvr3hLElrtPvVWCtKMIXz5
f2vLN12/KlxK0foHhM9mAQ5JyqKU1G+20ccY4gST6lTa6i5kRccO18LJNRpDh4SbLZYejbo28D1n
pDHA9kJC9XMLzu6e2OvDgbLe1EjIGWjlqhySQlm1Ji+n+UnkBR9KFYum+wokkeioQlfiHhCNFC1w
OiCZzzutghYbKdKOfEdWKi7vM3XUHq39kfG3O4acTSeVxKXMwg2JY+Opld+YoxUEO41Rtq5Lx689
PauRoS7hJrrQ9eZENgiU7/m3NxCnzQhuc2EzxN9/rgOV6T50ZjC1K10BdiNV86fC4xBihpTxo4co
mnUQU/Un5ujeNq9YV15ASkKyl1sNkLBKARNabvk8fftTrEKxuTi+hRbVjjuGzLLjjct5+xRyb+hD
RP1P1O02Xhy6W6K0Ls5OSbF8U7hzs7Uh9DHdc4iHkJT5cfhHKAHtmf5c3nBFl4obEe2d8uUEork4
/r1SRFfovLhAvlrlZH8A+WnYenuD7iUsV8xroPNeqh2oBW6EJ6R0KWQdpW1jO87qnZecZku1Npvd
8Z7JKSTyy/9Gz0l5b8zQvZidUDycm1kvRufzhGkZNdsVQCQmKEUicAKvwjYKu471fuPWK4k1MKaX
Dn2VuGWxx6Ulpj7UFlslWqdu+4BGAPGTWiv4DbjvXs+zAk3OrDR23IU65FESdNtJ5uDjUXAWeCDW
Gc43U8+KdMLde0x3sovfVz8100Yhzr7E47+uKhn7WnhOURTiMili9LyQNYiPCQWiYOQ8oejoAbIS
nYA4euozkPg4dTWV42d2ZYAIh2Rs0wjUr5jc5KuCxLrlo9lGUKJHDazefuu45x9X9JHZURQ72Hoi
cVdAx4QaQja0muk72fMDoYwm+T5JkF0gGMcfkFnn8/x2alaU30ylpVH7g3DqkEjgubf6mumM0cX9
jsbFFd6M5si5v64jfQNFy4eyfvQ08biTieUSfIizcnEHZn/x5pJRyi65ydJOn37hHXBYwTOYaHQI
wzcUnb6wYIIMRcC6AMeX0O34wWE2yRZXMtYqsmG1QUaci1MiSrX39SJpICW50EyykkEBSIIqgDpM
69JlC1cCN221XIMtrENsfwKV+k3dInu/YhY+6nSVHZlzpVEPIitYv8D1pL6u3Z8XLg+CCZUOyDFY
NzXVL/FshuhQZVw1P5ic+I+m9Y1DHJKx6Ws7t4hCxIDU155lCisHbPrMYsR7LdckO6LL4fiTyX6l
rNyX8pMT2she+wBrPKqIb4ml1zKTxqOckLJct/5i2SSwdAfeLwzzvvUct3qL0qAs+o5dFj048J3P
kmqOpdn3ynOikT1M0L9/9vkkSQ7980oNTuyK0Rn170+m39btzMOuVUQDkF0AA70UWFOxhzj0KDUm
AlxDFRsulhFg8C57efLhjlQNIHyM0QkYnRocY5mYrgcDZ1Rly64+9scBUsXhkArtaxe2ArPRyo8F
mF0xdyqks5SkQEc+lL2rEFOjNeeyKakcoFR0QwhVCd0yBguZ/Cld0yFJ1K/Ohad6Sq79Q266mHKB
bYafdAm4jyEMqSRKi6mjoLQO6dZOsvFl7KTnMPkVAlxHU9sAESgN3tE97nr3LUym/UYtUBtfvz2P
aMBepzSadYMHKPetZXs5DVh36sOiz6xr5rh1++SKv6VJP2YRutOxA9AJfDw+twdrv2mPR/TVpsEC
FZ22+PhqUIwsbroCFcu3JNK6we1s90FU8ReyK5YMsiBXosQPY5O783DZqAtAq7GnBwiQGt51EON9
OlT7fbSUfPK81NHbH4oriwjxLHD4vcS0vVlPFi9Re3YUIBnKeSFYnAJ1dg/r+EgIn/KCckw14eBC
Q+LUVD3rGi6HScwrW5VpcQh5ceiAx8fmBo1fUmFo5CqBJAl7Liv9NoqToQJqeha5oMCS/6z1QCeX
uRWrO5CyQQjWmufEATVWhMKVtn4KDW0iPg1/Wy1il295pYP5lDHi1F5bUtp/tPHb1V6uTSU+PP0h
HRHyqM5EC+mAOdVh0ckiRF2lBVwympuGhcgTJgcIW5wOmOqXUnojqf40Lv6w9OR2xP+pw39Kl0lE
pziNR1TGuHgnarYSEL8JUONgzC2H1WDFh3YIcFqEixo+9JXhKp9wnwWIz7fklBONqtzWCuhpapU1
J4BRTlvgXFtQ6cg73MfxyPbw6sC57RSEl9MksaZRfzpbwRCo7byEoP5hIopFLUKanFdZU6Q0787j
+5f4h01+z7902bjpyrKZyPPZkE34gB4aFLkrTgkWDaLmJVWHUALUVFj73t6Nkfogj6S/4wRqMans
PgSbANkARkQDg2g+yJTzSl7EdyHkcs5j8FHkX0RFhHnf1RGdojOzA6mjEn6zV5spwDzmCDHmzSk6
WRFRnhIaxZktUmkGxi1y2AbKogxlucEc3dP66DVcoXWLfN1QxoJUGQQ2ib6K1nZZr0Y6xrGlP9fk
+gEYIiI1jv3E1ZZcgqhjLomqZc6U9zMux9epbgSnz1uTHXTHZFHabtCiHiytHBAJQV2FPS4nqj92
2Htat+jjipD58rBaJPR/l+XvKQRDowOmPzVzU1SVxB/PxPajr8PdcLJHiVKVjTSdtgGvi3u6tyGH
6lDnNKWz9DnS9NqZpVL2/YEyHu/rGQCRigExmKJ4B07cbcL7JTyVS7TflJcJiJ84F3+Dp/7yvMxf
09h3OkSuGpqMDkobpCXrF/pKZK5p5F/x7tJPmqGAnfs0yaTiun+ONA9LxA6LHmsIKCEhGRcRS4nP
NZb9R+FTFC07KSXaHun4/aDL3JvJmhlZ6nAWYw6qckuNEM1AzNSzF2Cok24oIgAvzMMpBZGneyH0
t1Cfjb6XB6J2C8mjkCzEP0gQQfRZthTY4hNORUQ2Al6sffGS/sD9SxIdBTB13ZlHJrXHT56zNErq
QKI00IjqJzAkEj/Ubb9jPOPa948KzEu5/frKiiKcgPVwjaPGJDeMhAt9w1kEyrViiMjXQpZ/a2+a
/J61ZJM8QRwWWR3IuU1OHrIIyFB4FSMHmp6XLDr7Ztt9TJA8nFsDrbDBbEYgmggdRtjfdyJf/k3R
CQMZMH2lImOuOO8bQZH7dH5uSOyugUHo1bzhG2equzWHlxWjJnf+3nhpqbyv0TpXrTgstUrNkUMh
TSdW33MeEeJBdWTOMcmUmB0Rr+snUM0LeK0t4AVzPm1TumaxVQ5QK1zyvI59kSIl8wOb23aT2WJf
M5KFzGcTkXtnF3ipPRMKWbIzzFvoWaqL7287siEJjrYW/MDgh9VFQkjXkjlp7pC6XPWFhCwnpyBg
tkIGJl5PmWssDprYkgq7WIS5D4Ez38N/DXi8z2xvZo0r1QTLYCiiBxQIHPD2bgxLSxro9Fr8QTTz
//ujO47Eu46jM11w923vzmODhnn5mkdXSAiL+ZxJOJ1nv/AOyF5+JbvvQpkHXD6u6xBt4IgcYg7Z
OK9HB70oI7boFMDdBktpvJePXswyJ14U9T9gRfD4+lSMZIbg9c2OkJwuT8eTvEzRQXAaZx96ROD2
HCaAsf5QZTYl2T1iSOJOszbDnCCe9q9A1H3McFMInOCXdtrOw1X/4geYcRSJEWoxXxtVLCwRMgR8
kqevBNGcFQR+/KHEIYZlA6qw38cTt52T3ZUoxAOiSl/QrtUvKELe0Oym3kSw0kPs30G8NAG6RgpI
nG32ic7PzZZeICz4wYu8zoCTuUzUCR7+J7iU+AiWNLv3p06RRD6CoTgIqWNMaHQ4E9EBRAsTE1AW
vvDN/3T7VdYqo6+0wMtMNmi0/bcAltZBt+yI2k+/1NTNj5iLkpyu7c9Z5zAQIMAhgXdhNCxV1ShO
rmblsovGv1Esx2xqfZXrqOBJeDUwdWvin2nWuMTsAbE0RZY0fq/U0VTKiEj26+IT3PdX+GiGQoJR
bKBtKkNyJiIkZTjhUVo9gbWb06voOHN2jSpo2KVDMwBAEBRcmx10j59U9NjxjHKCMQhvfsMETZqE
2fXTcUfGBd/FCGMzas2uK3FxU+aD6ErcE+4aa6aoyjyC/urC85qE+RQhtm5klFSWton2xHm/EG14
dwJaTa6OkgIY9NXVaGbKNKnJvA4jvTHBM3VFGWNlFsCrEpz0nRcPWTm+nZIMgAmSDirySgnFzGEB
u9R4qbJDxyvKaC93tqrEb77eCHfUZUHy3AhhzkN54BJiZCWK9MFCiD4SQ9PuIrKNAL9P7vFDzh5J
kxVjftuoa3egJula1fjGFYawvj83kut4JEVyxm7tqZ/FoVKDWVgUV42j4/Lf8AR94xq0cxZGBSVP
4QEKRE2BUSH1BUSQd7ov1cvorePM57UQ8bX65thDEkvtXY0L2R9z2DUc8zZzS4NbeQdsVSKWQ5l4
Ke9qy7jaiUVO4JbZ8t+wTKgVhvGDg9WoutDk5PiKpW6NwQtLJoTOzKpFaTjDD48vCM5t7nXuYC1Z
uU6tEuyQMtA2xbB3tvH8Q0NsZmF9XNkCJjQRKHuDlEh+cADArbDpIrjwyVFo2n+yD3oI+Yyx29CC
WIDKhz7zT2fFJcoMepDixdgoBQUZ3K5HrAcRfjS8ll3yoqTQnKNN1OUbOtgFib8uHuXk78UDggpq
00lzKCYvMGhB6ZJjmfzW3c58X4XXIbpMy9/9ncdlrNt75GBQ8t4TOtI/9gGKUC6/u3CCSTKKAWGQ
NUjMexJcbLRXiAx2FnyvXzfr06TOeEX0JrkPEnvGHIIIw/flv7J74V91+VmikutmWT+nkXn3FJQC
D0W9fSkTYTttJ3zukciaJczQPaISf9fiwu4PA6efS9lO1yMb4zvF6SeDZnySJGDUz4rEtvj/Az1w
4aqM8PKKCbum91rHkWGBQ2ybyVjp3PUx8QKYOk9RFrVGeCU9JzdV4hNnKElU0uBAwwXhj7Qz5tSW
q8H/n9wNJY55q9DBbFsHI9kbfK0Ju2SlP3y9RvSjqnWK4Ph1eLi0qqEnQCU6qqgToQYqPihzEVfe
hM0gjZbbWqAdAFnlrlaDwWnZcF4oaVwsjAUbEc86ProtD4/0RaWaNZFPopwrhzHhF+/1HVoZ6yWy
lxyLx0Ftwk0XUSpufaAg2GgBV7+ozAZt5dnqJh450lAShK2eMOuizCh7C4jBrNZHpVKmnwAsHdy8
wQPeK/KATO87hrXuFqnq8HWMJ2r6qrz4x0q6UOhZgm1nJ+GrvmtxSGF+UZUE4zUGmf1mNEruITkx
PTA9vlBY/e4899iOSiXWpdfAjTIOaUd31YvcfmPe/KARwc0jVIBBAadfA9IIEm9qO9b2yGwlZnx9
hCDAesEg68rUQxmHkt3hVh3WvVbChpcrjdP4uWiXu8nf0KeiQt49mtyiIKMjMbUHMZkn5XWqkMW1
7CSVHYBs7TQYm2KgXKMUpZeLebqgEII1eIz34w0FvhZyK/+1OTiURFAGv+ub5Zp+oSuYvpbgs8LN
pYbjM74XyJhgb9AyaiIhFeiF3q5ngCtBu4B7Xx8bN8s/ZtbEpBDybuvdt5WTtHzNf3ZEL9YNOuzW
DLJ8nGSmz4DQjv5aoVTt+USN/LzfbtXz4aj/Z0iUL8jBdRf1rZpSEJDEE/lCiz60qdGsj66NCF0T
PXtikVdaXNb+CX4WJIAk5SxWtuxi5S7UWkiO9HJDayKEKflpLvVDPjztE9k6jSMrg2vpriUWY08k
u0IglYfpB1r/cMWmynQpJvnOdf7VeqLH5TUsCznZ1Ilg5HICaZKjhtyuTTsorrvowoM3GV+4IaqZ
+PNhzAxFauj7tCXuAnsgkVkSQgU+Q4eTuWOVJT+1/ILRvLYqlTMa1M0ng3TSUu+EGHQsDvHItbXP
KexYE3Vcldhz35JflrLdqpoInaWa1cmxC9qB4C0mq0Ee3idRTO7IeJlWajJvGwkUO43BHyqCfLSN
DoKRGZJWsb2zs/3IhvqeKcIFG+OV4Px34XzPb3PMoSypVj/Kvt4gy4Mel+UKXglRnUQ8BjRnHQ6n
QIhHYc75MxJHKtm22Af0R1ytDVyVvsVDbL2lB2rhNPZIhhBU5L86T+7Vu6uCQfLgSj2Cc5Rl6ZV4
wgbFsis44Jd8YiNDlvwyh7QhduXIaLMqkmPVVCU5Mq3rwhzwDPCU6kW/La1r7Qgo2HPmObb6VkpY
u4GeC4gl3jZoQ2ZTdpw7Tmzn7Np7F5QG16KY83OPTDnebuUxRWyTKbUQ57bjzsw5zMZdE5axEjiA
Cfp5w2m1l1pcW7PdUwUMtaV99Y1Qdrdu2+nQT901O7nBBzOlbfD9qthxKGQrOKntHmw2dKB7//Tv
FR3ltVZLzhc3zD7rK66ZbCNjhQfyDgCrBM8KNPl0U1Het3TAslF6y6maTWtlrFCqKhXIOD57aoxA
INBTP3I2EBeJNLGzE3QEl8ZBCzolzp2Xig5JyN4RKKXKIYGlD32I4Gi/CWEbyLbmeKKnq9mKH7TJ
UvgMo5/JvvPxgJ+wLbSWZA1k9smrUHnyhAe6Dacl+4PUWz1q3qpktW6BEFlUoqfBsbCMVA4tmHyz
vmDhrBR4ZDHrmtQ+FfA0BjuTEKs9NOXMbkjWNuQeXq/xqDNHxnIGjeS3NS5/5NW8E1MbKrM+qq+B
3jg8sHD6KkEU0TW+QoCC9AOvviJ0Pcl888DqQ196WMQSbSfYR/dcU+QM941c4+wE67VzA58aTOrl
DvuDUBAaXezxFL5CcVufZ7DJbaNbm1FEFfgL+lvuGHdRovFXDXIjLeYvHc/Q/HNq8UsO9zV3WVzV
FeNgT/U7ss6TQSgA0+cTsGECFbYoOOMS9l/GpUd251kYeRbkpnzF4AADB8qmlyJnZWusDSOcZ4Bo
yMj+ZUZPEg033eSXJdq+EVMLFfCawmRtx4Qh2nNRT+UNlOYCNrrIwPERXXomYxFHDfGtGlqJzTyD
wMEkh7JlkYz435dW08w20rtSPF1YSPaUJkAuE4TepcHJCVbupZo9pY61K5v/vfVORTB4tFX2wIAL
lY1Cu0jqyJOPjy29n3irotWb6DMF0hGikukmRqUx4ofWXSmU34jYYyuchr46ws0J0+T60pAyk3Fy
QlP0OP2GrWxN2tBX8aLflNuC7+n9HqB2qSEAjFCsMGLKxwyD1chS25vKghxb4TazW5llvaoKENmw
/qT36cRQGAitgey+JKvd47LIa7ULx88W5MweWLjnjlPATDbIhffwFug65B7JgxshwDiHJ70NtHO0
ZBcyIHIK9nt8wHnMiDf76Qn8DaoX548gxJXkrQT+r93nM97aRcTxPkJGvWLaaTokmt5CvjLkt7Ip
va/cDV0JiUcyNZ4JsmaTdcAA/gPsuLAsRjN+ia6ytxkKYYf3Q328/d/Ot1aFjwFFu2A0dQb7XTrP
I2KboYLJE3XJvLcNvirLdFaFsDTSx+ZSAEPMbTmkkkBqBBXsm3ZiKG9zJpJPB8IG561SYxQLXPQC
Y4rBnzo1GJhH/MUyRV6JZToc+4OTjAi2ZWaeIaX4E/3Ol4vxCqpfLz3mE+hjZ8vXdy3y3CHWxEBD
Al+Y3FqTkupcpr1oYlS4yxhao+H29ATYU1H2b2+tree6/fNhe5RAuuIVKENDEM0oY2Fxiu6rF6D9
vCgWtaWaKSh60XC7vdnkzkV8xDutsBzcL4pT5G844ulg1TIu158upEBaX7/p2vsqOBi+OL21RO1Z
FkIOw+cVBovQUzjaLQuXJhawl92IRgpzc9rQuJPp9mfbGMOZ1/v24wbRGu76O8p9O3yFTg2A6NQf
/W5znfKn/a7B0sClh/stqmhoSgvmZ0WMydDT5lSLqUwnBh3f9VroYAPre43TP2wdMgeP+SBF+plQ
Qr+CgQK7GQyho/HYBEUxVpXxYw6wf/xjWSYEtGaU8zvyIfRj5ZujxgqBuhvolNpl3e0buglkYLav
w2VC9AeIh/lqMn+XKwfBaA/Sg2sZpF+u1IG3SQ7XRnTTHH7Mm+70YxqfdYT0T0+EJJrkdG5OmAum
ZRGYB7dE4LTAnzHwsklmyY3LpXq13yTFP18s/SgPlmWvRKqMyY1ldifdYwOz7s25R+cy2bzLO3R1
yY7QBVJOXOgl/gEUFCgtJs4KNDS2M2nEJSLnrGm8o8XntuB7DsRm+7uBwR9Xu3nxE+bwv63RzXg6
YQUsMvhLapKc7ddf0nlMNX5Np5Kp/qqiLWgDfEMY+nUhC0TisF0Vj1ezo6tj5yqLrhdVB3AMrFrW
m/QMyVZzOuUuN+1ODKtJ/aPP1ukg2UsvxBMy9SHgo62jYkkMnWftF02RQ4GBuhHe9V8SYXS5u55D
1lkk83ABTi4TQz62PCEfTgOUpLOkOwrGV9adMke7Z0TU4cdT9CderxN5Anp5INVY5JVayAcZMvNY
wmH9zPg03Wrwd88IWZn0q82s8X1aDqBT+Pg5sGOC3OwHOwTrf7AFtw7M/uWnK10nvI6M9Da/zPsD
JrWSfockGpm+imgwpbyf9CbB6Y1kQKiddbOSGeIv4oncGf/461oqLvAXNzuKUd1A9wqkmg021xMk
g+5E0x9Bd31hTHqQM2Aqyn4VjJjbTJDVZd0gNX4YaP41HDmh1lmoYdlU5jdwJiLF+FAwSiOlWpPh
eXwaG/zwHwVMeutw7jchBA8j/49T+KCpicZnf+1ykGjh+urWmQ5OozLPtGTneRHrcwLrCW1X9ZF3
IadKTZNfFiMMTeLuwlRn8LZMVU/yIOaJmeoD/XeqxjMENLGnRwwzeoUlRBuCk+P+EOVKaGomTnep
8dAs1VPyv3pXAJc6auKmoAAM4rjwCqcimBnv5dsva1oFjPncoHM5lf9obGQUErVG9pwWrxk+gCx7
80qsSp/ACpwfjSEvhcR4Fmi+ATB/+1DrCutcUBYrK+hAplQBI6yb4ZoNP3fezic9VuHWb72evL3O
y8LvKkUclzQH9z6ik+2JeHJmFno97IcW3rKxTERgjUkAMHmzTO4kiNL5ivHLg6n+1a+KFCRLRSHB
k4yyaYl+Cpmbkv4+UX20pjPutLWTZnyoLxDhYtIk602HxqCEQe63z8pWDh71LiVtSeDDnk3lDGeH
k5FosZrkntC/kltiHT4YaPN9lNRVfttbyVSMuFcIXOYW0Lbf3CU5NczmfL5wHASrGyFUOU63hqjg
i5ZTYCAC7Ub5zgel0/y/FHP1k9Qv+hcltDgB8Va497QmuasQMU9dCdzsDd03b+CJdhGQYrxSMqW1
dm35/LLzgIlqFAwpE04vfVtE4LLMFcxuuWBWecVYHFqbg4cw395Zu37ir+uhkPi+0l9AjvIQJ8fx
ZZUEvJZWEVEGX9lTWvdJESnfEoV4lTRoJ6mc8SzrtobMamyRjPUhHIbF4cm4xVrup5gWJWs3RCsM
cdHw/GV3svABbC0fbZm9N8lo7q1foGA9wYy00M/OWTtKlpbbC6hyah5fOVyPgfGueUe8b/KnM37P
iGX6edrEv0XSjtGLdnIr8qMW4ZWv9ca4oNwslP4ur1NkI3E1aY1VVBRyAnuy2sI8L3wweSeg/m2l
9fkU4AaaRugl6/L/jdYkKtL6O+8oG2y3Q6a6Htw+9l626EN5cnVfiQjTmWMKWi4fzOmV5Jpz65zA
qlytwAjSM8n2aw5shymFfmXl7a49hKtjwghhrnnsCzYCNsY0nkmjJM4HeBXXtKMs+ETSBuagwiUo
zcVBp5vi1oyNed4q+iPLwRRSovv3BDkXoRx6CocxgVkS1aB5GnFm+jqtClkSCik0m9RIUF7ZBfbb
6HPWMaNW04vhXQqxmEuFlFT/02hLWboEby2tl7yzLHYr6lmrNjgxu4R3Zfw03OXQqA+rsDMu213W
8luwCgsSoW6FBl1Pr/kwHF5/AYOuzCWd5TR6mH3V98LWcHuPKdERxUp7S2qBEXIPj/l8kdesF5X6
hu8Xs7Qqx5cLbYI1PfWB/Gb7M/s8EXElUUTc0nnP/8oEUwbsn7gnaQHtkb/6XjjFh8vhHx68L2xT
DR0eBP81P3IweY+gQrB5NsDHuLgett0QsgV71kXnRvL0teREFeQmo2TKW6yyYPIwsI5zdenL+mBD
kJMx4ChOSqroqs7BIoEHvrWXm0zHJhKC+62B1hkRLCwDP2I4noE+3X/gjeuHXwXZNhfYG0igQK0N
qKBvDVYx4Gedk+T9jBQqgiyMN2DJZdvbqToCknU8eZS58aL8W2nTtpj3yvheOCnNiMXz+gk5sRiq
XahJ+d5sXc93V1lQv6C+O3jYI5RSjQMpDts8hxMGosXJnRPfLsJ80UIuukcIa8zwCoG67UeBamcE
yf76L+JGjpaDz5v8xIw8B4m7QHOdcWGs0CvgthfhvPv9eZ/phrzPgpIGLoKQPUYOA62UgDUFuyec
XUVRuAVAq/wKMsXJQl58jzQgXcxLVjXxmytZ94eNJPRV1oGa2iPzmGftb/VF+MJBhj9OFbZ/tvKF
YyrwRdi9Yfw5ov4Ufvuv2aABoPDAGDDZvYbRWelAN+aHChRtZi9k3jM+yOMnnWQ0pXd+kJ3Fncoz
Ov7kIKMHyEbdo7BNU5CGhgKV3mGoAE9cwTEnJu57SVSa4RQyV+i5jMhAbA/K3RUj0Nz5Z4zr7Uvq
2MYf14hd8+HrjHTtSSWJvayJugjXh4jQqJN/D3GgEDFxEi0aWTfu5YiMJzvCz37eWkJaigM+JbLS
cz6ki6dIFqJ2I9zs4Ys6Y1TcjHJYvs5LYiVPT4RqqBOK0gpYZ6BwQhLgNSFP0r3twsJa6BfS3EUp
ATuzDkUdRiwZghqk00m5zqWjdHa/f3Mr6BPktKPeacErviLzzGHOVFtDscbAR+bW0j0wDUPGAF0R
uy9KyTWVoy0MCcVNxKnTiR4kr/zX7q+K/wnhqij1qZjvIuj77q/FXWogDW/ZovNd9XOE5UVPhyuD
5yBqu6MWJ906tLN4uJEs/FxMG2tF3J2t76UCO5RMWZw8L7Wchun+KFn1Pgaj41USDM8zUWkJ3/dT
b0r5K4YcbV6BfIdup0D8tXS35T8WgMdzjaniYsdZ3Vuznw/RZ2msZofBMvzhhqG1kUJCYDgnFRF8
aWzkY5vWDq7Y7yky0GmWIPFNw/LVgoLx3VdxXJfM+CQ1CzvYvGDpGHOXnT75xmm+bDoGOSckUPWS
bCf5m42V5GdSCzRlMSSKfkmn04lLr0buE0MfTRAH6DnCKE77cakwz0Q6x6KoZkbjZyBNmO0Ue4XV
QUZtn6p9ifcCXfz06ei49wxtyAnoIrdhWmEjml+Vkdra8w7BEdr8esheomDKTw5Pbnu0MJnYdd85
JkQJ1boIopa0Sj524x9fTeu6rhpEnC6XcshZxO+f002RSq3LEi3DiE2n2UM62OqrpTVO21MDLqVr
mjF91KlO7p+zbPp/nhobRX0DO373kBE+OtiSnN3gcu8Pzxsrly6wukTk9zKzOgMAx3puT89Oqpet
HRHuJzbVWQIrPaEJ46uFK6fec6zLTybn+7EuRihwG/5iZelG9kt97gp7PbaokKsPbK1iqmgDM6co
d5xDIFPgM7y2Am4QPV1UD72hBVkpNTtziS0bmt9hKFTDorQwW3omQrJ0AtyeDmG4sPGXzMXKZViB
BrXP/gM/oDRxDmeW6EmSuFFjD5dXHTcjKQzLOqTpVtnoO+zdsoQkhJMwLZm1Zldr/vAhsnEwo6+c
kHJTWr/Ptuw5GNw0MU4m8GWXMXU84h4Bj2opsIZLBNhb9F8VT3BfxOrOaaLoymy1ihseHRLbpCbG
1ZJvTQlv9Ii0YKnhPuk86gQbf35OJQD/bKrYMtIffSybzodLx4CrBDUK8nMYvgb33ySueDUDy606
Ez3WrDnXsSj3PuLv+2lVjCjhyqyvwLNGVgvLg/JCK+Rt4UPLciak/u4I6EpJT39v/LBJS7o3XDxk
VTv7Y/fzzOTKLe8Yhjw4CHw9rJMDmDsKmaFk2ydJW0SZd2yH/c9icb5pcZCH7BHZq+u8+KomX9Lu
RvR2mlNK2VpKmOkOjGX52wizob+/qahjxLG/rSY/OLNdZKecgWcS8l6v5iMLVNvdehHKIez0sEm2
+OH2i/Bhk8GVOX9NcA+/T799mgJ0lD9tB4GL9rHKx5r66DswbYNki0J6wh0eQB0P2l1ralrEbdfS
lDkqUHx0akd2z3Knz+XXs9Np8ZsW/ZBn2GCSQ33MZULxLtAUX8R4NQE4WtoCyGKwmVFQHVidP705
XvJtP1yDQ7OebMM2X/K3xwwz1xVrky/dJmyzAOSxWV4HPRgrQ6CI/WDoExTndQHt9qaRpHxfTVuB
9sVALMHzP8ANJqPah7wA+a55axYoXRdrgchIQcjz5vb6pNNcRKZP3XlNw/vTvSBjLWarz0Je9Djh
37TqiRj5D50jwV0SqVBs1jDUW+3Wjd4qpgDA8xrr/SQLXtsW96gkzVbDKgv8gZlm9LJQHZRIKpgo
23PPTs27OL2xQwHdxWC4JKNzDc/m/upNvB0deeXqko+YUkIzWw0ttFZ//738GUNgYp5evcp35Xfr
FX/P2jXl7K/7mVULpqMzZVRO/cyBAm68uN7qLitgBERpHI428PUKr8dQ0zibpN3CjmtuyuhPQ9T0
HGyUh9QgrNEOKhe8Y3DnzjYOH7RCXmhSPcUOWSUR/d22SnvHD7xzIDoO1KmNxcLm1LNaO8JTkZCQ
76lyap3bS5L6PTpA3tl9/bc64jVoEK8JHxA2RloWTmMQ5nKb6PoNIv875nGBgvMrJVH7RSBHcb3u
1wK1+dUtm7HHmQPXHjhOyiL3T5LbOljU3QTtgKEOJynJAAgkV9k9+BE9oHDRK+m0D9xQ/rUfFmIM
42ZA0ZbH8CPPN5krR2WobbC8U5jqrjbdGKBj1n0uDHOMRa2LtPU1sBXMlzMrTEULLtTUrnEWqwzZ
d9kPKscFV01Ic5CeClu374jqosjUuZR4lTbkYTQVmvzCAiLmKk9FaOcYyFj9ckPVnkJoMA0V6QDq
rejr9ILjfygYIu1xz1SnLi5ELNA4SuXJ3aTKLsXTwP0WhZsop7Zt5QuqLzgHYygpiRfrrykWiSM4
5VPRKb9LNjZsJ3+lukGFjxdsYnhl6Zny9bnn1QIrziqNu8IbL25pZFwNL3MW9v5iH6T6ujtVAPbj
Moh7Bw9Zcs+J8AquHmncz5mg3HWDpc9paLN6RZMK2GHCqEFPNcbmVMvy1LeRFTbQ6M2Vz1myc3zv
5VRfW+IpoAbVjiuJAidE4fbkXWDGnsudhMyzNmkxUEM46Z15YXGnVZQ3mCsy6G2W4iexDwHgHsV1
Gt57hDwDKGSRKZSO/SitDHH5Bg4+kaPvVVILLe9a/W7QB8xDiyIy9uLsV8NzF7XKgJFeAg7UBsnF
J7pgdOccEubp5H0aY2O2Dg9oE6Tf2S17gY6dtyRfrrBE0HHWgRGaCu3+Wa/aaryyzYGnshsgcLYp
K19MrOCoNz16pZTa5eqljx4SJEn8ulk0iOXAK9DbXR8rN1PF8K/LWOuFfbgJuRBE/ekBw8VoZgQB
8toL1dYrnZqtv5zLC4yadttEqgHn95DYHJQ/pfdQsg5J9oTBojLtXTfX5pJf6d86GmUeLN/JvsaT
Lt06APt+B3wvE+rKl9EzrYnZNEPR6Vx7uxPnbh11Y82TV7YXRvY9KbZEUiICdiu1C4lJvGTifyfH
MsaKQMF84pN+Nr6QjIqI7tllihXStcdGUYV/wDSZafDs9YZLHESNKJLwFYaBTXrv5a1tMvKs+396
vdQrq/vR9rw72UoNs3zEp+Uuema1DJE+FZ1G/GwGuCliOt/bJcm+0fuwUc5o28X+GZ2nqZy9HN7y
Hm+PaFoaJiVbxMKuMNSt4WoMNb4rICkk4MNt3wazD9kDm3S/yiqeBk5GaDj3vP8TrTXjaRNGFD1D
wBxhbrswYkqpOvCh9T6F83cdR/yCDh/imCi6v63LZtkudC7GqSFaMcB3qseG3UUOpnUYiaeoKln+
8AjmyQFlkCRto6/H+tG3BY8V34bnb2m38X2ZrwB1IJGR1VVi/3VTA4BwdGeiH2V9VdxVwNr9fVNF
1ZXDLG/TX+KaCd+4UJ3SprAQy0yHkjdT8cimDoRNxJD13auWNaEM3FpwOgOfISq6pVLXSLAgQr9+
rC2wX7uKiQahpSU8qWHTbQ+zcdN3UZRyc7dzM/PgAzoNm+DdOR9j2AzMnoy8Vt3fYAmrUgdfAJhR
ziW2Ef65nG9OGNoAhG9VW2OTXNxaaRKdlG4iWdx0VKx7jryFCwoLJSGR1sgxLTMZMK8V/AQniJo0
MfaMMD1RsKXLphMRABuoo6ooqXU5/EvFjz1hG04pNQ5yxlPteP4bpDcZsfv0KUt6n9KJInzYpX9r
W7bycaKayopbwss+SqD8gGRY7YaVsZQwSoHGP+8tTYYqNLrbZUIM1+3doC8O+PNscCBtmsRzS0Ph
1gnu53UWNiyqrlKeHaq+o1O8FwebykIjZnlxeeEAYqGnbMe43ckWcipISnCl5faOwYTYV7MFzmUn
KvVXjUzBqbSvPATgpdKxdt7hIX6i5g/733cV4svnXOiZqnAovrYjTInJ5Hv3e+zBUDIt/W186Fdc
YBECpmKXZmkWS8Fv9Gf2NHRjaWRYeOkbjVrrDuged9Ln86d2SWHlIhMD1WgxfVglHlX5WsRt5tf8
uwuytOSkDDKebmH5jeTBikQnv3rbYbYXOElW6BhG2cgYssGn40kZ2vPxPYMsxRIyOUKmDLi4u518
0FX5ugZ4H3vo7cfoRj357JEoH1lFQJkQfm/DVfuBjehMpu59jFVO9L6dSp3KE87cGWpGeQYffmH/
kreN7yzepzJMa6bgAon8p4R0WzEPZxZno2YHxe0EfnGPmpEqETrXiTSeDbSXzkqx1Qjq+NOq14Y0
NCOp4AjdqMrRoO+JMdtpa/ax7+GznWJ4MwU+tMs5mI8mIsKzybHJZVWYFlytoPn/qgcB+h+XIJm/
TJzbAhwJT+TQAEtZQnfN0/rJ7NH/G0Gt4W5ftJyFoZrGb3YrbIkVBp8enUbuKz6OLflW3BfgMyhR
YOmLv+S/AbMo5BN6Nenxgyw33MiAAN1QYF2zvgRt109GHWJNj12nYB8TMI+8vVJiX+bw2UqtAM5J
2N8TRAfNgo4Za99cy6FvF0EGWiLQYy/Rz5TyCD1Kk+4dnIBnNH0GG0kUcgIy5+r0n451qBWAa64b
WZk3PdQUM28tYfcKhCt1TUS38K/UeyYelUNiQAXCy9aE3nFItZg8TcmIr2GRniYjDgOYCZhyHTZa
pyRQmvI/1rKBswDdXT+TckaV4hDRFK0xqgHEHPxBDwFLBb7Yiu0NnAQMnXgEzIO9oxUkIEAlG9cY
cxGsluFhglsTQygynVCFEOn8KV9Z1VKysl3sibRcT2WF/MEx0DC9PxEzYhtqxx+vuwgPphROniYI
5W32pIzgUMVVS3Gxe2iT03V1vzI2+WyatOV+ZqAXu3S+7MByCEdJqsJ8QKfPKwE6cTm8+ZbdYfd+
MP8n2A9U+fsNZ6XzbJ9vcBS84kp2acKqa+U9o5zWmbUwobUNCHtx7isbOPoJtXXDxfjo6xpzvPCQ
1Mb+G+jD6bywxg6/SVlAty46yCUAtz5McYknOohbKfwzDZZhG1uyBNWs0okTF2l4W1u+ED0j8vxe
MXAEXaCsk5PFFOpaGNT8NXDzHhSWmrsUuBl1PYttrOl/lSKnfZcSkMiFPGq5QlaE70tcinxmnDlO
nuSoOw9w2DfhQKoSU3kGBxVYVZjI6bHFHM7P+do/yhX/9hwUMqpLXXRFqxQeudvF71N/H0XykZ/l
if7R1h5kSmSWiDkofAtp6biO0cyNMMlA+fNEUQzaS4ubeFvF3OjzXEAfDTn6KzYBxd4e71mHLoMM
wD53KAOAXwMNRJkvDI4JgAjo7wQ3l3ibb+fyhbAw+ldx1xrg0CjjQ3Nj1K0KEbSc0ztJnljy01su
92bir+/GhcNPcYNTdE/LEgUurXfh7vaXBD6TXemeXD8zCL7RdevQEEHXlkOULVU+0q5pz39QRYN7
z5gkpkMz7gTu2rxbDTNHDotQtG6Dd0yulr3GLUfFjTXW0lIihISSC/FxdRQQ3jtQetYlOY5k/joo
7+W0JgvqWVnBQKit2G/B79KKWA55UOzoY+kzKSypd+nJJOyECoM0Ns8iQ0uPHAnZVvMkmvbVt29n
AUV1UKAU0b3n+ek4R4H5KQ8PrRlIbHRSnvgYYCMw0RcIerLDeNypHnURIPFu8DNwjth8JsXFVzVn
oCc1+VpYW2RgEkI4bPyW4aY7EEU4tTOHx2d+9hIMLfIGJ9SmwT5TCzUPCrKfjkj3j9GK++wtnD8i
sg1C6hs95gC+/sp+3818d2enCvRzpMFPUW1nx3XxSk8KVOltPvmJ/7HrPDt5c1AqoPfjHSc2gjep
A6wmgBrqWRVQnZ2GO3rLOB82+4cwZOsutm4O0C2Dpx8lOwgtDOoewr2HpauMoQZ01LR+2kRTYaPl
ezJQTM7V/VV+hP2RCYtqqULo0pO8MEeMpqZTGzztDay6nFNkV1ObkA5qAcbfypV5J9kQPv/BdNdX
j8IvsnKaVp4bhr3unkhz2PsuPSx4OSVZ08tiJkb58GU9vedhBox++XaHzPQKOW+z1Efx3R8yL3b5
q6rM7ak2O9v/7R3kslJo4/aljaCHRCmcmqgecnpvCdCcL0t3nINTO9K/6hoTKu77XOWh9I2DMhBe
zxFzUHT0gqe2e3iKvnVAbZEcgPIBPGwaTIKte///M+hTQ1c9GEwfQo1TWxRIHmRBhN2Hq11RqYtr
Ja8flg3Pqebwx/IUN6Nd2xP5nLmZ7Gl1jOQxGqGbfD8KrYQ+ep3NB776p+fWJO+qGMAmeOmuZyRx
T4XWTYXQ7dEjCiAQthQysYuxYrrRsuEjSMd6qoymIe4a4/CO2ojbDIfsYt8b/TtfIfG15k9Oi4ZY
Z299SgUTM7rSxouKG/gb7RtQuOaduztJ+GXmENaT+M1eNnfi3QhSX71Chi5LNJTPQlmBcx8UUKJC
1p63n/hXYOBV+3jsMWzTTRJeZ1L2zSc7vJZC9lWjTfCL5Kgxg/pDOlmNk416fLLltJJ3ag/fdL+w
Ej9mrCQd619jFNHrLeZ7XNf2tc41E/umeEm73vVOldDqtwpxmiiOoz+diICanzowiMg1BT76G5OM
hh+YVUL1RMZmiZBUELF/CpWQc8NlfKz62EGmDtFmBaz2PP6LSVQc1LxBQuG2fIG/ICAu1GFYYFxs
I3VJPLgmdmlE7OKZ3M3E7Roxj0B86pS2LI1cSnk8dHXDS44ut15JCqP4+OjyJtEXnOU8XJUFxqUt
dOfrkGFnDdGEZjmCQuEBYK3FM+X1HNF98qbFjlctPAxwAcdmIhUYl3YLryzECJ+CaLXyhE96WMBj
+GpRURW9nmM4w5VkSZZoLWT2Y+n5PT5vQZ9fy5GSkir/He+BrfkoBr52yfUJGXWUJgDwJusUAM0p
uH0ApNb8qRZl+7hQI/5VUQ8PIJJwfDrsXs1ZF7ZyZZ9gKhrth0Bap83qwk7C9rWvbLIQA7rrJ1BP
tU+g+ePbpSP8Xrs8GTqUTe9dP3CnPhHV+sTVkx1lfz2d0IMvhh2sDdC+2rF9vA4xImM9+Z1cLjtE
6QF1So7kkGRMbY3R8NFOEqSWQWWtwztSe0tRPqHT5NV6FlKweDgP7wdqrEOkkxVAIAq9nidaRlv5
1+VybuDVZSmI2qrQKmbBLGe5TxfMezrS2FAXXc4j4LE92PKj69VRyfmrXd2XCvhOuQHhUTirmyv4
viQD0WuOjIgw3CptXEZoWnlUJ8gvtqwDtnE0y9GZSky2SX+RUgfh0tXePwdQpMePH7QiF8Gnrgio
SRW+GkavdgddBCxK10xvWU6DQGZabgOjALNAZx7HCa4m1RbH7R3UMA7LhQiPsdPCGjaS8MWYRH4L
hKhBD8Jhf0OjWxt/08jgaEnkMlt67VZZIsHZHjasTrEomqhWSZOTZkvq+aTOuXJREdg2zEwjNWV+
giZcubbnODACZCQQndqDxgMjnRUgi93RKwxhhPNQKMF0hXfWz7dAvQ2DqW7wbttfLYIc0Fp+66gH
uKqBdrlDmLD6c5eA/ldaa5WfHbeq33VAW1KXdq70eYVhmuMc0ULGN7P1jo6/xgesOZUvZTM7I9YV
63cBiMItbQ0fLS33p8Qyh8IOaft0YcqUMvygXguQp4dIgLQy7CMrTTO+SW3gGQDT9DjcSY0JBUEg
Ad3nknu/I/l4AAgU3V7vn1mJqJRP6heA1gvYUZ5DseruirgucMkIu94mGCCaDErKi4fg29ph7sR7
nAXemqz8tPxqo3FZD8201H6Px7z+g5Jxqzt4z+gvzZfUvh5wDNilgWrDbMk+OeOE3xDoV+hkgx4V
Ac2lbgUeMSQygbmQ8uL+wVbiL15AZyrzjwAhR2N2RF+2Xiva7OPnDJlR5ANE2Ou5YJUkA7IN38qU
gp50dlA4d9F0Mcv7oOlYASPczuVOmhVnCcrFOQ5oSsHBNQmm5bTyLu1wW9bfM/dJloST8u4ot0Eq
2n8cv113TL1QxdPqbfdnPUUbUFAQcv2+zMqfxD+SVPLT8jODSRUS1OILAe0Hchx7fhSnFtBMcGYS
x+4ieNKMSwhRd60VRvu0xY30n9cHAy6jYzp6wnoD+uKxuJ8Qrc+JT7vCagyQpLV+p3WPvfRDJ7M9
qZrA2/JiZkR/3hy48i4vCSZhY1GHN28buci3MTNmjcSmomDU99pVXz90HpI/X/EMTUuGv/dAEdpu
NdbUrWlwgD9GHTWkXqdClpxDtfccNU2WISZ1mgw8qqUnkI6I/9Xush03i+qX9yyD7Oe5CtOOfxdU
1fqjUUQ/AtHBLjxbBMo75k+2F8HxrB4mAcb+Sql/BzuOWSyasa3PWHtpqI4b7MjOqzvhZ5DtQXB3
F9aYj/Tu8GHdiFy0ba11FkH8sZBPh5pXThmoel0Nzs0kgQyCUGOzJ2QnEjap8yhX+/PDb027qxGL
KhPrIOVerCPsqPWV1VN1XxVUrctJD0tmpZrXxBBt5/HHnlI8s2gyPghAGvH1C1J8vFelqQmr9yXB
bOBFolPC/pTh9LTOcOs/7uPhria5ffb6uR/Zjmz0ZkdaLZbhj0fErIYZrLCwITi/FJXzs0Z0ffXW
HrN4r7n2biRWp0fsdc0IHho4zwkVX2ji7p2jWQx0+6wql/1z11TxwlMYsCQ8wCi0xssj0tt3abCr
JEWCBAurana6mP/CdMmiUozZNomO9/4YIsgtAF3KnsyNNdH+N1BFDO35TuEkyOZXax+PHNQRc6bf
ATxE3piLD1u+AtNa680ZFNNMEymR2qHjVsNZF4aOdHRAsfVt35xwJbciWbo5N9K/q0wfVx1GqHIe
F9S5LtGCfXZZWbGpOSz5lPr/hmXMBFmICOBNvkMKVhdOHbVP9SJ3yVxCHcJ3h3QnwJgx979Yxe5k
CofBROixUXPlmjrVT/u3lmB7NKklUKDTS4ltYliqYUY+NR8oWaaVgTlHAcogz9n5N8HOzU4MyYii
G9thG0WdzIpvNpWKtviRo57g+o5+6nH5GPQz4nF/Qt6vfd2KwXXQCKsd0OCcYr6pWPORU3NA5L9Y
6v8s2QHHgseabslGfdR8TXPmZG2SaGGu6KTTfG/NUywKhfpKinQGS7uUWy2eckp235kgp4sYlEyk
85oqzgGBT8zgVaGQ4kEBoabuF3ZfiKdEIGLPm+LGfrCvJH6KQkJYRXdIMDzbxbfn2AtQzSuQ7lEg
ptApVIyeORB8zEksztqPRghmiKR5HomtXsRb72JQ756aM7/Y019TEMi/B5jMyIrFpEqJRR2NzvJn
PST0QKfwguKWajaXQ65ZJZAS1d82eAY5yQLOIKyqjB4OqHkwHJ1kCtSYWXmTjfmGIZBsTQfHFOUL
SFEX6cKJCp5mD8TN6BZjJ6rHAgF3e8TShBARPvK6DA0zKCWqkLgFDudsXGOVSanOChALIsAQl8VQ
LoaLJLIgrYviGrKkAioBEa68PU/YtA21qT7/zDgPBQHTvF3oushlavgIvXg9zfb6j2XiTDdY0Zdv
9Rkq9zBI5tgNgL7glYc8uivorilXFEA7HkstHaXljBq927mHfhjnOepBYAukJ1OAjMY5V5Yi/z47
zpkCXrUeYenaVXSm5yAdBG+bnhYb9H0ZohbEIWrA2+r0kiAn+tjNwLPbu56O3SAC1CaFiqu+PFkd
dG0DTYWlcIqe9jgSebjV69ioyFuiSghwp7kguQTfg0/UL41pEqHxOiYskrYxi55Gkctg0b5OkXbH
TOkpqQplEdEuAYu2I/7MahxAZmOy3A1/cHOzRI+mKcH7H+F7+AM7BJYyzP3cOS8A/DLDFtwzZy/P
SPVpKCkwqfiXTIHRShexLUAkXCcNsLLCuSaHT314HvWfwi8BMC/DbovwEcn1wntjqXIpF8lZhIAV
/XDsP/+Ch2SQOSaWEWDjdiisa3LMtt9Z5UycJvTa3GEawY3D6hU/Aju/aY1nRT1gH6FtiPpk9aAH
NATm1PDgt+Q3wfiznqZrezOT5nb/KHoL6yS6XU5XiCCcrkgWkfBs8pKGMSK4WKhXBXWE9/54hTOV
YGSXzAbvcD1XhAmRYcVUj6E5ZxgTC28vUKo8VBuH+2l2prruL3wFSz+0LLb1U9mTQe/EjX0fal3H
ClqaB923i+k8wqiffnnLNkMzEuWvreDvd1wyUy09XB3QFuuMxd6hwcIAZuRa5sRdyPYaeMTF5UE2
OeHd13BeP+pk1N5qQfODU0lA91CugdsgdGwnYdsr4vnemS99GOHRpr6R9RFOdmVL9qGlms1P6Ntv
4hDQFez8J+e9+57bD1mZtGBO2W8e4/3rdIWQjpZOtJor7bqMNCllPG0YckFesP3Ape82D17xIMou
v/Dig3bRIUTjYKNWAPLNcQ8V5dl4/ihke9EXBZxgu7DnfW3wJKAxTpvurPqm+w6qFOrkn8CFS5PN
FsiUce+Cb5Tn0ke+93i2Yl95xx3ND+TNKUeMje9kORO1LC3PjyTzPldboR0OrSsK2jpQLOqupylC
UeTNMHJG9lnTKQZFa8VGjDi854rFUYyFt0YdH+tla7nMNDk9Ghvo8dLOCS/Rr6tlEioqv88299++
tciCF8e7jL9tE9supAJ8b4RPpP0H0Egy6EPj+ThMSJt8/2Uysa4pZohhR/B1KD6iCBWOsieEw2jL
WkAAU4APy0KJX1njiUOBXkAw0am4Rvqp0OkcDO452YZ6eJAoFGUGLyo63mAM5r7TiNCThn0l8LYr
FBidS4LYaWUOgqQOHQ+0zFUlYKsuXN3znnUWtGuY1wFsXhSduYSIVBukU9ZfkKorJhmh/ku+dfk3
34NYmIJtQcJ4E3bejGMeVywV1+LQy6jj2FQO5mEc3tBy4n9BacYkvMIjiI8pQnP3ZRb6GI0WF6Wv
ks1NxnIFMmru4fpqfy0+Lh+BjeUmq5hM7psUVa//iWyOQelO9hsZmv8yurF/KHMcl1qOPIc4gOwV
CO5sre66RsoRt+iniOBPaXcQc8EhGNS0fWwnZ+w4KsR8wOxdOa60ewFy7gRJRP2JqsuEn++zI25l
5bLCIxVr9ReGwJFvYED5yxbV3zGBR3mOacV41tDsb2nPGUUZQjwA4lQIlMktCPuPOagjlpGpvg25
h2SdmgLFRvsg/R1h3RUez+IDNXZ/hH51vcjkBBexccZ6MNfgMD/SUdA1SVjsA+kuoAWC8djn9MTq
6HjZqKI1jbAZrT1TkuuGGLvLwNQ5AwhtOR/nq+CTm0pOz8+mvzingIYqYL2hStmscOYtYFCak6j/
5sZ6cJCHD6Ws2P9aafufLrHwvKuCyP3HSuWVVundrgRGxe/mKyKFnwhpVyFDmVZuz7BUMvNCzlzJ
Vjd/HkGOhG3CMnEy9yVJO3A7qr6oLUq9Xerk9+d8BeeC9UzSkRv1cH7wrA9T1BMkiVFx8ewhltCu
65wnzhymE9l6rXdGCayTT6dfHOQqrdL7x5Ndsp76cXmCKRFiTANismLFX8FXaocD1fPWs2fGfimJ
9IKNpqSN9uUtJ77TvLjfTPTV3tudBRxVXyoliGN/UB5EqgxMT1AQctngBug6k7orEMnSBzanTDQi
sh6mj/f582TRK1gA0s9iaC4yS4vQ/R61Tr/hPXDTDWcnWqEei1bRELIQLuT85bDxDtSNzkQ6D+ap
gkSDgwlqmG3OAjw+/p0S3uADQIdXbkOgiUZr9gH248nXaxdk/lG++PwxwLt4DPABoH30OinEtz/O
w7ygNQ9GP7uueqL0li085RJvoohTfW0JaqMBrT4qkyOyWA+qt7JrA/RvQf0jfQcBONwEZJLGvfjO
p3oi1s5x31byLIQ5tgFFLteZcx7Vm1XBDBQAgkZaC6KXRkwwBrS1wZiC72pc40GI3U2XCU7BY1xn
lCJSe0J7X10Og0TI64/jPxM+AH3PuZBJmxBMviRCh1yh3ifwoJqYCZnAfej18X2mz4ZAUWVNA1SN
P1eUnFgTBCqKCnwdNpqFfNnVIWUKPy25HQCvs7a1bXckbIHWn7PPjvSvz6roE5uZ1HEDOZtWjhGs
Rpml3iPH9HLjj+HVK6sY/EYvrArdhmrLKPPBt4vv7DGFCoKXjeYTrll9PVkCvPGByp08CY0Juu4C
Plp+NplBSY1IhBAVxz5xLkWrGuEH20isYmAprEOLs4h4l4DBlvzinwF/zGBJ2iQa/Al621uGlTCv
uwMekfoYQQQOHV65QTpOshg2M9lBSjV3u4jHDoFu7CxrHFR7FGqw3UuCc1kmvYfVDMxOkGbnYRdz
Q1+5dxLNM1S2LGw70dFC60z9p0dat/GMVQG/qIqZNsfQM6DzLD+Fkcu9NUbOFUcosxivTXvH5x+1
v9/VJvXGOJ3ADG6tNuaYOFRIGUTmLdt3o++x6/0PMv5sxmCcsa5Fwl/ZsznVudxMKgmnVyBsV3YR
M+VtsNaKI+tiJoDiBT02PtDpeLbPE6Qe9+AiI5izi+2SNE1Vvk+Znt7EHQFX+iWAasjDwY6XescJ
6Gpu15t06bVq6E8y0N5ipuWddXMpmtXG2KCV0BYHQJe9JU2mojA04NCq/ueqaTLlzCZf37nRKI0s
oKQr57kVavm94i1WofjbqofphpiucZuMd5lv/JDaZpyA9BE4rA081ckmotnfaSgPCcNOMtgbfO1n
z0a+SB08f+jWbe1wZer1jWseyBVdcq5oB2ig8vqirp2AuzrnRjhpdOkXBhx+bAmDrIaVBvbTBra8
zlQeWqwgsE/Qqbfz3pMQxlpsNGru2PUTg6lsBBQ7lurWOZLV42aFKet3lrgY/0BH5GWauFnZKRaN
caBLq/e6xyzhbKOLfoqFNFG6JMds4naZ2SqZZ5hTwALITCqZnWeQ4FGlxIpFNWyY6NFkwrWux3ms
vf5BePiC1FCKUp521jf5ga/zpoMd8Ki2W7odS9MZf8BX7orqTK/QZZZAExHRldiWnCJbQjPxIBlP
zMnhhMIlWigpD/EZV9GtnKBfgeynpmJFBrRUtOdrazYLPb1jR+4bKn11dmtPARNilnQ86wHWF2GR
Udl2sdm1QGe4IP+xELyQcCw4bAkNUmjx771TL33p/lsTNP4pAPTVco0WAXOFI74n9uwL24yZdAHN
uCTyBi0KOAuWKE3knF1TaAvbV2Jt5PBQ555hPYMpcdHutJKxvZFzwInUb1qMo6CduAFa0Ald6zEx
gAgcaGZhBV6Tzfd0WZfQUFaKNHzyzgOhhV+WNDj8okjeA2TW25rj6m21dwofblzBshjU/9Dc+qQY
CiMnLVJ5Ck31YTwevIF5/TrKSyXQnCo7/vnU9Fw1SaiyoSNoxbcMPA8m9ziKrtZ7n7N+0LPthfLk
nU1lxoyIqUetnfS/WuC7a/edyqPVDrF1eDHaLOrpkTU2N8ajTx13Ghi0ze5fHGVc9HcVUp4q3ii2
4iONYDRC6ZgaknMVn+HruWtx0X5sJQreIrEFX/2PQa8RFQKDg3FouH1elzpq9PjLgzE40NABbRLw
yuPH0dAbLYveqkHIzzBZSvLDb2+CLOvW6FdekXH2HIl2n7enKLiGhxlgdDsikXAgJnUwSZmm//Fj
ec8uSzGlPPTu7zkwH8x8L0WPkH98Q3FCnSsDy0yrGl01Hgubyie1c4rdd+5DcpfkZd2yNEOuesZe
ayZvUgDg3k3vRBQDZo/DuUuMhtRkzmFPWEuWgbJvmHfuxG5COVshwuADyI/+I7XF3678hHjm/KVb
IHP1IendNAZj4wla+SADn4628cmj5sbQtLKsKP61ZC8V7fuBzqMp0N/SrKN7H2GR7qdIt6bvUEwY
ITNMGcYlL3l5i8xuphpyNzFSYxP8luHR36AwkDNF4WP5hBGa8QFBs485dXWirxzlkZj4NzbSP2XU
Ww8t+BJOTsCwIVBnChcs6y1ZNDMjcTbvgfqynE1S4KMDQ+CVs+0IznVJv6GPbl3hyfIhHWuVbW+k
F51rfo8it3XtF7/MKshDRyzisfCl0Wmgq9cKsa00GZ8zZZ5ccS9EhkdMiCq71UcvaMK830RsJP3N
ry8rvb5QO5Ec9YhRZqWU3WsnVCJR3iGAHuQJVGgPE3iQeEtC5ed1sPHZ8ty3DcSDO7DhLIrIEC2V
sJOn1TeVEULWh2KCLxTHX9lL8EdIpEImhfKK+F/wJdwSGz3s3kBZUfE7nPykO0bZGGQC12F4YCin
ZAaTnfCae/MTJ87gwY//P/0kGCeQ5WV19nFW8u4ZxxMldigX0tDBLMcyX+gO657euoMBvLChKZCx
3eFv337lv4/C3j2nZPO10kA1bTmKkQNjEqxqcB7B216XS5G1DBAlRMZ9r/g+IhtCCFuGstKVMP51
od690noW9ApOi5cIa2GIUrqf7IXTI8TcMpoGjkKGTBnyRIIUFpD09KzJf2Y6afJ8VMmRz6aLoKoP
u2iz5UEeS8eD1entEoKKpjChuOhe5GWgT87XEEz/q7G0SyI+hdTiMj+hQ2Iv5P41eBgHjNlqxC9+
7Kl0dfRdoH/MmQqJ6Fw/tUUOcY34Byv3ixqw5YYEE+/Hi+pPfGlzRXXtPBdWZt4XFUBlU0vFg8zP
UGrskAP1QAub+NvlYS7/E6wny/dad3HSUbPlfi6+vt+o7E3v1K64xNU3BHzDjs2k2xPMetSBOQVQ
9QLLZmX4/oDohZkDAE7MVduKrCGBkubPbwLLUes+1NLT5ARLhvpVdX7AzRaJMqCjlisSPYiqaRhO
gDIovEXf5S1AvcKa+hbArj8r9g20sZiHgwr/h0fdjxmFcYZ6rPWxmxEEKmB1fL6V182wqSzLJ2Iv
+AOtQGnzntmA3uFX0iH6FJbrYVFY/pDPI26gWrOtoen5ZcG9B7JwSiwd1vonwv7ftDT4Ji0LjW8f
HtDfw9DFDIAeWsm/PeMD4dOomHKborgXX9epyD4ec6q13v6j/9JzjOzx7an6179cD2vZwRKxqsdE
0a60Yd3or2KNeLIbcCfEc3CatL85/H3FVsonKIMFQuKy2pwF5QRX2QJg2qEbL4Pocm5usb5fJV8t
fzDdl3+owCTf6zVoBhBQPwYulLHqxeKobEbEQFGGVNWxlXao7vREK8uqUPVgQHrNFutm0Im1kZYF
ab/8SC7L7gyBng4kLADcNHulqpfan4BgR0HmGQEKPrLUHDLYBzFobnX9TNmIylSf2ljpsoC4Wdhg
oBFiczrnAZ7eBVQlxTSrQtSPbjuSFN4d9AnWGtbaNqLwdY4e7YdyKaWbyGPoTvRykVeIc3lSAynS
pYvffxaGK21yYu5dG8Rvo0MyEgoocPl8RTf+dIoGTvUPk/01lhWIXoIsLLqMT69R8T/MUSf17HEN
9L+qInQSiTbeRd9cJ35bqYoUXpwvcgJhtdhKPdUXPLtWAl5682E4Mu3XnQJ/hhK8gozK0cLki/Q+
y0vw4YhaAia42KQmxRyo/j4h9Qtjs0B73AQZ+4POzKcAvdw9xjFI/SP/zH6poq+l4hC1EcrN8QCD
x42yyZ7+wMhV9jm4XlB9G3wDv9TsjfQimi1b7r/GVM7hbx02F6Wk037s/sO8dfvS2Vi6/h9Hra05
TXfIZ5Cub8m4lTIbhv2eFbeQmkaUXPliXJVVHJ12lR7Mzm4l6Iml8Lcvn7kQhpsTao3GaEmPLhW5
Dk46uMQqF3geyya7UypLXlkTE8qD8vYILIHTqYZ3y9+WC60AJtHjUSyohDEKDtRe6VuZptY1RLg6
pgZDf278oy9zDz3aodj8tyiN1xQ/9GJXA3nmbilgFote+jULnW95H0suiTPMWPgRfUsoTxmCYpq3
66J3ftI200FAVCUEz8e9GVeeZMKjaFqcDKOCheCCq/FrX+aFJhhllKPB10tVDzhUsIvxawPheSph
wdMrksByKMvuGsrLkC7KxxhitayLrzCiLdP8vK0KRWsxIQxjvsnWfDYNErMmWpnkLcEiQCjy8a/t
UdJwIYd6USAFv8UaFh44GAYViN3zC6O7gZ2RRTwsdqewthH8bcsyxPYVGxZ85gAmr92fmu0ONtEP
miXwOfiq+YqvzZ47SObCXx4mCRfHxEVomlmWbZoO3KN5aUdg2sDDXZa4QD5i9dsHcj8eSVJ6ol03
JeYgkf1f3XG5lU6X4txLc90vapc+sj7Yd8dOLHuUsoPrtocHZgRgRfPOQDBAXx5aplEEYmXoR2rr
7I9lEsyNBuHeMu9XkB9mYn864L4v3wJIt0mg3iCFOeXmP91YwgbAlP+kRlG9e1RS4DiCFoSQXpSl
lcnKjkI+5YLjw4FveyIVqt3SDqoMuioXqXaIB1xswCBaho0HXELhgvq1EIkY1IJVEJz01cpQyKeD
vjctdTfwbRNLRfCF2Mk89Bgp3jcvtsEbn0NO8Ik2Uc4c6EPbUEo5Rv02Wsas1Y8wggHR5B/e95+q
7Rlo0nAkd5IWPYwavdXx9L0jOy55bncxKj/oQhDErqF6XxTGrqoKgCKUsdLCKLrTkKmYFLsOmYAG
NJnbgICTeomNqxSu+XEui4k7ZSH/+hvmVxsMk1hRyYnCDl2gPIYo9SQP5alaQdZRlrEXFyEoGKFC
t4SxTibOoJgnlid1Zhgn9Ji0phD5lUH68mRpLrzea6r4GjEVE1uUK88hxqiDAfGhKrATfLtb25KG
2b++vmvcAg4MGGZzwShMGmqTGmHmP4Tx7OGmziXo4h/xNU0BYT4G+nWzwN3fjx1pv2Pf8Di8Ghli
c2To5ixdXleGIzbqH+N5BBWad6ylMNkJ8n2BjjMaE6LmK0418x5HpJVToAkneONGyL37UAr4jMys
lRCJIUZxdRsJbKKaMOPUR2brcvd8bP4o0Zo3WQuDIPJFv9DnAZARVjTkQDnMA15PkxLCdApqnlbS
gDdi+pDKKKHjCNp3Zy/gDJtZsqzMIcWZf6brjUy9EKKFFrq2Ta63UJkVdKWv4Djw2KWOpoJpIacK
2LplsBGF7WC5jW7s7CBW9+Dqao3+1ex5heWiONl9GVvCjGz+1B9XYbjbsNbP1e/PO5bpaTnm261D
X/Uptxr4wJLbBDOubJsEEHBCYDH4eMSYKFnBfvdonEeO7BzKNjx1LD8heqB9AZHyXlBelnht2s1R
IveStp9FY+0ZAopEhzRqMm9xABfbKDoEw5sdm6vKF25hFFWMfx8r1HIfz9hKT9rXssb2FnSaTtZC
Wy7ftXn6ezWN1rokuuGHQxpkbfYhAYwplchlXun0blisTLDGeL+49yb9YxSGUkbUvIsEaGv9xSoE
HalqAUzp0j7n2rj2XvD8qPLwfmsLTBlwUY+2DkZxH9A8h8cuf9tuQDP7R2dlCqB0cFbnFCdKDKLp
WYRrT9Rcg+17gQ8JVafHGXobVsEKFbrqNC2T+z2OZ1FYmwUOYMMGQwxD7u07sAK287hLU6deyRYU
iNdR4lhb3MZPvcKvSkmLdXss5H9npQR3xecstN6xLuCIor/OauS1sydXf+RMaDxt/NlsSH6xO8US
2uP5QekpxQEz6fvpc5ycgsB8K2sY56jO1qAEUIiGYY5Hmwup/nBUbojlKXE6YLHlvrWCRVxujxFT
UUw7xMZTjm7M9UnrMfSxK7yJbyAHw2ZorvwK1EOYDMx9/yn9ee90dGaqytkiAXioJdTSNJzz8dR8
A/uzeTnPmpWBiI/aK6tqU8X46BeRKNJ54Nc07b9twxln2kioVmY5n+EnGgKT5IO8kscM+ngV6xww
ByNH+0bZLMdXwYjk9fDrbzXTWsFFYS/7oZanyHysUhMT13nt0OwTykyOkv2Nv6CmNvd4yxC/aKH+
bBzvmdC2mpmN6urg5Je8YnArMI5F2c2A4HuR8BmK0ZAHIPPyZG8Mq+kmLTJd44cb9nI78mGQ0tdo
7OiF0PplhNejXPw7JfzpEuwY/+QouI2QjpUaP+FUq3v3DfGcKuEfGBnfuLBfVUtTr8oexG2kQHhX
ZrYwxmhl0qkYP+IR8lH0DfS5liuEdMoEcxlIDThxXRwfGXIw4xgw2/wnSPBjRqLoAHtFj1cjx4O6
WDsJZn6r0YTcq0M/Zy9TTyCyCCJ7e49hCnSA5wUeKtng5zOZHKenauodw/TbOlBrSQvf7c2K1GJ5
Yw8ahhv2uu+XyBiHUgmH5GF+0bErZuhH5lcHIqxqG/TOY5HzAeWRsfand27DLboe1W9lMiklXrsJ
0YN7Mgvmu8UqQNtpC+kFQW08Polyn8ytiG6/MorbGWjZMdOCsibpYOkhGzINxBgi8yW+5tsgi2En
UOqnCmwMnxMMecOKfzeupDzdPAh+YQ0NHLYaLF/eb4NVcU9nTaZfL0xyahW4WNcBhhWs/WQ4W8IC
2PG5SdNxIW6iKBbcl8JeHWg4gm4g5qtYwJR6+cdIWSbDf+ylWsBI3yxHr2KyAZ5bIjjNFpO7Yh0y
U4SErYXSrv870Lw2bsbPodM30/ewoYyivGDOpUqEFFzkq2dSRBCIdKrOzENqe0rxwAQn9O1Qs44K
orpyAxXZSTPfiCtvw1fIxuRzGLIEc/QhZ6LpYMtKT7nRgh3CJbUsyPVCHKUXWuZsl/JW+UlerGxr
ksHcuVtu9oTy7a+yfZ93swRYc+tlbsVr/CYhT/z43RzyuxR6VOofxoQrSEuvIn7Ur4GkNGEpC4vP
yKlr7sGT2tQiY713UGyJp8x1sSBpdF8hrAbbCc0u3UDKGz8ASR21fmkZegD8gwQSb0zJK+91bGHc
mD1F59M28KDjelbOtuk0J/wZzBMZK9NuwhRVTvvRWu9DcSz1HwYxJBLyv8cEGYyDBbi/N03ndnwh
SJFlz5Axg8sgdQ1lIRjd0pEUE0eXORQ5mtO7kSPYAi3+LBO37dYXZsu2V22DEF42e0w9pIQDk/kR
vy1JLWtXHTJcNZOT/54b/Z4+kwnEYwYY5m6Lk426qVb4foyJWegnnutsIa29CRh0njUFLbWtw5/I
UZl7kXzN7cpbCZlK6B3ottfcpIpxlFCROqm9nMSUWL/4LjhBj5ax6EmvBI5gm3DK5oHukGd+xQUe
ce6PdvVDttELj9jAI8g+3SyriytVEUDAnIx9vlmQMqRUH000tHwTkteBqTs6E6FZuQtXd++urUln
H921nzgAim7fFNJKhIlg5zvYGlJDbNC/ZFB/GB/vBsRygkMtI0CiFfFud6VYrk0jApW5x4g52VoN
4KVyy9+XUZ6pA9s4AQjdBWbpVl2p+zCBuEYVEVTdc+j70VR8zM9dRwaCUjZnBgU9grwljyhGyp4v
EEnAy85QWXO4A9IeyD3X3v7A+DomYloW9EhIoOFjmTKE353R9NhjtuiO2B4unIz0c/7wwRuJhyE2
lyerzEh72d0mnNtcQmg+a4zPVDX1S6gv/+iNkZOwI4v85aaWzuG/3qgQN+GQvJPlLmX0bv1jBI/o
6kAa5zdNn2uWlY9wUcEgvYFl8m3dJN17wg+sZWf5n01SFbHmC6eCzHpczhEN7AGSN1xAjWEim/2Y
VACoGS6UEWH5FkJEqQhSMOzvMDxRgflpxLSUMJVYzE/e513qWX3SmHXLe3gPWXKZ1vZeqiGA0edI
AYLma2REUzFAMdoNZofGN8jkJq/CrkVxIuiN01+k9lS46BXpeHeBM6mqa7lRyrnFf+obfc/LkOhr
oLZhhGT/uj24RiRdv1hP+++0yYv+6k8+TCFq8yM4GH3YIsOjeoikBFu72t6mKxWDYypdRZWUH0JF
tb+P1A1mbTpcG6TQjdVuZKMBWuL6WOHVrOKrGN84myXAMxR79brqWnO/jWGpCnVzDWCIi9Lf5GMi
UfoB0DmMkTcES3MsS/4ag7jMDrIVB+N7MWShXmeNwAMu9wzn3jEAlH2PdWrD9wmuRT7adjUhxNhb
QyYS5GymAAvCupKETySk0kqsa6gFC13iJyDkc/cE3hee0SFkhhSL6zT6gp9j8TWo/PFUeh0cQAl5
8JLl/7qKSEf1/UlX/owwu33HU/37QC+fAqq6mFgKwZbrZ2duwLTWGSsNMxGPzJljfVaMsgsragoS
8chNlHWHKChYw8cl3Tdv0OOtZjNIA4A+GIocAduWyucAL1sqT+O+Wxpt5PdRYTA4YSxVXJCWqR6+
X6GNMvDpoq9xjSD6JYadQ4rfrORuoUliIdMVZrrjpLEZoRaanL2f87DdFx4FWFASZqfUvzlx/llZ
3F10RC7yd4l6RELqVmdhYcKY1ykcbypdG0PPvrMYEfK5MK69TTjQUz7YE3AI2IF+l7bNEcgzkWTN
+hd4/b4J4tzuNEYGPdTj+p4gvbcbywpy+UDs8bgZDmlegiFPPdD839fEsAjPlB2D5HVpNoon49zk
E+gSulvEtqUHBz6EtbA/nM/VQnbD6Lydc+SiksYPb2QvnIkH27XduQY48FjwAJmWZ7z73nygWLRG
FltvrxkLJTq43uE2R/XBEZTYaVJlChplBa7Yaiak0kZOdG8ASMHH58momg2SiNM82fcO98NgRn5/
pJdVChT062bYslxEbEHabbgecDuI5A9p6Id6KGcC30qSlih/sOs+mvd9UPeIZ4ODIXeb45wOiTn2
a6KYzEDEo+Hr9nJr9F/E4Y4xykDtNtrKJPGFl8MIPvaVS1bkrVniq5DQmNZJK3YLYFnPG3H7Hbi1
eFaXlz/eZuNYqwShzF0tMSJnsEQJMjbdFFC0oCM6R0exFv71enaITXEL0drHKqbc6gohR30oSSdu
mD33cbAQdxNL3OkGBlllKGNiVPHnu1ZNxlpniKR5W+tdpLlPxq5WKi3TWqqi4hcDRnRt6z8MEUoh
hNS/MO7cPhowK4r8wtN7U3CDT4yjLV5Y2/utpBBcNUoNKankIYuJq5Wa1xNx7vAZzsGx8T4uvB2x
cE95RoyPNCO8m5CP687mLjGj/4aSulhQPVwRMTfVnRNhoM7Gf1qFnTOU4R2UDUw4O9C498pkxY9T
5Z3GQev/ubzpM5Kg4naVYY2E8PS8xkR38vsWYw9V4JQp2z3tHhviWjwaSLwoAmIwVffat2gZ48dP
h/tPVRxJ2AJwnrdFvvaoYllX4/qGn7oWugEWm2UVJO7zoTzSPmK4d/jU93TGURdSCYch/kPzjY2H
hTCfTcclv0mkgrH23z3EDnrLOpqg5XD3JAYNEZ26YXgImBZTYWvUnykmuDpUpNxv3Dmte+Cdm/ac
6QLfBvnlnjFZlZZZUVng12nEqoM+nbUPfSvFstoIMPJ82pW8ijLGlLlrTCCNGQlmReUVGemSecmQ
T3LTDENLgBxVSJenY5c8o3oWhEMuMv7aeSn3kr2PIoFVD1WJZFZEor7cvrM2NZbxOCS3e5OOOJ6v
8l8srC6nwe7Rqt4gNWBMT6ZvmPEwAud7KOeOPDFthtcHuOryosdayBKQ11k1lWq+UQyK3PIeJUtO
1u414bVFhgdED3Crj926ko3QOwC6vA9RVQkatpSz5z813oZ1hu6S1qO1QL9BfqimrbRaCFf1YRl8
/3A1S3TVQvC8YPv4gfGzXnMLDe9BfzrhL2uZpFzeJYxYhKD65ahQs4pyefbaCxKoMLpmV+Dz47mY
fDg11ALnjskmSG1Ds/HSRJ2n+OWeB58yCIBGUFcU4j1LXKbl/1RQd5GuxJ1ecL1cUpWLsXP3Uokd
L3mTVcKjv/OZWmXiSq0JS5ePPSZAGvaoZ61cd2L+qFPC+JYYUTNLG9lk3/TFt97rEz73dIWlLqo9
EdjfZWTKpoVx+QBThN5annM6sMQotMarrSC/6Jn8qE999yGacOF0wB1bIh7DtQZ72GQXPmqeCAw/
zZnoMUbJ382p7kAdjvFgY1lSo7bZ+cCPqJERSq4PbMVf2o+2IcBOCFEr+mOZrGI6CbAawV8+C5fb
+eGEOPuMYsMddjd6ciQQ0HTGqEc2QnxBOg59q2tBHJq7Dw1ab7hymot4KfS7s6dZdHv4BF97jxWb
AQcPO3/WEpO+JcaWjc2p00HwV+b0b/lgrdsEnqIvj4jc4iOR0D8rTr+Q8D4VOtkvQAWConLaNhN3
qFEI78tnOaiwXu+fwGzv3WA/5ip50/MHpn9BbDPbSKA+NTaoNizhPjyzdMeReA7Y4b1s3XvotAO/
A04lDy5cluIZPZTJckFDKBe02a6zb/psrdRDhciW9+84mi7U+n71sgtvADhonbFA8zzLcfWzx599
+WRf/voTftm4WYzMkvKIu81rVi8m2kt+bHPFtn8eveWj/el9Mng4rgorZlYxcj1sedb1lDnSdN1l
O1Gez2GWmySrhL8R7+dA+r10Kh04E9Rc1hLFOVkSBK8VpqLAlNB/Bi/Lo2S3Wy/1lcx/6Bkp0O4P
Ys/sjClp8Wgb0Bwbkh3yXyVd3D9+nVoPpNrbDV7HDcs+A3jDrAtrrO1ZkpsaZxycUVMMeD5o6D7/
kHvSdODJWPXpUnxQfvWWh9hZ1gLmRMrigqvnprOXjLSvIJepbsuJPgSTaX3R6XPEHpwaHZJwjvLh
lOSyBsYIJJEYm2CzI8r6DMARAiQkdUjSRxnDrt+BxrfDdStLJoZWOpZBHh5X3YiuRa9tq4y4VsGi
XLajqVfChR1PkdbXrVYpCWF8xoi7AbTpcODYAVZIjTx6Pu3DzlqUAjEZgUZIL8jV6Zfy42LPpeJT
MsNmDu5ltcUL5AF7zkT91qluPeVjDXtB4XdpaN5zTWb9bqyZOp3FgXrTmsxxScLu/Z52uDSFD3v1
Z+b/xtO5CVF1H+j0K+WOAiocEIz6JU128pgo0YTv0nqJymEVr8oJiDi+uulf+P5z0MYW5x4QDgve
mfpTzco3GnkEbOybFKbC8mFO4m3TpEPF/yAdnp2czTm9eMI2DCPv35qHfDGP7ye/aZ70ddbK3yxo
p/ucr2d6BJaOHdx6eKfxZDMTVDV9/p0kNaCIybLvuteAgfXRoBKRpP/DhF8e37lJy2oAcRC0TnI1
OlmG/mvFQZxqOORuKNKub2IqCtM6P1DvnQEhYmzIl/8QkKNcv7lkkpxhUNicQW12p2QrdXWP+U+8
m85P7EmY+b6NCMPSySjBRJgR/OdW8QwUbKpXgnfoWZ5lm6gky3YHea3R61jGcIQcgYHFhE1GzOK1
/uIL/k5frbCT97yw87U8y9cfUMz2KLCPJlfXpIvP+JCrDjVMMWFLfGotLmNf/VMjaWQZN6s8nXXk
dTpDYi0Ue8iaRA97tQsY8IJ+Mfd2cbFRi2EqJrKe+IYuu7EeLV8JqJT50+klJ/obOUO5m8F7K8Q1
mRamG5mAmrNJ012ylk/1GwdG0vs7AvHytQWkBmSjuIXtG+JOeNgoIuW+D+OO6KB5bJ4zRFEQNZST
eMibP+J9UqvgDjAK1B5z7YuqDG4UaEO8uG2OIGGYnLSukZRtbXEYQgYRuRgdVPg9yEIoHp+yXi9p
pfOvSrt9cbx3mF/uBFkYa24ioFBGY9uZQGded07XLHB8aVS9mQn6VlXgLxFQ+hE2toyMH1SH2us0
EMR69CxFhA6EufnduMhnfHVNxwfPoQMGTXL2yWiFFNGWFQK1fveeMG7tUCP+8uNgR2hHLsC3vqk+
7u9XX0kneOam24BZ1dy1DNoWZXSMUy2RDAeT8TaBmraqaBQ2xWWPinGzZYzDS6VOo7qYa/hzRbQl
R8tdWBk2YEdCeNnlhe3/y5QPK6adpFI/agoTd3xUaujgrNDBmG8mCkr+YoruOdZImb85KXrWUsCX
vkHF+Ado4Dy6BkgN2BCd8LKiWaoZVtCIFLmdpMyT1+rmHXUGCONULGxPJpVzX5yVTXZs8jJeS2N2
bN/fZ1ZseYlSEsR3fYKwDMZcu+3GhYROy32JT+KOHTX/rKLlYB5IQvmnPYpIEttxe5UGJZ+9KKCz
BYOzvU5pyuizi7msH/MvS8oojZbMzWxTYWibFDG0zYMx82rZMT0u2Mc8QFV6J4vWpI3FFIqFvzzx
AF+tg6/uifeI2n9pYueSWbQ9QMjgbWm+1XN2uc9HoNKHXWB0nBW6xJXRiwTV+LFNRBPbS8WD2WXR
9iL7BJ0u9maTdlZkUgFVz05tN79RKEUzGRqt4Dp6cbNMJn5bmCoOveifjrhHUcZynvumgP+gTuPU
GP1DMIUQINKPvueb439b2fLR70YEaDC92GwMhzFfjh1JMBxwXXLISSAZSk8O4vcRlR7LgVzfxqcw
+DOWXaNniOVg9p7y5GwOLQuZiMh5vKilGw2QzTUTnSRTzl9RoK8ehxUK4Zwi1z0HqIusgtBmUqD4
Xlsromyb8xSTTfphDwjavsMthC/rFZCNO9nNyWUdMKPljCf/I1ssoCBjeH5rAvFYwuVIGnZI5AHA
NUy/oF58/DJNdCCC28JrEtjnC/ZSYEtt8D3LY4bS5CgQzKwz8udF850Gy+TNcKYm364xLE0GG1sv
lyHbBNoJPHDJHSEMAfhhFrZf3FSDLU6NeHaQDfD7UsNM6NycKq2YpXZz6nG/L0rCFDzkDujoYc7j
u37MU1Uivo4jpaxXbpLWospTpYPrqzVzhW5FrfE3xbuNZ1Io+KWCrpoXYAOpj++WEsWOki58UuK9
jmSIht0N1ZFRYXaOSoOZxFjV+Fvj7j/MbJ+EKmy2b9c5SV1j2zPIXXOWHm2L4bKQ/6XSCLYt4T5F
BzV4Kc6nmKDY83YDzWlSdRkuGaRWsrPDMoBksTFOGnifM7zsP8ZJLC5igvXcmJRZg0jppN/IAH/O
dZlG0CATfea0mLYImt4zAFEIFFeRKrx8fxv5UP7HnTal/BV8gX/2vPv6EE30XLSICs4sicE0SZze
T3FLENfXPDM2RoTO20CXlYIaHrCk7HCcq/igf0rNU+jyGMFyPD94LGRkvR0L6Y82V6kd87B72rz6
XKzgfsFxgyglxDg+aoSgoNzc+dVsWxWFrfZMVd4cwSWXGrExbF4hFXNa3X3bOSq8rH0BhPYSPIS6
wWm1N7ZnYymtU89KjTMAg8BrGMmjtUvetVcON3ymdaDQrSkonhBWvA0nozR7fbZkb83H0z2gn9AH
X4W05CIFn0oROswRFmDRPg/yvFo9+M/sRIHOtCiPJE+zCNi+3DVBgKlZ/Ww76FXOwAFJgq5l2+js
gS6vE/x9t+OkW8OTmEPgYN/+GgPrf0lpSAbVnnRKNLcvQSCWwDom4Kzm4PTQfEkfBqnQ3XXRwRgB
ef/vBRVvQx6a1/nF5RdK2x361pLVPpQ+O0W+WATL2iCOQcziuqMTPSrs4ahomMpXkySqDG8fCb0k
zYC8AAZIsTuTfwPf6i7IOXYGhx4pRQdpE7xtwkcsz+AzSGctYJblW3G9zakiKb8GNtZZGOl7Al9V
nJBKqaTsY1oMxhCB8YbKRflEa6jeQ3GvPoPh0brUw1QT67yu/PTztNJhCwrxT2LJwqyKo4tGgeIy
xHHXn0eePISATHjEts7Aw5RTlk5OutSt86QGX2kQhNEPRlu2S45fe5vHH0ZwHAinj3kBr5R7WCgu
y3Q8dERwIsuicwBSQi0CKaaj2u8bc+9mf5Ldehej+7hLjcTuJBeGSmFY7FP4geGS/kQ2bFCCXcdC
9FEvLys+ttteUv9jOTpHIkFJ1Hn4Il0N2tMqCbTxDRomV0p4FRYS1+p9d/vbgVPW5EPGQJMTeS4I
Q1h4b8nD6Jnym/5vdgctwsYsAYKc9lVkd/66/I8ykPczYADdLA9jycxmOGALRAwGib0atUP6yC/J
BHU/QEGseBuinKZauTNFw889LJs/8oy56aob7c1+YQray/9lOHexhSQ0MNiAyP2LiL9hEy2rdFfH
NhBEwoPKdMeE9czBf4tdVlftYSZ/sJPZJA5rUSeyOiHrcoyY59r1OKzzU+4KnawvsF0gQ3iXeT4+
rI7EXCvn75NKOHHKBdWJhrcVZWNAZNVvdCXkkbpiRh9lf160rzg1edDaALwF8SJEeqwnQQGCrdWu
bES2Q2t/QPL0KMuXssAHkG0FzHU17Pf+2tWrigu7Ig17QGMt2smc8EBv3c4jvNnRDzWLX4KjN901
6cG3mNZS31v4UaXb5JXOzXPSo9OLd4kTR62HIAXupnp7qsk4y/7ppEYt1rhktTE2bEDSrcHtrpr2
ZQrh0nxSr6jUWRJpZungu3PH2XIBOab3GHjV0Bxys85h6oi9mDxhAuPQtNLIr9LA8fUhzuaVsksb
i8f+ibBTJCE97ht4hxHJHyFyi1Px1iyVb8GxLmf9ZfK2iYD0M+MMbQzD+J/Z9+B6LHrFbqDdleFp
/AuSrnBjDpbDzNhOZlpXNwJJpOIfQY3Adfv4V3BmKYFk7dc+ZUhfhSz3dgKOTZZf+X/lB2HUeLTI
p6Uk2dFN5a9+K6C17NHHQcIQoUJI0Y8ANUVE6u5bUSaSPEQqyPeY3YeNkcjYdvKoMQcxdawYR8Po
+0mm03A8sNQU/gFehu8D+PjfuOIGTk9RFEXPZr25WJ6utOxwmGzUXXZu1fjaRY098La3GZ/XkBe+
ZbLMFnZsDeggw3JCYDhbVcd1FJ3x1exLbB94qmb/imOQA7fdwVbe8HaG2jV4fOCUW7Ki9/H0eG5B
BJj5JjX/j4l7Uag4VqkLXYoUC9t1lbIXkaDXi+gBrNwYB6473bwEMfAGn0Ax4AG1xexLSxLBQFLm
sGzol/5/kFaDFoc895DItlJ1Kl8GM6NWoVubu1ZzsCsytThrJvk6yhI8G3T1Q0N8yqVREKrau4rN
atTyNLjVhHZAGKaywU1ONziZLTE2PFMWLaqv45ja4OVzozwVmF6ghM7ka8z9YWwkCQdPODj6koFj
SMi9ak1uqNM3WDN1DGc+LYwF1f/kAJ7CLSWtsBbVyihUXssZug8cPyg3nOM5kZ505uXqdnmSPPSZ
UNFzrCe++gMN5zdNyufH//FYqL3/rDl1/ybtoYBHF7WzXX0XH0orlmlk4Qm2c5CoITnEgAXMA/vF
za2FvIFKCHG1E7J1A29rLnnzx1+Zy+K2WoRJFJlqzcZ8pZe/rXK/SJcEwwegXZ/qm3h/YOhEe6vL
zobdrRnKcDSDlSdIy//TWLc24cb6nc5L3EDpHwO1fMQX2WLxj01W+rP4bmG2dM2AKlpLD7nswT0r
dw2W5ECu7AK7uoVNb1oFgUtxQFgwmZvH7uAiaVRqAzyMy4fo6z16Tmt6kCFSW5P+uQ9/CheOmfZ+
DD4GSDvb/RDOv6BvNlCAwBfZS9keBHtOMuWVZNq8swiGE6L+dlz/HmRhf5eifdQLbKsncaiO0sO4
XqmZee+fgc4ONQnZJM8PSzBD+5/cgXWX9KQ6Jfk7owWgvm0DoBjnRzyPDyuN3GEkdB/d17ISJMVT
8bn+Nw74uw779ShT/kqWZ9KfW4KK5phIH1tSO56S91DeQIQyumPFikFvobaJCJ+bn8dIjaKC/9bw
eMl5s9Un1GZtDf5IqplMOdTC6ehfdqZeQFT9xxK2+rMoXoSKBazxbT0p1xh5pt/Jrfid1mPWDg8R
vBj4tQtbtIEmxUswRNBS55XHhuIYeCIm96eMmdHcaQz0Yg9HaKsOvzdN6dxR/nRfCFqy3/UHjrFO
eaXrolbUrYWN+AV4XOqGqqRD9OwUXtVCsebYu+cyWZJlEEzVKocDZHkC5edgf+dqXSK7Ib26+aiX
UQt3S/a6EclBa+xKbzVqpWUs130xJ2sJfJ44iiyE/lDGkymKwXau8WZo2vfZRaoOb+RQnfsmMRzD
+4/k9XhWMrHSTUa5oPItH/bzlAR3IxWWboJVeeoK/nyZFx/PDupte3pLnHfwzycZNFur58Upmr8E
sPsZUr6EnoHX6wpmvCTiGxmndv6RZYVTHaOGKr9kPNx9xcnWNKeqk8x3gkrfNxOSpoS8OaX1ctT8
ELTuCpBqmKi8ZoMmmzrGGVLFOoOb7Ag4n0jhwnbXzfdv73N7K8JhgIRrBQd0kJKUnxTIceebrtco
/2attv45Iu56Ybv7IjkfpWHzH4vTFTiZZDQl02xlyDV2sO2GukcWVs8SZw1ZVSgI4kA0h5ARWhU5
/2rvP/M1q1MoQ/bMCEO2dWFp/VWC7JeHmkqRWQ9V0denzPndOhQwuWuSx5ExcCCOYZDuMzJz7X+I
Qb2qpRfBivVGaJxUrfB8s27AeE/aISQhQpet85yFSP9njioLG7Brbl7O9AJwlPuLrUOsIXyNacAt
FP29W1YzncOkr9UhopyEP9PS1m/ZdT6qn6k6UiiGBXEu1OZr6qmSqwdBhzyViwgj8i6sajNGlurn
vdT4ids9ZdlF/wXjaJUcUs+SIt7pzs5rqouV7jRjDiUQw6uNx8znf8S4XAR1BOfkH+AJ0OnFKtm7
iH0Z2GJTb9LJwwfhnnV795Dd4DY4tn2vLtHnyTfE0EYPDuR4qWpyiszqj4kH/++bceulEk1A4SB8
CvzoDMTLeDBjTC5YSp15hhAm+UKaSLf2m+SIpc/dM/YmsbUXtPdwmpXu2HI5gQzUKWRRXkurXgr/
AYgujvkuQDXx2dK4JltPoTnFunYJ1ZLvIJB/2+0KL7b7eNaH4droleTO1hboESDzkw//vk8Z5kkY
ImkuTFDgL0NGnjj9TFgNqLy1h6ch5ftMYweWRU/iXxBupocqV3aomJgz64cKF5H+WOUUGXDFLoh4
eBz0yQaiawA7fifagUkS5vya3DIsAY2bZB2pVNmZDBtgOegf98zXCBClW7F0V+NkRJf8h6NicHVI
hBiaGfaGrXXjlxC4xnH95LoVEA3498mCH64cSU46xW5x48k67F6We6yB9oNIc2bQYXmun2rckUG4
yVzb9VsN54+gamg7o26a5gDeHspwwOWH3P1bDqx8Cb6jidw7gzJKTkdEKkXKtK9LZBSoEKZ7TRyT
7YEKte1ZjhbMh103y647ObEnycu0ju/Un7/Rv5eY3p9hHTk46JBXobxgAMGwOD4m9qvdmHpyMTtD
GGOD/aW90h1y/7sl7JldS74yaxP8IZnHtrlK+rDmqn9oDRmtQAyfOLcVVSSjb23tNCAL8bXGUeRf
gIVYiVQuhPVVgSx5UUusUqH9xGA/tHGIPjW/VjhGhu5YcNJ2mk1FAtGe0SeigIKNNOcKoelOefOo
VkvacTxUyrbELkZC0p17/lGu3G5/vgGCi/IZYOwC+oYkzaTsBUvThgzOiqPjeg2E1N503tnCZjVl
cw91pmF7lKQz56DFI3B+44T7q4sb186LUjyTWwoUfFM446zM3+Y6QhWGYZfZZJXM2DBBxveKPt1s
9WZcmYJptjZOdSUnQMffFuE3SmSp3v5P68gyRF97moerqX0U0ZhJASGR2hKlPOxa5/XvYn0ke+/L
wwtxRFE4npvYoMzWYsVVHDTQQnYKeGuZf6isaQ6fTPIMDgC4AuSQbIRWKux+WxAnxWH6n4mDAKK8
DmiIBWeBNWZNZ2impq2ihDuHPQ0BFsr/qSfGYL+QCHxZ/Qkv823Fcz3r5bYMnfMp6/Wa8eHurBtw
VYip7yCqAebYd1bBVpvhXNF+8o2LJlhcWf0Y7imQJeRUL9yQ0zkH0F+b+6tAnJr6Ba7IpSlX3R2u
8vTQCg0cMgQ7V7K4YBEtZF4ulHdZHUeCmqqRwQANHstl5+f+j0RoqGAZYhsA3s11RTQvTVpXjMku
r8wUaJ0F06YqvbBM1+tjQNRVAq1jMzpo0tdLqRvjghCCn+q5zZf/YLIoP+agmW5qvbX3KySUDN5j
4IPSwuuOHasFhXGGCpf0GYodin0+ZvyO/8A63oLAS0FdDYhME7zsOsG0GtpXWVSrTnh3khl3JUjp
0tlaZECGqaS56chM+MeyhX3H8Pd7P8xSCh+j7vaSVdU4gMroZlVID6S+rZLRUmBeNsY6Fr/xBFMb
R4OxsloB61Pznh5vV1fyTFmA/ol2GCk3pakdsu0dr7KN5H4Mn6a5SFGITOVkOowVQwGhUMAATbVU
H/BG7HKAqO+Q5OFGCz8Y7epWd/kPDZ+iebf3ZSPri/yF6ZQk0JtK3GDWyXH11w1Oisp2vcqjhHz/
+Jb1YdCmXuFnJLFXTVX8fm3Fv/N52LWxYiGqAinb63/0/xYxuvtyKsBLLqfys7lPMKTRYBLaud/F
Q56GLnsCKr8+xzq5AFeC9XOJ73O0FM/Yym5SUS1skLG7dsxJFwIj/8wq+Ksl6K6eDPu+0kg0xPf5
7oytgkpd0taTxv5gzpcdZ0CXLyRIzW4M49WAakPs0ioA5mDCGhMfq4k8g5dhEBOJImzfZoC+oYl5
0+HGaZNVxJ0yIGtg0paLu1lfTTR7A7PqrVdqctHIff1Y5EIzhalgf+DFzrUr9SCpJvmME318Puo8
5QqizQgB7OeX5U72PMQyVcVIzWeipwqz9KzKvnsEi8uJIZoxjq1R2TfH9RGBalRfWzSDAlnPMIdh
BBjVTRr+Pd/N4MRK2uOAJEhHwvg7OXSIPjQG1d+dDgrBYQ96UJ17mMM/rxl9BlQirAhuULxK6fmn
2dM/egN8oWtiCqRx3MCD3PodaOWpIPLxsHiq36KZs0H8/d8VtEwaJVEWNGXWZk8l3fkMIrZ+iZou
ZfYz6VMFHOE9irM4vdIircsYhCFyF/T5MltbwCT+1w8Bru8exrlMYcIYTkLoYyZEv9Ui9O4YXu3h
26ZXnlWxYRvyob52T9LbhggACv5dwmT8PvBA3JHnTl+YdwenUQIzynupOlaZlCoAAlwG2tJ5Qy78
JSFQJG08brTwbNOPNRG/O1zDUpCPf3NGUStoMYjExDngXFllQIXWlBKDUDwpYz+B2PhLTpU0h/M+
G7ZrmW9E5gTNCzlCJmgXNEhpFyvH9uLbn23cUhnWZpJwQvx/+2H66hxjJrzsmZfYnQwTHXXDL71q
RkkDdnsiR2RfLJuF+rRwnWTEWEeEDFKV3+wWVLUBPr+asVN621kdyluszVHzO5B1CoDtE69macTf
1lYlhW4QB4lFXox79gLNpj7bXq7MTG2XgfD/c4+qbPG0ArNaBlPd3Bkd9vTU+zgDQGV6sWOddrg0
SeohMKbO3eeP4B/N1oZQ9qtUnEpt8qVIVdCjB4XkIfRKPPnzks7NGXoAuLC22LDuAQAzGhvgOR9/
j39LwLCZVrfGWyTCRvJVaNC8R3q9AuWX++MrCTBtypB0TAs5h1BjUhXwdtHcv2Zo1tKCDC1L8/ai
OGujCrWyZxpSQ0RogcmH+DMNYjArmYAPZE9SzJP2h+033pFssI9RWVgIWDMWEk7AvmmzrkdGqu7t
uX/eebzFobd8KdmnJgV+IWfJdv09zKKCOCfODuw2n7VD3STeZHVxpkf67Mwj3OAKgBaeOtQFimRC
sqBaOgyHUUaR/aTQM113N9wsBIDUfJ4B2RTUXFX6em4QAT/XI46lCrTydeRbjHU3qVxvpNPe2aA6
Qu2zlIBpbRGHBjOzHagdRZ1jeqQ4q69RAgCJSro4EI+OJLQ+D6AuC6TmMd+YNXtQPx2W+BY87MrP
Pz0B2MKIsRQH+VEpJeRfjHKx59pB4GTjGejFtnFAt3JMfGpsgsJjWziiBbdrX3W0ndoqxsSK7J3A
ovKVv+Pma/vKRahUMNrcP3AUh5Kuep3LQ9PyM4qbgpWZWvQE043VdVs/HX2yYXgB2h1YOp0XOt/5
BbPM5BeSUfbi5Ih3xgfNQ9EWldQAG406zFDKhjeNrk6ka4clhgI4Y2JTClZB/EuSXsU5YYRhRkEG
zuzLIMrHV+SA3cw0nG5ereLSTIuZdIJc6ncFSN/WJnXYQI9YzBV+73+as47z1y8UeATArLx+rTg9
J8Wde6GLpB52lf6SENV0nj+n2IqN9PJgdT9ih2FoQ6oaiWSdJL/cRuR5sbOwRoCER1sPTvs2O807
MtYKNhqGa35K7vMkZBexIeHXv4Uuojn89C4NjINKUExOBDRqGW8D662oufDNb6Gke1mKoC+jrd+S
EX1uAliAxVco973CFk4Y9VJMPwaIKBnPimBC34qVZdWS3cTbFSXnm2MGGI0GVhRSLQ98KA2iFwOJ
ikl5Xpl80jshz6dnqTkeX4niFD2tp9e7d/gzBzaIgp2le1SqM/g9QN+waPvhCmUuM/L1u33lZE1y
0XHjgyoj+bhzByS1IWPNK1701RXZnDctugd7iLMRlb3CsQn38E00AKF9i7JHuSwb1unkqwDxyoTe
irkBApbsjFIEgSrr64QPHgLhIJlHCm0IJhXAq7uGmkpeAlbrzUXXcbFnc/H5nq9pqXa2vvjVhBxw
KeyFm/jk/szzu5yHUc2p+CCpPXcJV5B5aLcZSfbkmS+FqSrwbeIxoL3RV6UuGAtBJe256Y2W1ViF
u7fHt1JhN78Ihu4EWo1jkUSmuBA++S3v5xA0eJvRIAcYfw5dE3j6huyoe9zsGJuGP8v9kIo6djVk
J5FpF+ThqfBFAW7U+uTfz26ns/lbV2tIr7uHBg8vOlz5cJOJLDEL52m69uLJLTlDe7lMlPxjWG2r
3RsZPJhZsy4nJAtYUowVs48QGMd4BCnA6NykCaUW+3Mq+BYrHCXPMUOX49yIUAUeLdN/a+rD/2Eu
NVVfgikN5RwYY0q/yU6etKb+7qvnjJnQsKqm8ULsEjmi9Imb4ESuN5MyXMsPNXiXF8YfSkD5BnYm
VzfWltIdE6ejaPEY495jCnUbLo/DCtymHz1WNGbgJs1NumLTdAfhi3kLPZZXjk4Fu67Dr+siYkHq
mPNGIf0NbOsc6gSEtE8DuEyKm3YlaLTuQLACAX7mNa/1lj297uA5Wne+PAELV5f9VouIjH8QIm+B
NoaroygZqQU42/Hc1ODqC3j7R+I5O//70vf94n+LfrOPSU+qiBfbl05Hfu3cUe7BztE8moArxEpw
neGDTmN9J0SBjevUm9R+KAQzHZN+gBgkNsPB+bRyfSkB+yWR6p/zLmKsniHEfaQYtO4YEcYVBs24
UWxb6dGReOTukBljP6MusAXRFIuXZ/7ZIV0HiUCYL+DFX0Tgi6vDry09DpMDghuMFllx2G/jlGF9
BNJgOyHZPTi9zCP3OhWhaA6LDSGUUn537Dw/UVnWOkgdUvhx0WRJU387B8cCk5FwI+dDYVzpE8cK
h5Sw+lfjgsrizVU7YiQMX6VvgG9VFZQeU4ihHmkTiuUPp7yTMYOhTPnYSy9k6thbPY2d1Ta6IoEh
Nhmf3h+rPkQ5I8r1iM0wbY2CaUmbRyLRKMfmqcsWvKrq6vE5srGMyHOss39qKJwyDbqTPGCWMtOO
lrb17TE56trBfBzCSZZuyHErtQXM+mbi051rCw9unVsKwmrgdEHiCycleQpowSDJai0SMJR09vDS
YESMXUnRObTaQbry8KwhRl7IRv+EDtnkNnBugDCJGy8RSVmgvDQCNUR/UciXq9q9tl59SG7Yg2x9
DKud3/mLXz6c5lxJmAenkNgELbWbzUgUqBS8NxxIg+pwDhgJTr/1Hh6MZwYHVDuhImKjzlfl2abU
3MNiTtuCKQ1t1VAgbTDrE1FkmjE755afjSgd8CyxMmZJ3WgYFgiKRHWmRKapFEH5TKheZ2NSSBFi
1r/4njbODhjaTYfIYYrztoXhGn4xDWFps4hqBU0cIwO5BG+09xwZMR6QbunM/AeTYD4U8JW21J8J
QmMupsY2E8Ikqn9xAuURGTyuBsBKMZKHXyKVM2rDe3iUKVNU36my9rq3jguNrbaFF/llRWmaGOrD
m+ZwIcfeZMc8y5V2bBAl8iUwvSOucmb37T7/IXkN1Ac2pHnJjflQqGilSbT+4/dPAUVl+oVk8wnZ
wkZkspWq0CFGYnIt6jLDjELMARZHcm2EbA8SAmg003pxRaxGxaciqwCgcWRe6z5QHF/PnJOuzW3b
Fm/JTuSoBT1WqhTxa2xkvvdyTBh2FdTod45DnZExO5thUXwldJXtVO2vYV3YlpeQiuJAU/8gjoUy
E1cKXxh2h0EJwFPRtMm/DXlvF9OpeLQ4zfRgCCGHKH5WqE7lOBMIb96VXmOsVGuF84onp7ctX4vG
lJXAC2K5dpO4NllClBw0He1H1lzXVr8Ra+iuOq2ZIqWSTVhdBMTquJBUyBBd/H1ZDqu4hWfOQHhj
gPCzOzY881E8i4A1gXJxdcM0QtHlad1x9Bol5ueY1KDOrK+yA3C9hOyvVK2u31kgOCz+siPo0G+j
k45s7uOFYAskQWym+A3CxVHrnkMQk4UZoIrujo713hUMgRjtB2PpPMOF+mapJdQB2ibL+C1gZVz+
5FpsNuSCq1puw8TuUbAnsQxOwZFlN88VDSN+D9mVdtRfJyA71nv0vJNTYdrFVd78vxC/06dDjByX
HZDNl6tmN6gWRV3tM3j7qZgT58MCKuggR2sltYJ7PIrv5EdfFRKsgXQuCH1kDtjMVPHIo7Z4XBbj
cLA+K6aOg1kzCq2u7qZnrvu/1DbVCVcit52H7PZ6Gdhm0hQR6jls0yhbXznWiHy2rbhd6xk5tTyM
z9E4HkZBmwRffN5hM8n6f6ulAPJZe4ZWeC0WtCajfWel84o2pVQIh//KoD5eLLSga3rnVu25TqZn
C+D0EVpjURKUuKnBmEuEa7d+slbEDDxEhzKoku50PcUClLuFYqpNt1ya9e1EWNR+chzMwIMdSX3o
rHnU3zASRzhPLJs/EcfLJLjn+FxOaiYo1JmoY8sXRL80ABGtSvtrwfHrR+NFqt22EQBZEIqsGxlZ
1QbtQvYNOhxxxM9xOBPVWorgKXnVe+YHpH42D+PgiVZo/sFw/jfzDRemAstQ7sGvzT1Kv9qHp618
pJaDPEF9t6syZ9yXZ8h5//tcrLkf1ZXqYYUoBL8Yz4DcTPeGiAwUjoLPgLWpy0t+pi1Cfta5mV58
42RSruf9AMPz1RUQ4u4mwa/JVblcLAS7LtL97deqwuWl/84a1kr6f4oLafw2TJKkkuta6FFh+aON
fkX1sgMiTsxYdFCtZzdTh2j9KjZZCXK2q2t7nLRPPNw92DgKY4/QdU7rD+b92BxonIVWSLOy9plT
6EMEW76qH1oLULeSMOzOGtNViqjoiWUlSEIGfjv8clfoey1dPkIOKhwx+zWLO49ep+jnDmgRuCdl
krTQ2Q+l2pNVvENgtMrMTr2Jye2k09G31btOvKDX2Qxs+rImj1cH5NnldtFavB6hAMO2pT4oVBMa
uqxG0AxhgUqOrjicmU6acf75jkCxsIOapcIPmZXs82FJCtYTenJmYrb1mTqTzw/m/fmIbHNdArUJ
Qi/8RtXpzk8v2DQ/m+ucIbiB2eJ3oNMlCTIoY/KnR1KFlG8nqkmd/kUNsUDKeK2+3XMfwUqWTP+l
djzftiEPRsGKI2Zo2zRqhFAFzSU+zSJoRys6mNzgprLz4gMuYY03LilUGKUv1HV5S0fMvt2ToQnr
3skjmqJH3C0PQM+ggXQ/kEaVzzF8J7wEgVpsBsKdqgkysf2KF9gV0pAghVJJVFOOZ5dPr77hIfAq
KTRZMwioG1ey6l50P7uG88aa0v8917cobVU0n3EQImtefNAXxkN684LI3AZrv2tlrDJeEle2AFT+
PXGaKRwxHwN/LjT3v8hEQTpjH1D6/ZINtOwN6bD21/tuuRB3OhBedpC9NownZFuikT4Lu0hfyPFI
AzJ3A24GqPFTNC8OhBfg9oaRWZ9UKgm/bL5ujV+fJPi99f80fBxSncwoW4XVgpO2QhYe60/GJTM+
NZ/fU7YbrVGuiBlV4SR7EPH6mBVnLQwkwMBrVVyY3S9UqwlSnQE8g57hly2n0QaE8mXIFPRx74b5
LgtwMjudhXedE8OKCBaqP3TD2xL4bC9DkoAN+s/VnBLoWqaKuarV6YXJF5pDmbe82S9Un9fgAMqh
9q29RJo/TZbwTPa7MCz+orybvvEXoR5g7gVQqH8k+YaVcgXCUHjmoE6bTH2pey3f4mOehPKSsXOk
GGzUODJU0o8U0BO+BMcHXlHJK7kNpNueiChDWU36aGezrRWdvKhi3omUYziGaCM5gMjdYG6hvZaE
Yv8+ci3ic5zQpwvebqmfpfseE564X4Ht7jmDfAgwzOsKn+n/ZC1u6NlccdjUozGe00pRqJfkbz8E
mtTaZqeilN4FpJDQpsXDgGO7q+B1Qg8827CDB/tkg37NfbZltQ6kxWx9P12ToRmz1fbAOG2x4i+F
UPEWXeK0SuiwCWuBoaPWKHzUbfeVl5Sd4VFyhoZtQ4cmBZTSirfH3XvIxID+C43xTy2HP0Ez4KMv
UvdBDDz0MOs06q5uqMCoiGhOT8ElCclWAlt20MCORgiDTltT8u3567mq1uRwb5JmlP9w4YgT9Uwz
53KDQgb8rXUgcQWbhxuU7S092AX2kA1ZpUWEWuM6WvZedDTCn3Drh79DBvA47jNYhzyoZnZxTufG
YPSPuqubTzeNPphdRNyyUjfMJYHygrfcU39tAX4I0J2A7Ey0vAgTGvlFtYy3t4Vas8NJ09F6wDzX
IUmb8W0Iok3+77l1wBQY01iYn0DICgZMOcGxIrOJXDXWwNreh9p+1qhvt8UnxOpbzmJ46xiV2db7
+RywPYBA37CWzax2z2N5DA0jyqVbrJbjP5IpWnH72supXhz83Va6LOq/cUG1eD5uO6PpHTKIjPly
7Xf0TGw4xicMtKu4Ny34IgtGcExdA0iAypshQSpdgQkfYw4NCjvcl2vc/B7QMjVQDSL7F7Yzyg60
dLtjTH4vFC3Nd3K9U3DWr1YhsPArxQj0cWnJT5YR3/tJvt88GX/2hWeDwi2CGiXGhT0ncJsvaalH
++X+dxPXe8tryuDBQTEwsNQOI5j3uXpFaEwyEWWdMblvEZiQ762GKWS7m5/kUn0U3m+PfazT+JKM
JntXy1kHGWI8ji8Fak6oylwVL59abyih2HB8xymg3vUwLG+e3Ru6d+0mUoTX1QN7VnvdTDb0gbZ9
ZJGju5vyXwcwuk2N7Rl//4Qrx8VX6xcQPgmtr3qf66qu9TyG6MIvfrxpqIwUcVV95AWRA8d3t8nG
5sru6FZofUsccVRxUCdY7GXsh+L1p57xI6s8FpvBN9e8/QJPWLharmxb1xd8rGNm5RGF+qZL/VvL
EdFbeucZ7F950dip0ZtNTaYWvkx2IFJcX6MqIjflJi/E8i0nFdZxEMnWYvNDg2DBntDJJPboqYIc
17r5pHl7UmDVEMPdfkJPveG7fMPtOJsvqL4ZUsoYtgeUrM5SSgVusJ7mzLUBaa2aEKQ1Fhm4wiMq
Gls7pT6PUU1eTjuJGXRAHPPeSxAH2Jw/L84g0Rb42fnPVNq8zUbjbBka2pLNFbSofhZ8hhB2McGZ
6D+C0AKMlt45sXvs6G7lTIxM81dNH8+PEoegcujeUS2IdMOWRKUqJ+WuRnHuq7EYs3j0wxkUINZe
RQkZWkzP86emQ59xOZ8W1UaQjg+NVa2KDXmTD4S0dExyL18GK99WKTCahhXi6h7uxXCT8V2rigS3
HqGjo6BFPfkPKFGZ8WMFYAjiD6HFsYVxj6g7vgh7l7C9wAI2WKL1v3TR/vZLBs39iHVRg9pVLYLv
oe0S61uU/FUtzPK4oSj8rdWBe5w+GxRIFjEEAhNlhq3rB2iA8PqXCdKBOh4P9je4RFy1PzssBZ5b
l9nZhcKqiDpjCSaez4aw3+n+HUhiXqity0EpHC1AN+KagT1GQhtJEvvK6H90+3gOCa+tOh9Z1TDw
3mk7k85+7P6JuqS7BDo9QsydIR7gbE3XULMaHiYRw5n0D/0rPt662+0MCi/qKyaRXpW2kJv18Au+
YqDp9bQDgqovtf8pVqhLZPqGhbrdRcjpGnJPHh2CJc7Hmusu4m4t087Q/r0JZ/rfrky+/13x29CQ
9bohuQyp07kljIisGMjC9yga7ZGL1ZlDwE2v5mtaLHpqgDpq2V3tcdoHV9+uRvMgujdhHuCgkFmq
aw14BtGiW1VAkhd8pPkJmmPmRItsuV7V1dOdUKFf/6ZhP02iN5pnruy3Hf51Fo4g1D2n05qdu5l8
r9N+yFWNm+dYO33mW82aCoqb+56ROyZwQRwJtuJn658yjgOIKOPu8hyeMdSTPsc0QlnQsMnGYWvR
jXsIta4X5FPEFTJxQFErE1FU2uUxTfuFaAiZ6C5nQb59RdKdZ17BFd1s/w5+LA780sqfDlJjHeaE
nLbq7mew6LQ/qN9bdTrPdcEFYRsRb6GIGvdExHA7FtMXrZyJWzm8jKAcoPOSavufarvFPUS886np
GDLEDvvMSWN4JBp4uYgxIjT1wo08tF/FZJqnWyFuP5gP5I8F1XWMmi2u+cUMWUN2kNCIgj5JJPzj
TTLkcQ2CZD4/6WpzHISVxQnOB+T5Ky6mHYdJmr0vchgyb5I1MBveQLbp0129x/t4DEBadRQP0rGw
aA+x7bL82Vwj8Bzn2hBf+tqm+5xvC1LYSC91bwcp8VYdE+YHrWOKBir2WJowOF2+EnB6ChhWKSlq
IKuQlH5DX4/QzFslgrBWPii+pvfpRI+UtR01PpnMmfiJcGMsSc177LVnjiEXKAzjcMbweTAULc2J
zBX6Iy8x7C/GAYGLUO3smzk/1wRyhLGpDryHgOH4AAonc0An3vsf1bQwcL3vF6cAHHV+mmY+ijuZ
dG8gFjlH5mCwd6BVhSkqkdvLgERw5/lZbK/v/954gUfcOOjeu4acvsbHwHy5h7XXDdDcfyRUZFj7
kcrDAFab1MAmJMWXVWJi43ZHNidDW4PnTHdvkg80qr8NIJSxMdpOEG0Ft8v7d6G0OqlvS/Zha5Dc
X+clqlQjzsIjaM613JL62w7zKSv4h4QDP4g7+1BsD9zqWADWhzHazJdMUH1no8Dh9aM40qSlelF0
q6I/0ZW0hTaaPPRcoCzUPv4BD+QTghjymTG4CMjP/jYzSMTHnXzlUSPu3QFp1LQCMahomVEc63o+
sPuSEoUUbefc+k1R1RcJTm1TVCAgixx9Ox7xru7Hh/FfqRwaSxsadkhUNMmu6aA1Ilpa993NStI5
73ZArNZRUmQb+6M6qL6Pn6HluCaV8OvCywdDUfKIIEtm0Pu2f4PVefDP/IKtAtgDUYLwFdYZOHOA
cHk9Hk+UofdePMydrIpeUuP8pDioZigw9pc3Xx7ZcjDq8t5YAoDpCRETxVuLUgktvI7j8oXKoAOC
0IaumWYA0tmuoeG+ayZGeuPtjdd9xGR3u3an9Tf0zdWx8L4ptucV/aqgwhusaMgHIHcy+N1Dcl/5
UVV/vNMxVKit8fOZEZenbvOJKxZOlm3s9nn5LlJIyt8ayZl20U7kJplfamTn0+JUYAwMv1HvoDkS
/V0wp3lTMYTKL9R7oruC1jUH4UsxilPmiW/IKzZ9L2uJT6kIaHxHutZxasbXzefSWZdqPAhJSW35
YaNwZbk0LPwoslY5a2LlhYDGyZ/ZelH89wZsl2LQS/37fRpD3A5ns2ItwKwTnvRmDmdKybtXVrdI
lXiJS9FVQNvEox9/envF6ukaZlUHzfADI6ySZp9hIYmk3ZrXLGYJg5CuiFX4R87keH0KBFOF7IaZ
rdhxjm5aLi7n2ScnjCkN9nPI32fUMkt2VOzPHGsuNuLRINswDjusnUXkPqif88YENDNd4sw/1KPg
FIIEp65VG1ZuSsMisvOLWJVPq+BF8Q0SGPqj7VpLUf218qhAc3qVcM3NPKRie4cafU/ID8Z+LWDK
M+PgzYeCT3fSvSkKgHrKP1t5MxQnjTUPyVN5PU1m4gl72BXicmJxdlIc2TSLM7Q81dvjbdBUkLXq
TZH5jlGES6t/GE9Cyj3XcbX17/tsngLDKQNJYqrs/VZdWoigzdle4VjLQ0olljzMe9gLMuIVfQSL
9Cx6zlCVqWraSKTCTYuHRoOLAj9AzVlL1WKgSQfL9sm6RmgQWvpZ2kQi69ePgQiisNXnfm2ku949
AZjxDkpXBLhy6URPlqyts3dot3XcqV52/2ixpPIZbEFQDsvlrNZDHch3l/ky87ibFjZS1rvD4EOw
iIjrVEfkXhsHMa0qAqyh+LUC8jkDtXdoPao3NY5VbS+xCbzW9BxJhMbnYPXS9/Lh+vKNCH7s8xtE
thB7cFzHBL61gCPa29LaAxrSRzpFcCsV3LMyuDhLpo5P4NZPcg3TtFnCOM/zjNhou/aTPzq6SSK6
mZWgZrXCzzMEnQOfcaXeZcFg+A7tjYgZnsv9D5Xjv5843Ib98JdDu4cjqlXepMAe52xo56pJxSgh
dPFjA+UOyBv1X/LarlrJoAwQ8h4iyksbNoXrSLzAC/TEY/O/y/QCUQdGb/UlNu/SuIJ5j+gQ07OR
eqzw6iwUAY3pI1la3mXbuborEKnuqkOnhra7GqNYN+q7mzjERZjZ0x0zB14QQaSJ86zYEvGlAZcS
EiAMvhLS+SlTXFmzsklzhUGENrSETusTQCH3CCZ7BepBf+WqHoy5e7c/3KerWuoaX2I5wSV01+v1
bmJI8HRbTKLCfjRcwwle0kAASLYczw/vemLtwRyQSznOQRyqQ/sgvw7TDJTVO9UgQ8OkxpkBUkRB
5x5moFKZr5712/KYgHD3mOHbLejBHlyWAk4EipfxHXGm/FJ4oJFu8HmvxEmDsi6tAqhRauAd+D0s
z4C6X+N4IZQ3OEgl2Lv/5/gJnt5xOnG0uT4pa2QrtvGZDkbR1rhgh8KOyqt6lkcUZH0DFF87uIEr
GcWH1JdJ+WvDehAs/0jeziHO1jkaywmlJWLnGDWOX2VK0pDCnJzSHjYKZqWlx364iXUHDnXJRVPO
sBANJO+sGtpJD5qQS0Zso5DJkXGkoIpk1ceRc1C1Z3ZdSb5ZVGrvwDqq4qvXBsvBMlh2O2+AJqAT
V7Gj5gKmyf0vOxcxmJjMwses6ZpfDKo5lAI8CyJXaCYhi8TguwHzZKOTgYce60KJVSWHKTRQz73v
UNcw3CIvkgKHwiAEs3moMQ/fxtLf2ZLW8rJB9PFTaQge/Vwl6F1P54GIThQqavq3dFveXlXNFaHQ
WvXEEhh3pjkqNmh9IHiwF0kv2c+mzxtSxhAA5JRE37KLBDRHrLZeKEIks0RaX3xb0zN4nJjwLpwR
6srRM/97jaQT/NSoctMwwh8xUeQ3iytarNErhktQkkbEgl8Nd2per/BoshXTdzYRuqeItzWdWZRM
VAN759YZZ4FB0cKYsy5azsjlJF1x2G3zOuiiK6eDD1fX2cxjMSYMwTnKwP9N4mcGA6qPgu6ToAq/
c1SjGrgnfMM1hRqg+kC4zLAF8wta9nLwylpgmQtlebmQ38jkavsesSVorJ1KWkB4jqZHslYJIS9L
Pn+YTTpAzIEqmq5X0+L5wno0kSYGml2gfSN/fDOnetas+cr0l2ObycXUm54ZuEnD46/FUHQ0f+6f
Oo9bD2Oti0+OOrt2TKenbWvaTkEHvMQfvc+5OUPd4pILJXMiBUM2nniTzLAJ5JmN2FNE3yI2DDWF
hGsPP317Hs6IxmrSqzwlpmsYCiB4OsCLpD36spf8uF29XPypVNctnjMe0aqQy8kZfgSXR6pBfQcs
X2QMci2gN2t4y7XYUGk2qCLDbthVJ6hgnT8XUSdWC5uPtjfw7HAZbV1Ii3vkaXitXzdYSd+QMZsC
OqiFzvDH4YedpmjfInzaaRvbWyEXDQhJ0Tn7icxuK4blyH7OGSkmfr70Lj1b496RxgRZEvq9aGmm
uEOh3RA7wSnspTHddSab5n4ziqLt4DneopgYcQ8nM8qc6uGp++0ox9Uug0y/bLcpXTq9Z2FPIYUU
+EXqmPsb1wapXTE/neSGtr7yzh4DHtZ7uLVgesP7jbyb03DXCZ3JY6zRqOKxf7TtprFbks9rTj7i
2f7qzG+c3U38XsGngCdUPYuaA7UmCgoCtyvrkLn5dVyU0NcFyHsFf5Grn2C2CNdqUEaipQEOiMRd
fUT60o39VVN0SKed9oDxLmeDUN/uI4QqvwPLjwpyGPWoZwP3B87QulsbHdE5vKzE7hOJPeD0iUkp
V+a717XFj2aFy+FhVXhMFcvn1eBmIhm5lgmFGxJm/0l5Y8/vC20DL5uMGEGuXpoknSzJGQBQDzdf
K/vR1Ow6/nm0kkYjUyjUS+tDfBhDFK8e55zaEZXU1gjb20rQ8JGQsVTFxKjBnj4r9TgMk6kZMv4g
l5LIEgMon1cnxmdul8W7WL9D8TXRt55VV9ymLSrqwiJ4ukOAaufJvjJnFjJmE2Zlstjp9MXnqfca
gTTwqxtnA5IinPwRoUYGGNzPwyGVs55m4yIerK9V1QPp+RwfwH8Y3BEdCaW/CMZVYjq6Ncp7uaO5
bEQSZ8MhNY6ot5YaBtbiMXDaGaBGfYULubjF2os9bii5+F2EUmLIi2AGB9LbNvuS8xdwOghevFQ3
aQWxEnwzpx9BkwIrySwr+KDTgwaCmvmVVA1H4LliZ7m7KfIxOLoTM2ATu+SFldlr4jJNz4dXaWzu
aH4gYUz2I49mjiXtBd0uM4RP+XaLI9A9+A1NUjJYhtDo3mQSVD0xFCVzYPSotpDat6n/PPeu8hOB
lfWrbwvVw2qWLgoYnN+muT/GKVPncGkuA1WPO4kth+l1PmAXZB8qa2ech0YRtMDirCFjHYZJ4HKH
Gh9E+OdRA0oQamnvtOA8C5Zb6O1/CNft417UHYl+KrmmBmHLZEIy+fKSEmuHnEQHsgqb5gSMHF7A
Vy1qGOXpGy11EQOafhpCl+eW0PS5mIaMcHGLMDXa1Q3ZLcJP6H4OCulQR/I5ixl0GiNywWe6Ibgr
GCIU+XACjn3AMg3DyNCJ9tmi7TQFOvcjUSOSf/34i9rHVCC2nb0Z6pQZuhFAeY+4YyDTBVh+Sq0N
zCEp9kDt9txO8oKBQND3yLloEHftAUMOvvcW42vqWK0szuVEhraeBF4zmxFjySx0xSnY5gQF9zgh
y0D8VG45QcyufKMLx+oMTpW+dyxGU+RpS/T8KlaadKFtJik/Ey0/PXyLnnPeWluXJnjDWu+sdsoo
0KLVwP2vcR2rP3126D3plNdFjIgpA33/MRbtSkL2D42I2i20B013d5y65eT3Dbq4mOVimbJU7dxl
8G1iYjS3XMJbOt4oO5P3jspE4zZfGxdNTy2UODgk0tD+bjNGQOi0ilqHoruvIszoRuj1aCqygx1e
l1LSiGdrlzEqeqaKg4w5PQQHgsjxHG8/feouGmAD9GslYGjT7rXBM4+r0nQcMPynUyPHq92Rl/yF
bFKLb8WQ0mvmwOpnr+p5XvCdlEuOSiRHyctLvJzn3MFnzSt/koSzSnDvm7VsUxiVo77YKBxTZ0II
MEN1KyWF8wyMDS3RrgL5Kv3pMB7quuETJMy2S+JYOdhMplZD2szjRK26lZO6fXeaNPxmPMm4gGuA
xSBP9Qf6zZlSBSn3r2AZ0ByXdxS4uM4hniC5+pUzeaqiuMe4+WhKGJXMPcl/unnbG55gUmPtAR5t
W7+I6ZcVai5L01bwXDPPFc72sYb5QhlUzvGsuGa1DIxOZKVTKiTjAkzff9DxDPVr/j/MFVWdBjSf
S9swFxf3uHorHwL/ELTmeznZm+PON3vU9x9h+952HYEp/4QVeiFOhrmhKh+qma6eaQQPesfe48TX
0YrtAItk2Q2Cn2QI0r3A0K20nDuMNzmkexcDhmVbd7Zl1d1SBYGgclsulW99LQknfYl38AuBQhkd
IOUC51BDwmjKzJRSZvOEqSqR/jHOj3epuUpnIqtD8jJymX6tdJkCSLWFzeEVEIgSb0+eYBQjWyyq
r96vmn/ToRcTr6PKlFkIcA1hq+kYd4gnkE2h/bbvCuc3s65Y1ldStvoifOtHsvn7Md46Mfg3nX4m
Zvd9R7K8xuEHKwGgtbqDyZRv7Kuk+zPaz0hG+0HBb+TZXY+1WSLWwLof0eyRyJvMbfZfFHWuR0lO
KXR2DPf58rY/NYkN+2B2gOU5JY5iH1eu3h2wThc8ZzgoCxDRx0AP6aXzxr3SqU0jPyCNWgmP9h/x
9dl0ziCTllNq2OslwC6cnPsr4FyIhaZ6BVpcA3Ge/nAwARPYloJKcUDKE4jJpb+2I3uoDi0hPQh2
Scw8F0+98ieDwlOIT+HoRSIV0VPLETHG+QSNWVRTY/MLiFrmrMssqE/5l2CZtDOFDE+gxwM4Spq0
2Y7pkwacCKMWOXRSQKb98j4/fKZ4hLfhWWEntY5ymQipfNB6cfLVLGfxJnP9WhVUV2ldgj7Ak86E
QrXkEqA7GAUG5wP27tNAd1Q4C8WOKbufy4g9xrgL/E56v9IfoltT6hdIvnCQJYzE5+nzsIhH3urp
ZkF88fokvi7/4dpc0pU2spUnyWaaDdTr0njZumkHjO1mB0azxo4j3bHkTxlU8Rl1Qs/U+54inb82
lPsdK+RMvx9Um4lJQRXa/ifNlMqnFOCSgpDMCr8EeHerrxcKsz3Y12xnFtseueFCfGPtCQQEyImN
POVVwkeDzgwg5vBRdaIMQsqwUQ7y9tMCtsjw8+s9tbzf2T2t87pPd0UWnVutiyvQHXby8AbM6L8A
OgoJ649AcNZhJcowC8VpBfC0S4GvW730u8tU2azG+CNO5azT7AfK6J3tMPsOUYhi1fxHI291FSOL
AGY0qPkQuFUvVdIRd/Bfs3XwsSDCDkvadCweQYrxC2rVzEw8lqSS1tTRLLqj16yVTkYaBUfnzVoW
0SfX0K7wu4d8s/DIhR/TZAWA/cekbr0z8CinDwWjxhaeNu90AihjCDhh2RX5Q8V8A+ZM2ul/1dvu
qw5DDCV1WCMBStViMemSZs608jg2orSgLqpZAUD5XarM6Za2SCZHV2JpWZv8LBmq+yQMgTHD8Pw1
49mmwu5DEHAKiZLKTHBnZZe+EP9YZS7g03dDyquhtm+JXEcKHKq68/kw8/Sw40NITsCQObvVhdwH
vaqBRZn8KJeffcYzQvrCODDMYd59PAkW9Elq3er/2XcRFs/O2gOrOdIbXrzCUqZ73cFJx5f2vHFw
USS4Nw94C9E9GBiL/WXKe6D8hF7/ZOR2xxjK8oTYqVFizmMVQZvCeMW+kl0ORzDuz3H2fGSc3jK7
khTUZkqObXnBFJ8gOS7iy/qgmzR5NPI+DGsBrW8aUNLRPcWpep1/Rqi8knJtbFCoCPkEuukNb+1C
RbnegEyo4LV0zxYxAvdSroE7jieop0e6FHKOIoJ47nyuOYHrM9UUXAjzVlSFtiPrJyyWzY0u+aoV
ewhohXTTBgHrcskt3WBOn1Ra0jKyqyQxdAgJKqUmDseg/A7oaD80Lti5oLID+h8dKfk9JddnrZIY
FN+B7h6p1LkqkmBio2ndQY5JMZ31lhN19AYJt0izQRy/TNP10tQDnJYUvEn2olYF0ydVdqdJ9bH9
NCJqFFSshpFCUGgRzqY6Nyql41BgITBwZZuO7Nz+U80EBVHlVzMW4L1+ZKFkjcNR5uUG82dAtbNI
4AC8kCh7kDlYZFse9Ka/PlkVojnM3XNf84vYZ4w3wEgJWxbBofY52dltaMaj9PoTZkQ2gFaTvfew
FixtPL+Ncaje9j7FxNFXO9nO1s6v+9Ea52nfCegH66j/3T/8P1+WtgdjUArrorT0TZkwTDRK4XaR
5Q5cYHqIuJt0Rkl52/CFfp1OELCkVkEh+XZJxuHYXSVbUti1ajZSGUqCpSaPh3Ocw8qBdTVeHfvJ
fy6UqORDsGaZlZJml7wyEoL8O2OOzbda+eQZjR7vvem5Y83aIGR+K++X243O255nScIp3KeDr2Ag
wX7TLFT2TRxyK+QIy/L9dRZJML7edL0N2VnAmEBNdvSRG7+9Pan3BautlyF/Q3sqqaXza01xA+EE
zKL2P0XFISIk6sl/VBM1vFRaxL2yJGsQB+SWYgUhL1OtICrgfspKsGIj/kY8c4pvUwAPwfanYYNW
uJNxluvyzfoWrpA5u4dkDC0P8jfzVzl6YsWL/zp/mbUs05T/BlcQ2vrJnLMJ8/VBI8nDsU3zcf2V
y2Ajyt9G5I7YjI30ZxyCtAfk2TOtOqBoSIPIGgxOV6SRpCnlMuxPZ6PRfwDOTMjcZfrE01su0WdM
ZxviYKO8t7FfpDXBHIzuCvHjHJMOCybPOn9NmnhxkS11UDlixOaPJoXupPwCWSWHZL+d4k04eKfF
yZLD65q0pygxZl1pIYSRvXhYaCx2etL3ZndLBPFWNi2hBj1CdBdtF7wetUB+RPOoHIo/yFQUGrRM
Yun014NyLu+k3wLE+3CC6hn89MVa90ZJFER2J0nHDh2S3jUu8sR+3oTHgTlJmqbukSzuQnR48otj
Z09AjIlbeX91sKv0q7OymN4zV6ZuBzmsG2pRLGrAVcflT8JcmqsG1f5Gsj0KJ8OIFQemo8QxatpX
YCQntjZCMYTHDAFzCKJRij2xa/xPCusXZNWno2tmzoExAbgCrRWQKpAexcf9oCn5R7zoErDNGjS+
SwNxc8Q9kZHJRTAgIoBrAcvCB6JrNsTQHa3VsrG2RooWhST84Og/x6yArUv2pA8aNfxkXyoGTK4F
2DElJQTj58dey1um2IF6sjgQplR6ktiKRPILMqojNWM6T3mj8hu5xffmMhwthpZqXNG6FaaEn1T/
wzlSvmqTUeQNRgxfSDdghWVSOtPlZOdkjEzjq3O1pwr4pRBkXPG7+rWCUTYYLmp4Fzog4MVHRZ9m
XgzDrpt9SM6JoHO58fpG0PzE80q/H5ggsf8jPWIQtZMh8l6q3HXgVvVAfAN2YN4ybjaj3k9uaqkP
042xoduoK68gNIHpU7FRIzIn5diZBlSKNd8HbEF9RFNRgElK44Xx0XPTQpTto6fgM4xuETyHRl6Q
vfq4zh5GFwS3jkgEIGzipATCG5N6UlpEZWiq+/3VAGhoXYG8LqjF4PuIen1r84DrH9JuwObDH50d
+F+qeJXkSM2maHYmiDVGFOAAY2ma+zRTkPysoPsG5Xn1Hw3TiiDyc+yL1rXAY0cQchQk58xXONGF
CtqC7U2BO7GGfSHD7shz/A/eK2O/6RdH63ycfPTHy0MTcuCar47YqfPQZe/WK1fNTfJ+aqnlKKA1
4Zh/3cXGIvAHCBswl+Uz2tQyYdl9l8dpbLHdi50k/blyLjZhsokzBAWnVXK3x0ws6s2w/SSqW6bh
FLtWyrCYCyPwDb1JHG7DZGnJ7VWZoSYZK+PIw3larQo9Zw0O6akKqXy0wf4AKDisIvJEEyTR+VcK
CXfHqY4zrcx2UgUTmkeWUhPgcVIRDo3IHt3s4Z719thrvFc5LPWj5nvBybau7FbwY68sMstSs6O0
d/cYJCRkbjeImWD1cDn1V3WJtelD/rqTBWfeVnx9QOcT9IPVHXgf9fu7UreBLPOLA+gVnNH+jUUd
YYmqDYly+mvkjY/VXpxUI+Byth5nOfjvak3aW9sQmWmfxZ8BzEwq+eYtarSrJfL9KAoesAIWw6jW
/AYZIb6da3fqQg6DLqJfxs/TsT9lg1o3zM4YEtIvUie8IqsQdG/hb7cFUtDaqUyoq8w32BMI2Q3H
Jz46rNlgbnECqHsx9EpIOaBH61cW1v3OlnPFVw3Qn522EgPtbOtX+YF9ihhX1djLFOSpopyb563m
gJTDYwkRfhv6D5/YonWtvIifQ0kBlS+7YSwqnWYPJCNpPs/2ec1Pq8UgRFd7cVmhgjGsVkKDXvxr
hx0UoMG+q90EDbh18UgCJEK2LZNY+1OBexxf54xqwmSYfskGiUEzuEZheIpYlhcC92hrD+8/Xxft
vXCfjNa7ocJLWz+AdQnMrGQ8fEye1IWC7DPnTRKbG90k8qmfL02MqjQOtVJ+0HkUztDeT6CcnrnJ
G2IG4ecMB2BiZZkWgQ034XN9R1GTslC2Z78bEklamkolaBgrYhJry/IumZzItLGyrATCW2AHQ2uQ
JGGNQjK8oTys9/tB6Il+GuX/wPsS5Qny4YoCAE8joYjEAwy3RArMpgq2qDzOXnDDfhW5azaSWke4
c9NZcN+Tuv3KtQfhiTJzvirLXIXHXBBHDrNlpqBfS9g0yfuKsAKw7HvQaPhoNox+3DM1TfxBZmoG
xir+aeUVCtqUZP4r/7VKjnU+bdza2l3Mlo7+ROyWZBx0oDd1ie7aBSrNs66wWtIvfG34YPHUBJbH
efb/7qjx74nWsVC3+e9NT409cjra3YyCWPrNDnbICPJLGmaclahPbaeMOHsDcmMAG0EdFASgtdP1
D3ze6CQyo1t4rm3tANuVJxsphE5Twqr6ZuUGd3/oOC0JKqGvZebcbVQJlNhtyQ7b9H3WJvY116VT
N2PP2EHL+7JpbDlHmUPjlcH6a3Ybkjn7XfViVmKlPDW4MP9OpciOsIZ5VGekB3e57U7wozRcOAVR
e5WoWgmlLKwhPrBXf38EQRCqX8OuASopE7+DJHl7Eh1Is6qZq1p3TFO1sssnhsy6cj2xBftv+JIJ
QWlZqzyRJ+VGviO/QsThvwToI0ftsie/loFYZtt2pnXadaX6KQfbZ8T3c/HlcxwRlxmuWRZq5+U8
CWMueX9FRPS/imycxfgxUvRzHEhOFUDBEORSqI8JQIQ3r/7OCPRWWj1EcOdNn693XJycm0GgJGIo
jGjfEoO3TPIt40CKN1XhBYM0kGPc1isq2wxjdyZa1plBpAsMjnAVkTwJ/VzNxc4RoY+U52sgbvFI
ExwKZPXw63nq6xtzQBEKiKKp/dnJJQP7XDxtdvyMpG22EI8qKW5jTphyDsEgGSLAeCVV7GbjoYAh
AvlCKgJ/TSWNI/ewX8gu/x/aNRS6BjWTJO9DD1FwAFDlg/uZrxpPdw6Un5UNFPF37WDQX+Yqi1R7
gIJJ5ujg3qC7G6SmZH7xUihQCzMmhxWk+QQWw4Ci1eSKiWo8fP9DF/SVWojGn5cS4c6t+Vo+tWhf
YRmBxtoDDhXonnjmy6dHPtSBa3rlk0NqN4uSm89vj7W9VFHxkl8MoGHOPOxth2KEbK6CIc7g+BOE
u5uQBzM5djWHzNgGlonFomGgxlIVMAdvsMbIUdw0Im0KgstsMyS2ku6Spv/+i9ANO8qk+BKJSwtc
h2cr3/yKPW1sr7XvUB3Rt7JnvqSNlXo0GvXP/lt4PeAzu+thFFQqI6kyUiccTktmipVkKE1h4r97
YPl+DRzG+pK9xlX/hPc5VaRqdOKc1cj+4iIeCww7XFhLDsrCfR5WkoXrDtFpq6JxrXfoJVEF4GLF
xHCO3ctOnK8KbUGMhx4eb6IhLG0jtk0uyc6QJpe24fD77dh/5GTI4sb1b60d7AHDxVT+S6IiW0b0
y+Q9try0RgpRQk3aXvibwtEcub1xGZUXwceHxbqI5Un55LyMbmHjbkjNlGaX/HzHxLpaqpxTcGq1
n7ltsesZ+j6jwYyciNMKho8qM1fyq12YLSgqGJagrg3lDdTpcSdnC1w4UGBrssxkTWsshDQLzIXu
ATzwF8J5kT5/XkFMO+jRm/EMjxPB303qx6XIgYFfkAvaT2wmoSkZL1cpY9OhiDWhsZOHXfMtWKEw
3j/R1CGfPLecxVFuttboRbIkxKP7cQCDyN6JL2lVn/4ADXsdwK0xhZS/PqUAv0f4+tc/2oe7UoQA
XiMwOBPtBtNKAUqjefFBbjFJSa1jrrW+0XPMHY9rYmm40nzw/BodvaGugYKNio9IfFbPsMVkTMSs
LxAKqb8pxeR3HuUNtsBlMh7iff9aaN0Bls3ObYjKANmYewp3YzA5RJ1wU4cn5IuU4btmJ08obU5n
dMKAgf7bsHUJ65TSK+vnIRSGm3dadfcZ+O9XVjjAhViagNgBhDHHuH4ebkUx8Ep2w/waZBm3D5p0
EqbeY2mPqQQejWPVG272NYTUjsMk84xzpHRsXXTbJYUAKPcyBczAxD/lDxhfZViPamuw+ME7GM0X
gPkPNi+njbZ+hc/lCudC6cK0xd5YkG/KnRMEJ9ip0SyFBMaFYcjglB4c8tgNImTAESvwc+NJXSSq
mijy5aG2FohZMbcFJHSQXvxlOX0hXgQniqGL6Fi6RqorwYs6rey8OCmCcXh4Uep71526qGFF52a+
/MRxkga9FusyTe1POPAtX+gvCuMmleXurhKahRsWRrl33aWsWWi8oGXUk51f6kFu5a0XenoWIv86
B4vpHmUL+8QXFI+wqRY3vB2o/7F325cng7WTPHsiEaZcGPPS7SKWTu//HdAA/qP12JCye2z7+WW0
UhERf3/s2ygaJJjUBqr0qkUyzRzwjJsbr8hhpj+q5lYP0ppjpl5GMsMhZCQXltA00EzT24vrl9l8
NP3zB4YxUatX12hvVZ+LRsgP7P2Ks3T1woiSm5J8aAQaNFTJiSUII0Bjw3+r6cRSLjAM27XkPqUQ
o1ERBITuOh5R4Nz62o8tBkvxgA/uwG5TADIOTycl3jcI9C+6Tpu8oc4ZETKjPW7DmuWhf71tGEJ6
yTdqTdHpN19bfXNW8Q33U0yEA1aQS1QMnKl2CgFcHvclKWijI8hFVmLJzp3IcNiX4JRQQtDCbUPM
O3EsuM0UJaOVtRI1fH5lqMxZINWt31nXcsiMDfiKcqpR5kjSaE6h2iKqFg8vbNZnkAChjX/dWjg3
L3cHiqRbODD8705Kug/8n0bNLem57Z1po0t/QbdX8ejFTyvSf+ZkRBamg70qUV4hsfM1umC9Ffcy
dSDRY4DwyLHWQFs0DXpBYwpIMp++kjkgdC5ePfQHs37xPNzbGn5cXGzG9Vtpz95+5Pp5aXuDxMRp
S9hwtmPzwX0pKI2nSJQ2enacV2suI9gysJdIM43mNHjfecQeiZIZEB/NfQUYJEFQqOCdR2aaxFXO
NUeh+iSccViehHxJSfzDBjpWIKykmoUVZaMGgVGywiGaodvoBBRyM2sSs3NZ8QcsaNzfC6PuuNxB
Uz+kyjV5fJCZqnYoclVg7TlJe1EID1LLOqEh2c6CN0xER3VFibVqH6GA3XlccClDyr3D+Z8bsRVr
JxyHRDGVUm6Z38mYWaZqE5bI43Uct3uYzmMZWDFRgfSK+75OfIaP5x4bhyvoASzT940jWccFHMQk
pUG8861svE5hKz6zTGDBzj2Xpf8x7nPoqpKyjCn1xGsqLDZjEqMvrkXyXgTgy1MoIchE8MwfEqv3
zXL55bDsVFs6WVDu4+cQUw8Kknc553vaNAj4YduuXZfILTzBpChrlP/BgvErYsgsDNuVAKkH98ou
HVY1RI61ptvJWsMMSg8qnNcL81y5oJLEEa60y71w9BkTVQ9AKQIDdPjpNyLq46hpe+fB4UrxYf35
QU/nHBXNwAXz3Lgie9Ic1zcpqKoXwLOtAuX3Uwy9X1SxX9NwY2F91FfOL4IjenFO+D0JuCF11HN2
QPeVz+t/uodC/HaLhh3iAkoCz3PqeTRip/aI3A8kNnYhrb6NFcChKc/cSmcTb0pmIA1q2B/3jxta
5ZMb4PdOfw8O9whGaDbvWm5NZCr4xIXdQI55o2DPdOxA7MKTS2TcRdVzhqNHD6hmQd4KZ29lzc23
EH8UKk6zcke7XXIngKOaYnLXyHStuKDt5j2tF686AGZGkZEYR5szMH4Oc80dZtknPjVZ6eTr05yX
j8B0jQJzkFNX92RovYKYc7SY9PNiYLNVwx+6T1G/56enbiyxMLq2XNqO24EG5Z9o89hZuR5WSx3u
KPcJhPnFn72MBhnEDDuLT3ynirFATqBNa2NZaNfV54BO+A/6V/9Zm5CIgm62IvRBqt41iV5a+S87
TE05Pb5ECa+E23MP4cIe6oY9+IwxYDdFUr6JySkAqjv5yyGZJoVa+BZyICMuokDlGt140UHW67JH
BRCtd2vYmT/YJH6kR7AS9Z3WG/z0VA3wVXD+JPj8JLybwg2B/aL7O0mYAUYWjqD+uGwLK5uLouYg
8Fi1+zJX1ktXKKW1kNlxxWd139S/as354KLHYpk5uXwlCLsAqqvssxGLUOdtpG0h8yB4rx+Shl3j
90AqQ5zqwIGF9wwHMXya3nzAtH3E6hHqVKVbrqXCTWbLkQrvYJP6ZQnyqBiM72pOoZA0d7JR46f8
ZMuUXnlsfhOKbuEyoJnGgBGaZB5yLk/KC0LeO7ZrjAs3C3S8dU1h3u5ByvrbiOcuf+VCeGLAJab8
KFBsYLaJElHUd6ytUYn74zcoDxeI0/ORBRes2h7dhb9gBMkPlAa/wZl80lDxgvvftKh7/umocQDB
uuIVxFQQiIa8DHQ/2diX6pFeFw0s/3/KgyDmpnu3G6ZxpzyK7wjRntl4onddUchvBnrqa6cinrWt
oCq9ySxHMfsE9GbnuJjNCMfTuePZTGdELYM74JN5kpHI87Zq4bscAVL+jQCVVNZ7Ro5Z1NyBC86Q
pwZBpVJULsFA4vMLla77/yGvv9/OMHT270OX1eOKcT01WAB6sCoB54Mk0J9sOJfLlxDhfgFM+UX9
dBC1Qog5OD5KvkVBY4P1ifBetcFWM/S2r9c/O5GmRoRHlUd0GJEvPJeAHFnwVFmLk5dfCCPzQOM3
KnvZ6jDTtYnrGUHR4P5XmdHVLot6XMOjnKlZD0FKGeR0xX0QqaHrNHnftFKedOl/UvAJ58QH0gNe
r/tI9A88Wlx6OBZFslpmRgtoktFQjQU6a9y3gPDjfl+Tz/d8BgCZE+DC/1WnBes4dBdNu5HIAMyU
pQPLK/3JFWXlQTQ2JypCLUErshDFeBPC2zQpJ2otCbC+0YWQTKucQvIiivOQuyTi4uZ6bxHCuwxv
CQ0baAelu8qfFJtOrEcq7xrYVRETfEpHE1Nf7aO0Xk/JkivFgMrQ8MjJ0HJ/3nk4vIrNBO/tWZOd
Ymd0/B7EWsyBNzdgTxX4KjKBuE08RZd4JxZZYu0SUWeWOm6IW+OmfpWmleYk/QCYUYOUlZWVpUKV
l0mdoOSQ5TX+uAKL3X0lHhaDdIn60ZKiHMdrryxDAv5rH1iOIMazMS9bAOV9l+V3lBxSoh3dV4xT
B8gz2/efSjXYl2ePQ78sNvRjnZAr94W0qFSfcmYi64yAsTKe1uAwkV5yUl9N5moRBQvjruIxrh8Q
xTiPuFZ+jUN++OBKFH3tsx8jiFdFfv7K+J8GJkJpB3/kN+SA7hkBWyY07zp9PyLpCof2nbNIxE6F
UyAxFbYin7O9W1Ow8AjI0xBu2Ua8WSLRAXhg+4zIerZq6XkFlNr3ugO8t4jnOlxTeSupfGD8tRnG
t4FZHcqGTgjwGBa5+Y6m1pfwu25JFcYT/MmGJObHFvl5LQ15DbQ2XE5gpv66XkTWzHyBfnFd21qV
Slvi+CPWJyq5jFiGobu88ttgN5UEbfGpu+NWCaYlfI33O96BTiRybYRlxfTdU4rCRtgxN4VFn+gF
It2G0W2Et2toufb0CIGa5BCAQfhLBJyfXfzHmTSusxjrfEtrc3O19ihX/0tKih1U/krathIn5lUs
rq7UE76bgg1hndeHxvNfv8ClN5u3bbr4PgJNloklWfRfzoCPeF3DNEWepKWDkrfKpl2y36P/aCsf
vBGkywt94yvtC/D5LHuNdYuBsoLXIgSh0XeMB/Enmvyn6iJ1rmj5Pk3JoBLP+Rok40yh5NKRqNoa
ySD6r3r7C/ZFGhhnrX5H6G/hbTkFPNpUgyytd1PSPYQ4oGrl6aZapsRUzSok5WMSJQVLBLrN2TM9
i97B05OVN2BMmE57SyYTn8tAyzUzhcorx6jk+4RKlNvZJvwgl7tzZE5vOxhHFjBQ+qhqlR/fWFUI
MPZ72GCI6Fa8rbkTMFcG//UY99OoYr8bnePNDIQQOvhA+ShtBWu2KFp/q9DE01HUlDwxtDUGDJoU
7qmzZSSlIJswBjpRPOigaRDGcfaTdBwXW67gAt573Eu/5eyMgR0rd/xSD3/3FYgFTf7ac6N0ZZKN
619ZrkTd4ddzqNTlQQuaha4946DOg/PpJLe3H/R27r6RpRzX8+cc3T80NlMx1ZLeD2JRYJUuOp+K
w1AYXO9isgZA1i2jzUGDsllydOIfmtWkdRr6uBP4AjjNknrCoX1rgQRrpUY3BLcUa34LZyc+kCYs
YlX833ZVoB0f4vBmPLV3hgw4Yr6KB0+MVu9ETGYarFjKQF8P6Td1QgDZJajfXu/hPEqYPs89FDxr
J55dMb3oafY1nOtTct2nXe8622ExBH3scNQPh8kpLYEJwGmwlJGWW5paX4Rs+lMtlxGzGTHcisB6
8EvXZv77O4ZohJEUhRanw5oRBsO+uDN1VfIg2hLPCj+9agiQpSGQi22y6/uvQdtDcwuAqefIkW5v
VJmLREIN+UXJXjpWYYFK16MRC4k9LkDwkF4mLy3K0rT7B30De79SrfLry6lH3i39Z3vEZYuPmc2j
tsQHf/TsNmOyD6pbt/Vnc2Q0jdCrpz/1iLtsj5BI/z8E/2T56la6hjPWM5cCsfXoDOjnQuR7vyBY
+rDJk68p3gq5Jg0kR0dpTT/zBuyO0r8r4rBnBcdpd7GPDmCS7rL4KwKtoBGsRccDETVzePNGBjGC
ULW5AJ++RaW4v/nTxXHEus1DSzR5yvtyH0j9IpNpDDm8sB5yvdLwA3dqWs5PsXckjE5m/vWT5hQK
7a3V3XFORrOCvPv9wT+OpQp1fawqFKvKkXgc5XRD/OFnQC7dunpHoxYt0Lmljxi4k8DpYSpZtoCA
/ol3V5Q7YZS03Hz7Q9tVf0VQNTQwTBonb3bU44UWWyfu9f1Cg2dlMiQztdfoskWb+iFK+v/8GT1d
L4q6cwoWdum9MDa4Y6NufVOa3C75/kZicNWjF4Ep68N5yr1vUNrePO3f90sjSqPbltezYdx+VOvN
onhqbYzATHTM317anE8DGI6wx/HBjq8BGpt4NVMaf+mWMrINN9zagC9AT2TC9VO3hQNoYW0U+7yQ
Bcd8/QQRsAJld7DTyJxmYpzHq43hu9MY8/upu8s++fvUmC4HbxvVlOhNF/t2yMhMVK3ZpKGFSBzd
1WRbWfbmkoqf0MDE0FYDK5yby2a1+Kzv8//E/2fZTpKPT663H9/GWa5+q520grVsjMbeweqepmd1
Lx3AvRh8Oz725xh38UbVa8GRAjn8FB7n/TCa1T8+mFnLbQeEd/wYC2JOBmh1FEHPVbKRiI+bVH14
P9rqQaKdCFXzqJGWe40b5hRBsFE98Hl3oEu51arjsuvGEjEnoH3/5ENqO2K7gZtV+Lkq/aV1xO/h
7DIROEthR1+A+iX29BJQB3dcpC/2pxSHVhhM9w6uyDitrKbQEWW0mskx3Lhed4JXjwcDsg/aUcVo
UsSjXmD+XtlZms7FbCmMjTvVnsqf6ltTc+s/giuuudBTKN/ZDqf8DihGHo71dQmjyMno5M3KkeSh
kSZAEhuGBuRsHJJZWsmeLFuS5EwlzI7ZXLDfwTehqwPYspjpiJFB0oGJZfhvHccxRF82s5DJfiWF
h97QANQALtUitCEdE31HVEmltAGga4WVicF7FQocGVLaW5ydWuA5dteS1k/HV0HHdN2aRxFxTeyQ
PFK+zr4pRLs8CthNTS8LTGSKWRLaVCxejaolhdW2IqvDz201y/CF1rvu0vSEeS/+ZV99G3iDrS51
0WG4pp3VZUhHKXbXyOoep15PPi1R9GY9tpq742uwu+pOf4T/aA6QjKwuQBceh12Yfe9qaHzeEtgN
xmKIbsqc6pLQRKEE3xrjBzg+rq4H9ZXXoMpXmFLuYUEprJgNj0f0DJkhWWdT9z5fIyNsgWEl2MeL
kS2naPtpMgxez7wG/7sbuL4+is9NdQGSTNqvQ3H25gME/b+uyl31poJ3YfqKMO3RIsXUjsvodAx7
2/LlPkzTFefi21DZ2BKZ2RjlgPNhuWS743DaUTTnn1n0uxasXePJf6hIN2atb2f/5XiY5K1ODx3x
OsINWIaRAAOock+rCqQLea1eMoFys/lY/9iDBUKyrEq/MkTWMaAHTYTohzOIxF6FhpTUT7nPdRLA
RLAHGB/JcEcJCU3d93MEwipjHJruZYADxSl7KJzvYBCW0GnocEdQ6fvImZyqOLZIH7VsYW5nB1A4
Kww1MIz1PlVLRQ0JCxIDKPIHCEq9uBM4Tsknh56bLM/Z9PAFBZPqFgJPMj7m/y3eRTq4xKpLtWyq
hrKDumlqtYa7N35UjgzwvoiQPdGwNCTNVibV4h43RfXF2X/asrmA0gw7VlrVksJVKbUsrq+wbveU
T57LNYkBP4ddRvhlNp8SAmtZZGy6xyMtnFrnya0PWwL1i82dLeIE4Rdp2xYUKNO00xjnCcb4IH0j
IF+jXa21/0PhJkrNTsIinsInGFK5V1cBm2/STPwZ7381ZfNNFUDGkkhP90gct/utSQ4f7CGwRRdF
5uL6ototBUcfuOcQium0JNRV+S9j/L8Cd0ZxPKkG1c8kkqhZ/QnJvRhZZutyHQiHaTrTlfiAMe+B
2N9R58ApOXKV1lqFbp3wg3LVS53k2c9aAhmoucCHSpLPDbY4yPZ6xLxKDSOZ9jvwH0pv0bwa3LYw
jeWfMFUhHl5tc614pPqP3VCdmfKH0sAD2+v0sRly+iWf1YgbabX028LoPzGS7PGvEpOaUay3wCha
cqYeGJKVe9/SZBRQbij4vRqVrOPs0sTT5GZnG5sFMXlDQkCqlHg+5QnhoufVqmzfZqWfkvl9CRY2
Hwg7wt3SZbLiFjqmXl/6YaYwBz43mk4WHuQpS8sf0PbfPmoJrKKtqnEiz/VHq5yxfKyRsjIU8DmZ
zzzdD7xnxTo2U8LqX2NR2Q/gOV7F0kCZIMRJCPmUsuZsucAH2DrJxgzq07wFQ3hJw67nCPuuJPzM
v11SGHxSL2bRP2R8BV3avXRiOJBm0LnR0kBVpca/dv0cQwTOMcXvPWfCpb7GaVXAB5kSDZOrzDR8
Vt483fcimNwMdGcysNK/4Q96u1WuMbx3C2lvvOmOmVRgVUu8J1Y4n0avW1Pn3krhMr1LbzSNIbQm
v65MYwbbHRO4NIm+gJoKz1AsfMZuPfVFIx//WTBuF6jNVxOyRaHLpKnwOri50AY/xWjd2bMf/NVc
O6aEz5XF/1Jt/1pUlGWqRwgFsYYTAD+4ZYOsitdcfRI8TxF8t1+6JrNKkqU1GjQDnCcvxrnPjeIu
0cHoueOJ0v3eSNOPO1dw38yPRfbo9kNRbTrzp7uHe8fXoytD95+xpej+xKyFGIQsFu7xnpc1Q6cz
667hjqOIE+0SbLBCODufk5j3mFr5b/mtxgRQI4r7z25qmyYcPCAfCkoq3173h/Y/nBgnTroyf7kd
dgaXvj1RAmQdJPvsvGIWG/z+jcq++B9HyvEjIxoHbHKAJxz/lqdRtI5Xl9BGzCczDW4HlIQNTN34
CNT6pHCLKttrl2+ErjnAiXSI+w/kJBO8Znyrpna9EDyEWRfXlgRwtRqAMnQFwzBaNDnpc/bOkzp/
WxjRmH7+aBsUk+lBlhGzbGdo+Kj/yagsSM8qLFHXlQCgAeWEni1ZnQxiBNgklGx+dy9bWhUm89dk
P6ZX2yOqSxzjd80uzXslrKiXFc2XqixPnIfa/4/4dHCaJq7nzhRXkWb1KEczn5zVjGmSHgdcFpVl
+BCxyV/NiZ5EeWL7/3WbxhsU4KI31vC0RimupqYprJveMPjZ37m/oL5fnEfJ504qcpSTutbU0/Qx
4HbH9yd6B4A2RhvqEgLy27cXuv69toiVA0+DsMwLS37qpjEts9N6G+dh/JkTYrNdWeG1AXzPUMkU
48loobnHb3Tp8ceK/D/aJmZ2tpJAA2yHiG8Nfpx+IhB+1dgJoyA43Knj/ByD+rY874LmfYM8hx7h
AR9T/IzFYhBd+DTEZGdg76Nl7y0TvXrXyV+P5RSonRSVzmUhfjAx0MppajCStDKKwaRqseV+kw66
INfpYt6NLA56N1PNx3TyiRtN0GZ5iYR4Jt48s0JiHMwI3pwZUSjtoVSWmLlKI85F9JOPPzjOumRp
P/VtAYrKyow3mhZHK7h3JyqO30vTiSljNyLKLdludYCH41tlErnq8Gku9cFukoPJvHsilXXtlieu
pnfqV5VgoqAY/YyWQCisDTln5xWheeBZLPuONiytQtpJJSdw+YNZBCTup5NcA3xFfsqwNvwp1NQf
hFB1bidRk1z0B4heIhTSR4VCNXtRYiNVfkpgWZ18EkvJDb8u04N2mLv8VfhKflyS73ZbwtT6bSEL
DQXXHvGAVyHQ6MuQCuBLNCl8nMhQZjHRNBrAz/MV/tm1nraZaB9ly+bdf8ZFUTzkLbucP93d9fSw
JrJEOjUyVoFI++5D259fWBlnMmYtPR2DZ7ONYGPzO2vHooPtMHonToILOs87t6WIm9+2Rih5WltH
9Y937KCb90vgbzCiX9OKR8l+WwGTqFNXZ70gfEicVf9RCVZxsmy5w9XViJ5c3uwFVwDummjhp3N5
vYzjAxXdBK7WtbywDfb3adGZCmHAZhy/Wy2PTpdTzGav1hCfZyFNqjY5qEBgPVTzDB9+d6LP3zRs
/4YWiI0v9fBmniDEfsWaYk3iKQ/paKehC5DO1n1dXrSxb69Ko/tjZj+ql+p2jDtIxGnWepKYNPDT
8p0H9YgF4HGj9Nl2JNinA7SgmdZb5fa4zKQpFlFTQmu03mWh0CG9em/wJs1u6gKSNbPQ12b6R3Ov
ITLce0MbCpap/+G9SfsShojA3JCMQDffp16KA60hJVcZjufBq837EnlHlQMpZWGAFAEB3oLOLc7i
9b9bBPypZrZF2ndQtmmtBEsURlUi8SaXHzy+PkLkRzapvxd/unL8peuw8UPOw1ps4SDxNrejSLrR
vyiYqjoo9zGITQAD4JlsRahwvVAGcroWn9ogfsOU1jILimw7+uNF3MdWoZ/MTPOEkYBg0/BZKcdp
tzxIYCTkEarJeEnTE0nUOKxC3I4PYBLkoScMwJwfAttSmOeMtvJ0sEfH9zipOKGbN/YXEmRvphoo
ZfxX4g68570QEqpye6DW9CYnNwiiyXX+kj0nPO3YCJgiFxtlPD1kfTekbVjjtDc400G87Hc5TWEk
l0jp2Wn35LKT3X4yfbb3/dDc7qSU8CtX+r5wAiUVEqooC9UzeOsGYVdQiigNt0vqsOZ4HDHn+T1L
YIAiZ3LfPu523vnUxu/pGpyDkXQUexqcj63hSyXKFdIhuaBWg638wcsRu63a4fkU89JPDVKPRGEC
bOVuNNkFTIpgAh6rGDA05jlvZ7AXO+JnFIgpbRcRLJkdiYJHLbMDrq9/qXF6R9lk1Of7zGi0kpjn
uqMFW8u9NsMCGzu5foEilZvxivKGNpg/taTOibH1jsXqPkIL6mtajT8+AyhgSRYSPdmPEzgQLihM
GgSZgTM6cB+jIwIrduUZpiblPUxV87hFLjgq23udqM+XVq4NPrxSXAOC3aGurYtZl20ZtrMMzgVZ
+RlnJUE1uqtbS9i4JJflYCK/STRnHac2MXlFZGBGCftX17PfHm+g/zwgvXht4bdcYIGH1S3Ukca1
dT6DeZ4HUPoGjV8d3uXL6plV01UL3CKxgXrIQXJG/mjhiPztyewJKcQIEzkdIZjmCKJ8L/RgSChd
bNytowtoK4gS+DJUQPYMmdle8wQG14/8n2GAA53y4aEMtPjGMiBQ7TCcUkCDvtQa9o3Op1IO7GNw
l7RJATnT3Z48tEUTFtXageJlyoMqxyh7P0jBzr8eeisOlXIJm+xUIVAi9srogsAteoPfObBHMGKE
T6ZkM571sysb328qDY/gbpCrtD0EIubmqwhAkyu1HvsaH5WbTKktmSuHw6VHEalb0SmPoYGey6OT
e3wbIphTpriXQxz4IWQaWYiZHAYZxwpCEuXuiEIXUehjTVtpJJX7dBTwClqrvjZ65+T/OyyDDNZc
tWd189he9AqWMfwWzQT7BhDV7GQsb76sVn9nEsOgFUOsY9WO3sU+iYkelKzYWZ7O/VeKSYojMPSj
QLvk56aRN73Fj0bZCw+VQuFm3jvsGDdLSAxh7veB0nzR0APrpL5BsEg5z+H0Ju0Om/swXbeMybyf
Rxu7h1j3p0Av2rRRjGvcfSH8GmI63Wx9askqscb6L0+8QGUaUmPIf0M9Hu9fvOsPd6dHqJeTWRWp
QlPdOcWxegaBazzUJV+a10TUsoCtHhhQj56nwz6UkacKiDPuk84AAg5t07P89yz+6H+VgHCgHv7r
mKRsBlBM4eQx0tsErzEIFuaZ3v4ivV+pjJGaZej57qXHZ/1CkOo0gZC9XFkJATM6ikGi0Dxwccl8
zBPTXlQxftvSF4Oog0fz9tDa7roW3x6vtLIVomV5KRxCb9RkvEwd6hIeO7l9fIxZrlMapaOStfiN
q+ezVSfNiDB/9+Jcwg2BYPE4IddmzqjE+mbSZFkKs0gQ+SPqkGJu7EKin2tOiMMxHgWOLZ3guy4k
oVFKcuef9m7i30Woi37Hu9HnAT8GFpuuL+5T7EAxo7J1rQouwAVhpu3flIsBL7GWTfAzMaPnNv2A
l+zoUfi5njl8BE5i7hz6gw9hASIz6JL5m+4oPkyeoDut8AIfAn4IAwx1ePU8lsOmytO833rCnGJk
z9/SCfrVHeRhXAORr5P+eN5cKBVPBpemhO+jYvIBDM3mWPFBWOfDs3PijgZb/bRae5yBmWwg8rQS
K7MrC86rQYXQv6ZrnxhbTiXZB1K5A32+/NPTWjervRl1dR/p03GACShXV1FYxDc6qPK0GGI4Yryt
gdxDus7ORTb8tgkGZvJEbGA7cN4MPjeL4VOoUHktsi500SlNvA2mLnpiIWxfhb5ppjVHtUZA5PzI
vmDWbyofKvBfM/+HHJETh+YUQV16sE4G4TIt7BM1AJewfsafStoFW3J60ZMJri9McsIw6kDUatlW
B/liHvzEcmCwxUhLnLaV1GwYR1PhW2bhn0hGb/ByPnsUCA9odsufFlL68p8gHO1Okc22T6FX2nKH
RjPsGbzmcfalesEYtwSa0Lilhe1+tRGcib2TEmH1U8Pf61s0QrUrdI/tmw8gRJ0RszDUxh6jUXZs
nLwDgkzFBmY9nBgb9207uP9Y6Hp+rpfU2Z4cX7z4A8AyaOOJ5KcIg4WznyjVq9H46oow4p7kyxHP
rTI3u7Tie8Z0NK/QzzCCVXd9bTc19RgdVUvI1RsH54+KxTdunKeDSMdwxDL0VPoKWwoHpVib63D4
pVZtKjy5yB0u0qz+nBVBmgKsmmadBBym2c5VQJnEpM8bdBOht1gqpAZ67LZSuWeLaluXm2O9MzoT
qbM0QdmLxPfPCAYBSm7lao2Sztn4xiJy/t0HYb2uQZLIptO5cy6WCUCxQ7w9b3lMav/HqIg25+fb
T4dnb1isPRaX/sLy3pEZTnxAoGcBBL7ZxtkXLqXl9BPM+8OVIlYhZ1tM4t4C4wRfWda2taanO+/i
N1RvY56pvkwDRmOMqzITrIcGq6TuRn7ihVNGzwAgbACepTYMriMN3pwiuW4JHR4Vhy7rZ0UKs6V7
rCU1xnJ0HhG/LuUmhRuQL8NdrBy3j/pqFmtXt+TQOs9GjTYx2H28V3yPlU3mNf+q9nFqXkKHj3IM
mf/CZV4Cmt5MYFbKtS5qGWR4Nr1ddqszsISAbNQ9hTZ0lF96CufTqDRhi+fjbMGIkpCdLR2x1zSF
YWn7ao7gx/vGiX9DzRxo4u3DA9EbdA472DRNLSIcs7ObgerVZb7UF/xImGwnNFnCbsTZ0Gyu8f/X
y6Sc+clco5zqNoAHaa4RMq6KrH3QLXbtbahOpGEB7zF0uU66SbcUSgXRG4o1RBf6HU2f+ucS/hB3
nWyzvreYEMKJpGzAHLh54WtNR9WyBa+bFriY3s3k/BLP0JfvUtrGMcy1aS4eAn3U+Np2ZG3cPW91
JwxaV6YN7rjptPibQhPEJw94iVNLiFYv6WuVJ5lsNhtXK/dg47uHTjC2sXBwdFoTPQWnl8PuRlkk
xS9r0qCGX5nxkX45dT5udJoCIdVB+NezjApn/dW2hrR9xa73PhPs1yx3DuzzYCgyGMW678N/vir9
RuppHwIvUez9aoz5GKbn8zPOoO90QGdWCTJz+kDb1cUP2oZhORUx2gEdEZfhf2qZXK11cRptWoY3
8nIGfNVK0q+IABzcAMgZd8b10J4Co45hiCTh3EzxzmayiIw9e44lqdl7cUlYLmxSjiOF2MCh781Z
s5qn1lVOH6PHh6NpGMKpPEgryrxrTsTIaosdcE8jZUDuPZdLXl2F8lAvVdCM/p5RNd2pnmmn5kcE
sJGgqhTM+wuFn3CgeFQqtGcAKw4Bmreq7eTFr5hqHJWNPVF7KJ4/pqumcLJQfJD6M8IDcKPwD9O5
M+lzQJXBqzZhBFiBtdj0FKa7DFr7wdT0yQ+G3VtmB/1y/zej8XCqRujvIX3jKfHDqiDtmflxaGCy
1lXkYIgE2THc/8jah9rJY59UF5iYTDG7pdbNIobV9DuYY+4d7sZPO6icuZzAXbms6a4ToEbbscc2
3iumG7rE07USl9MFg7TWtASF7f8l1BDV1z9c790pbra1Yq2KtjnsjZqS/0n/hfUDil4KBGM2DPuF
XmL5m3cKl7kA7gkAwrGdHm9MeiMGOXEjgKCmAKJuuyQvGAQDdOs+VqsaQtAKLJt8tK8mS0oO8QNg
D8GkNFbpQfk80GPuMZSS5zOqhylNGdni+L/lgD3/7My5BPIYJNWJwxzm5B/k3EaKDfQwTdcfOZJe
fILDfQKbvEaZNdcajDfcFqJG/rkosq6Pf7DTsKNcPqmItFjFli8Af3vsEi4qsAMsu7a7gK96YDYm
YeOTmBWLwknwI73be7BwyKyw3dghRwqoGBkW8u6h8MYnmKnivN2ceT0W8ePw1hTpChbsiKGLK17D
uNM33GMHH1kBzrkjA0ulAfHYzD0b00CEFE3I5wGa9R4EzmhJ32y3BmUFXV2aJgT+5vzoTsHAwCGP
79eRZ3LXQs99WaM2N/jMunvfjRhFtnJc3fxlIC4y8IXjmF4sZsPu9PG6oR0RraVSQ4mXWM6+Ozr0
GBtNKRlgEwNqgDGb0GFXR61Y1Jk77wozeOb5EiaEv2w0GvvujpB4qIKUlIQaZ2P2f3cmYdsOgPbD
olhTAr6RWdtkjAYNbp1Cco8HFgav+rh/EkwtZoznIzK5M9sflFkTBkD071RUc/pq8CLpsf1iegUm
eWcJtuo37+tEgw+qVbZYHRpbvrVzHUk2h8LzybZ2mEuFJ57LSV5zIuufr9ySDrk49hRM4GfgVJjR
O6mq5hpxb/AUGAlGBgrbjsNYOpN99vCQQyQZHnuhbuva36riUEiYk18yt8ncXQ86EmbUIa7qCcfT
w8uxucObfkKhUHnhesuSgYz0KgK8HMc8QESn3ni1IPHm2PKz2SUcTcE/sXUaAREtAfADfck4dMFF
kytS1ANw8RBQMwDWxw33RQxgBVKVyoK/XrpblHU5aIunGO4op1MlzQN1d+3yYqyAZuoxIJIlduXR
/35EO7w77moRtSj7ep7JwZtnwsZRlQop9d0R/jPIU6PHQvloirTKrpDpxyT7/h1o2qaCIBKApg/f
X78O1YofbvLIeAj88WVVvIPa8xsNhgJKy7MiwpVx2zPqzd/86bKd8zY39NdzPIQ3H3lJMRQ2IVH+
oVbhgyWVFsQDmVBKFdW+Mpg+TDNXEKFEQXVvw4unTooLvysaTQX1OpeaCI510d/TM43eVq3pgLc7
y1UnxWht+tEHEDCxUbKuMVJTTtjtzCOlJIYZ6rtzKVsuIevdtKVeCoRwa914ajZYzxPrtLHilZ4g
NLkVkfMR6FmcNl96Y4XjEAqoWTUIBl1ngt5VDQuoRZ/255k1HEZvoKxV8iFj+udwm1wC5zGi/ZtC
DgIsx3Y+0nRYuRBDJcJhE5lNjvPvf277JQmYVqDzze6shFZFVuB3HuF1GLtEJhROTZwVTrcdP9dn
1UZ1MkleSEJ3qSkmZZvp+grq9fX5CDVoC7wzrRClGFGOnXhS670o3enrDEGX8nH/1fV1LKl4ckhU
743rkKMvpfBA1qoQudhoqaL4as1RqdRpwwqn2BUrA61vjvttyRmnnK1b7BCuUM3U6VTAe2VzJzjz
a8GwHcEmrscoeIZvsz0LA2001iXhhQcH6f9Ee1Lc9Zup+oAfexGAURed8QdPkFI9/s6M4hgUMdi/
ScDKXJV8fdAYSow7u+uJ42rtmLtn+C0+qbIz5RuY+/jZGilDmomloMIpARK4z0eFt76D1X1IXmh9
3LOemAYoVOG+u9mPGwETabvft5YIfgmP0z4TcoFzIAxfq2B3lDCj9d7YNy8PlPe1DYPyyFGorqcR
EuFuvpl7Tne+r/W9MUUGhKyBMhgeGTeR/liih49nKWT8aXdGAthKrZOPVucbbbcWXjzPdXAk2Z/Y
FDfb27an9i5iBIv74VebEZin6uKOm1xiWb5rHyc0lzET3q79c+TfmdN5ni31MlLLdJf0r77cFXm+
TZ1Zwm6v3eNOvNPLda8wvebePaOSE4gLKB87fUpWuqw3Pk4wEGSOLxTLGFuRCzToNmHezwsctK0z
mDxmIYpWfWavUPGBJUm3+nRMkJ6hB51sz+QEMXGCXuqB9ycBfK+WKuGqZAcimXMQ3YK3+Ep9fTWw
9PsYx3uRoWXdCW9iSaF0zEX0yJqyRyymN3PeYQrHYoARBg43tdnUBK39j6yRATvYpEx4/5QdEyj4
+Dup92oBeL+soLYPYrbu8zyT2PF+FxKJItk1kbNCcv+VIQnKk+h5v7Os9boFtSA+opChoflGUv3m
V5FycDEnt8JTuyjp3e5IkH8fsvlzBRxbeDeoe2X94Cg05FsStu9ThHp0WFUoQoNGvxh5wlR3/o/n
rySm7qLU27M/s+HwKe2aqSczoQpXbzbH90oqVDtXArShhzduc8gXhXRcYsIAQ15do80UBWDf7jn5
z8HUDJVz89xjiiB81a342jIUoCB2PisCgsjdHljTv/qoNaH0i9mSjMipIil1MFVqiRoif46uMOvn
Bsgp3r0mnBqt80mL4B+DScbk+IvAnmj7dxajr5HtKFVIjCMvzdVrKTIGyB5hqF0MuecDtqyOuw3s
U8YuDuCcWi9H/SJfs8ycVx9fQF/lB0X39Kj2bOWkKG5Gd6ZFJWTJ/SEhDTnUSkZeo/l2iGDq4BAx
w3wAU92/fk4e+Y3p/oE1aX2fPlDb/0F/PMwgqZIWJhJsub5PIRe6QuqypY/7RjMTSNTtlq5wK2wJ
D/ePJh3mRn3zaFhic517oKE9R589rZPYsxgpyihvPmD3DtzXSl3zEKmyMGwAdLz+NemX8mbhuV43
f9CoByPpjzaQreNLBwT6F43cGORquzS7Z4qFVZm+v3l1hxh7kKdgaAai/Dc2yBfOt0LoG+A+xM2e
atxfKv3RkpfOxF6IPRvAxsWo95tUGh3/mjzZ8BJV7fa0HiuuRmoq8aPe8VlC8SnulypGLxCtHsoD
wP91UiLCHuDwOrN4qnfhdDqfSMr2YrYwYJgcEVn1bV7xzTPXAItx9v0tWJhMarSXyQ63oV/8J5FB
cW1zPd/HAEHTV9x9W3xnZPKAOLJVDoJO1kI6NNpntt3Lm5qH6CYL+z4Y1uWkNfvwXkgmRMc0HBGd
j6WKG8SaQzHUBvYsMl+vXKQlVqPQWU1i0Dn8YW3rytCvAdSjAiTFss0z98txzgx9kJWfD+Isv9RX
8DBHqgXWFTwY4pGjUP7lCijh4oOp1OQ2XZtMRc868F2Vvl3cJWg7+tsvUZeULOYjONi7zrBteIpX
9c/JTzC0XiBMn72mBIYEDVqLkjylhUSRH2fr3dZbt/8lM+CsNeBdrFuD7FN63fzgCLAy2EnTZpW5
fl8wYllE4mPkdHGzcfNZOQfzBsc9enDqA4p9RzpT05APhudVDlp9BYVqJ3d4RIsOyDNdPAZn4HwI
L5TkF8+Fgo6jtqIwV/7e/JcnkRKRfR3hbVHupMFu4+HXbjZZpqSsT/TfX9vwyqAgpqX4yAzbHIM9
F1/KiPCWNEkrmXL02E2R4oqCXK4TIErSIzC8TKhBfilLc3evbE3mp2fIautkAld1QWqIklES4JLX
8/9vEURxdB6XFYIxyzZYw1IOeVusyH67DTIw8qwUPuo4UZVKjBtdqr45y/D1GUc25hS6MlQr6x93
qA4kEBUt0r3Q1p/aQp1Z/zdmbByL3rlN8JbR+Dw3tcf1/8qkM0CGnLIXXd8+gji9DHDTfO0zd0Uz
989aGJZmkgUTRFglArvGty9PIExqStGDVsTOpuDUyYaBMEltEOhtFTkL7zWHhFhe2kc8tbkmLoyP
4BhyF82mRRXeo4LdXiwoTkmMBYxj4nni8yfIlA16/W3gNop1nc7Mjyuc8op+tYrUyRNyfxHzreRf
9OKJHaY4We+B1U8OMBXimIsg3ysMJ/I73Csi6Duf5l5YUFEhuufw5X/pV0wztrGeygMXIWJnmZSr
KW7GYyUmBXw31kGxmtGAMVvOur3xH0u/omIQ3m4KUqVo4iqMXWRyelGya/1V7sYyHOCkGIH1BTxn
YtT58QD6yvR0hnk5lLO6dCN5Ir4/JH2SIzl/w+7JpAsDDq3kYz4sRJqUEBBgjt3jMiAKhS3EEdyr
VtF71L5XdLiq1yrWwSgFChUsNYGWzN0KN+zhx2TwaesyoHAs7uzHLq3OOvm0TxvHT2OZvgpgvRcE
sc+ebOdHMxNSoF8zSiVmbcg59HxJn0zjbJ6fS41yamefBqoh2BUscu3LMMwSxX4qevbymSq4E2nL
lGkBh09IIqAc/+454WELn+FDgK0DrUYwvBX1te5OJYQJ1zR7QLNS50X/qduM8mGpQjjFyDPVanFE
9ZEbj3gwux1gqAgkH2q3EHsSmMkv2ln4yVsfdHT1zQ9uieeEdljPqCrGPOknN+h2MID5sAiGWdl6
XhnPap9C5CSp3GvRvDrwAOm2HBCnR1d2UV5AnutoUkM91K3xB4gqwLBpB1EGELqv/gucW+eY4cEV
QvLR3WKDn1mSjrztZmM3/Xx4CW+Nn4hdJdN3brtbURZZt31Lyd348GUeVhOuNLflnEs1zwMTqT6c
QtplPF+VyVlAIp+HtWh6rLEPifdWCcipg/tSoSF1sNJw9Oy9TEF0N1DvCN2+S4hlbZXvnu9P1EqQ
q2SKTeZ2SqHq6WFGXiS4Tdn2Iy1jjdl9GcbJOip8MitHcmGEX3v9KdXVUJUpneW/Af6VPgFDx1cR
WJFbjjGf3kaglCvmpdfzW8dycwDBElhEKY9zaRlz7qHp3anh7DuYNoV/QqiqB6ZmqJqI+LSxW5iD
n+QQnNomGDRfN5ad8jBSqI0CVqNWH0Rf0vhJF9AYa8Hd+tOe5O23STxFHoDW75OhaWzUhym9cgIl
1p6KBQ7oXlQFaoAyKP8vps/xPvUnlVxMxkfbJXhjK9kYUCiMOkczOT3vML27MljYBqkhxsbGVLb4
dcOT2eg1Vx2vW8h4f9hMQfLv1zBoW0h558KpgUwSLULNaWJMMja1BbeLkzJqjTl8jCPdgXG9EgEV
wQO/4CnZ6kOlxO+FE44QiDXRfsUndziIlk22LV7KBcAk/Dont29nQV6BLcJCN5+S4A5daWFImgGO
/9+Qpzoo4WFO2EHTbj48PVAKqZkEnkpCPEn+RKfbvUuU31xmPWLrwmGWrt/CIIYRR9JkBs6w2Ypq
AWLrt5U0M43h+/3rxOSSl9LgLEcF2LV8NgumobYMjapYfmtzmqEu5wM37jWBtnCib2GR3BapLn6e
ZAWsbbJnrm0qaeQrnX88+oJYucqOp4LA0vmokyrHVnz36wkF43vu+Oi01tcXeWxifOZFbjXjWcus
rMgWIlNyEjPotpttBdRPHO1qujD4ejY8ZyFKyW+TzUfew2oe/9iKydUTZiBAb3z6+Z5kIqK0sKcI
RDRQhmzfOLJsJdeXH7bhxgyks69OiHHKGK/wGOPtTVyRCthqZzRaIxaC8nKitnK278BSN+1au5wH
v4mI2J6jkcVI2sowWvFe+bYqteJ9NWFnOkY3+228d0/BpW+U3a5eZUJL2wwifdzG9fjqaElLhrGa
+AccA1ubycArt6QRjYygRNcDZkeoZLAPeRRI8POsPejSGSa94Xene+QNsjHWMcUHgW01Msxy36rx
xnizkL3nR4KlqZbXUbb2djskO9Oz4yIEhowQyfu8iU0ibbY/ra6+K22MQ/AzKe61MVx6sScy2B9r
xsS8YdUJCVy9UagYSDFdThXI/tu+n6CHV+HQEMinD3NPGdHJhlhBNs0PYrHvNHmru37j+Pf0iXRq
iD2kpshEYtXREs+fghDQmal1Rd6RWSAweJA7WUZ3M+axa3pnprvmYDbhm3gQvI1GfY9mVchgrwLE
OiJlsHKGIbCTU5N/AAhI+gM7IVILq6Q0hEAE+lF+3m3ksZQN50vt9o0XFmTvxVFhSLyXk3ZN1UXj
SBhk4+MoW630/V8VrKgrrCh4KzmqFillds5GvZVoH/tOiRntT4ghqNQmxDBlbwQ1Ew3KsEtW2bYX
5e0GLJBfRgDWvP0G8Um4W+7cDtzlyWhXGuqNh/MpBo/nrRCjOoWLCBY3BOi3rGAC25QMRA2L3WDy
WPjveR+qVCrHak9wgjPXpPhEO5mrJHCdJLWqQZrWPhk+APOD+yjw6ahxhHmypKs2Wz3K2jdaZmT0
4NtEGJHfBjkxDaYc2c6QSA3Y6y1dmPykbVsgxlx+2dqiHz8RQ9D2FHV689+uKninUETpx0GVaeWY
SalFmE5MEPAV1KhMV9oV5sKV/GIyy5z42fLV/c2Uhy3QdUmySflB1z8PGcaVe4gaCQtQF/EoNvjU
R2R+rkSJKpncDoRoUO5NsZ3bO3Ju1Jd+FFmcc2B7tlZSh2KrQZb0SZbFtTo1d1pvSuxKLG2Hrk3s
FVz9ymY+1ZZRy+6CwH58jWpyH8DPXaOZoLL3IfG1Ee+3I/nuNtp1H7B7X2gwmKPIDY18TofwVnQ+
jkYsVA4WtZVg2V7mwfyGSDZqCHDyGUvwWMZsBdsYU7XzPIg+dJLckSyHfRMuXxH5x2h+9pvznKOP
nOCXsInrVWal6T/A8ewXh+CkhiXTxCWQhN5a08dMUAQnZxhjTSJBbwrul+hhru6BEEdwXmc0hUYV
/9NFn4crstRa1YvwI2cKNTvFTUp7R3ThXEG+EDpuzySidLzNeeHvCA/IqP99uFqDy9X6hPwW6/Fj
0vuPHyGqVa2ohvojL0a/CeMWZZlnN9kPbWjkiTOzpfNFJpdxrLAACKoTnaaoQBKWSm0yUX3bDQcb
1LRp2w+xf5PbdIP7iv+mTCzm6RtFw7Lzk2RB04UFaWWsIv38uvNIyQXbLQrHlslRXIcxIKxCLM23
Yb0VWuN3m7CeWmEqrzoHYD4ZM9wAn8R0XYf8nzckdK+dG1PjVGMCf7gGANwF5hPvLriowvwn04YP
dytZe3tzMMiTlaX7MeOYcgZZgAoW1bQ7WvGUt2kXA0In2ZoDmsGNmGCuw0vWQH2HIX9wcN9K5QqB
bEcOsV4Q9OfedqVWACTBBZZwfO5OIViXa0Omu3QFVXae7dz+dPHwntdNgBsHeUQxJIgMuygY4FQG
nDLDcsO/GKKKkkUOIE/exTMlcXkaDz3dV24mF3AJqz3EnMEll/5yyX7zcp92u7xx//tA+poavmob
5cbAUa47Lq0rknvJzPE3AWnAUG/bGMexExotuLUyO5pSdCgldeTxL7CaeWm0MBauDyZLOALaF8An
t2F1zTBaDDWoKb8lxv8bJ0ouL78jmkGP2/S6WdMs1p2GYnfV3puuPD0fG4jl5UI4+sRSZI6peoSq
B+7nxtl+JV3d7e/b2D7VvUDf2gLWHrz/H2luY/iFLB+B2e8nWlhwgPwJc/sOMGvahUb0wXuWj+XE
6JFPkACinZj1KL0tLGLd2cdifTvDrZBgqPAoe499eKxYuQnQTeYzJJbi9KtCcq3c1rASBpDleTAH
9dqR8QnyhjH6a1fxQAuzu/NDcopZjd+hCmwxwkoZpcFdJWFS2dM8q+bZj5CbedD4amD6d3EO2fut
x0k+yISJQXewezAXfQXX5DVvmZeIYXFd3B1Bji/HlkfuVxG7G8/SG1M0Ufk/I1zUU/G3lvRuVkVx
4OeDCqekKPfGFW1BO7FWU0weYJBF59Pjzh7r+T/7+z4G8lfxPPAyqd4xbVdoC7kpRiqDsH3ZUUrO
7Q6Bva27RUJdP6F3V0Pukpjmwnso9ggQP9/qSr52J5x7Uy/MJDwD9IOCQhYpKUhfBTcWzTLhHh53
L4UYpyALiB0Z9qOWCZh3DNfIFPdoj4o+eAjjjVrANs53rgpE7ExaCt8U35APTgeFv6fsv2/maU02
G9A4QGGhCrOPGCriD7TIcK0rwwapvPJ22BsNZEnx2MVTfjNZNNz2QD3jNQNvph1o3uOtD4K/9T47
ezzbU/dGA66vChxs4O1pK/2lUhZdNqWI91jMsspPV6DxDRUWTb/0W/T/mIaOkkGltsZkiMhU0iJx
UgI9W9EEAM7m67UfURbZvCBmeUq6b89Lu5k008Q7kTY/986/CbOwtlYVyiw8S87mfUR8KrDL5wK8
HgHMasXY0c3yODdbrhA8zGzOAWjyr1jKGCPeaaIQ26i6GBN8aQWhWJvWArduKn4lloTYCvUmBENw
k5ZTRhXcUUjK21G+xk/Rygu9n6X2hwCULsiZDXOi02DTjVx9qrOfN9d4q1ydBrT5f8nQGvp56CzP
CeGgZr9iEf3R6gIsHXYNc1kupIrvhYyx+Y0wykQIsqAgRxDMzt4Ll+a/XY3tHzVIwpG1jFGcUgsS
n1ehCnlJPVcU9MHc4vmHLEo4Iw4EwwxSKDXnBMo3ZD4iqTcl7bwTpfiKA7vWjcE4APb3WXLTzctM
MqGN2GyZgZzNNBi515BtL6/NuYYqLAXMDsKjCa4tg6BevAXKsQBkRCBf2/RdI9mTA63ALEP6RqH4
ssYce6p48A56VT/6nnlVVYkQKGU6d4z/xAtGqx21d87UYgaTbKAHfa+HOrnokFCV3jX/Xyt8c89Z
E9RGjZUHBN/LhtvUFjzZpY8hbuM+yOWacOpYPTfDKVnoSCzP78mcOgHqAasNl0ia0melf2j0rjx/
c/huLQgRLDpLDnfArsSW/1tqrlWqZrCRG0N800iHTWLXrxO+dpsp3CZQLCdyuPV5WVuOaKH/jqBH
Z/mUX3bSsYg+hLtR66Ke/3NdkjeCNVaQLqF3OA0gdeznxTor/4m9/93RuOEc4wfIpYPlxHS4lOd7
79d7QY8XogM2Wi5Lyn6mGFmN+KzTB/X0xXp2J3V3Z2qm9yXOy38UJxXM0YnjaOd3u5kBRNAzUu+d
v90foTUHQGB/Gn8L6jzZTzyKKe7CRt4aU6N5MrFW1pV2p5vyn+aZi9+4Pr4PmQM5kUhZsrJlCH/l
NAA0fk/a765k9gTS83NeDiosesHP10Uij1QfhJPUGgoVacewKu/Gp6qlznGMar1d+z2G37jS9bg+
R3rBSI1MTOznetM9qtpuyu65CJk2wDWe5Z9wyQy8NoEL4iHYHhovG9VXYpIqyD4ZvRS2LZsDnDp4
TQNAHwbuSExm8JLUWR6qA4Kl4AbSkzBeNnU6v9f0WiCrEckdifQ/5LzTLA5HFiYhgJn+gEJ/AVBU
RUVEy07QlMPFywxC29tLB0+kjPI4egrm49z/6/DDrKMi4goJvGteTlztulsnw4PL+bZwbemHDppc
QfzbQQYeRHYCJ6xCr6FEydx/kHo/KRAReKDtGn2kb3CUHm+Jrq8oJ90vrrz5rhpPWleRlDQaRniV
6SuPRb+MMN0gSRDvCEvbnkra7gTXpmyezuF+LoMkbnmHUjBe5wJly3yat7XK+U9gaatC1YTyKwwK
yArqxbvUN2Svadr4K0GP1M1j9ocg0ZI3/VqLDLDh1euNRsSHjMlCLkdBT8RLZCo8lnJ+TRVbpZ0l
lG5+5Ni5tHjgn6xkcRa/mBeTQddp7J01L8uq6eJgQOHyPC29frrjSiIJORYQZM1T2puyzVf7FM08
A0RMSlyyooqtrEd9cm0LPcNLBRg+p50WFZWwlxb/m9+LF5dN2tzC4X4NypJOFQz6/yLUH6IOB+54
tzpeAum0hRBc+1i5ZWCrh+1epjSCE6a4+7YvMuY8CfmOVKztRGX+6p502yf0dKjNWOibV62XL7g+
yhoUfEAL0Ou2SCrjoEscm8gfv0yt7OeLATjgWzWSOhUK+7J935i1epROjafu45GEBpLFmKtOYnnI
mnloeoFgAARq0YSUAxYQ1nOw14MyxBuJFwCSIzN5xK7CENUGAAqnyTfhmgUP5WsRFHQJ88BSF+bO
8Cn7PEm/h4bp/IrdlLtUPaS3KtWrQUvqDf+tjkd+uczCJz5CAyNqAIjSrthvHoPQvuq2Rbqpq1cc
J7uoaY4Hcy1gr/kgDhPPXQnpuu1438O96ZlASzXqzt+jjqcaMxhkdRvcV0JgGlL4ttKyzBP4j0Yb
zXsVamfU4JdSRcilhJJApkU9WkQLOcrV0zZgZ2H/+2/1nVAmrBvJkTNILibcfW/q4pgwihfdPCvz
thxCN9xsSEfbYFTBUDyQu8MVXCFQcTAQ6P8Wa5E9OumAmakH0U4wVytbkjl07x8YQiXBJNezP6CP
jp6jvyOioYThm1RUWgKG+REarsRUGUArYV/iPA90v7g1T3BoFGU0wmr1vvsgkKUog3tl0TeN2Rrz
DUi1U2Vg1LAt0+Nfe363uSLlRJvIZ1MniWcxCr+Ith9/Pf0PsIbDB8oy/MYrXVQUEKrJXo+A91Yu
h5++phpr4nnI/43hBV2D6B6y3Cx/eOE2vKGd88cUys5rEggSU4QQrbsCD4TWQ/djDO1QuVSSnuVj
oeJxg4dqglc9I2vkg6bVHEwWWx+10LEmsC9bIqqliwkbgcgNmShUd5Vlp+CtmB6JYfXYa35EPg3o
0suPmAQYOxIdsnMqOG8yTyRIWj75SoV/yC2dk8vfwb8Lui20g1FAUJaO3G7wTPlxjd/RTCw+Dh4m
9oC1UfDKg/wtn0wslQ4ycLVf/HFZeed8xh+X2gVctXD1xJXfgZeSo+H4NbtTz/zL9UEjXRjbBO7P
xmMzGNcEna3LR5o9ByzmuhamCax6MqpUCkBpghHk7f0d7NnxUxSvojIO6/lIzKIVPiq/UhZ6caEB
qCR1CXfmKIzzLqe9K15/SSkRZeiqdEjA38OUO//eU7Y57A1KfyMs0rr6Pb0OuzudW/MaXsBz0CFi
bqpr21LJCDAK/Ih+LCNovMg9Iqe9LWYH+d0SDHegq4plCRLylZkr/gTHbdjchRAkLNpqiZ2dpIIv
bp1zHwnV261EVehtp6OtaNFDkAn/0I6iG5Q2GBKq3FYmHlUV7TYUMn654bYELBdS5/MvWIcI/Qjo
wpDdmkiM3CPTDQbHmrP+OeahMfmb+r7TvJ4v974BxKw3Arh1jbXAfrWej3xvCkOwm5A5w+q+InmL
FQmAOWYxXEbStVWOyT8gel6wLroxw5Pmpb/Jjw9wd+263DAJVbQ361r/7Dc8eN3+Ke7CAeBaMqa0
LsJqyP85FkxK63fKpQ3rk+WhFCBS2J1l96YwwlmQ4PoCM05bONnc8Zoc6j0lKI1LjW2QRL1CMDtx
I6oT90ZSebtudz9hNtUwCHAHZXXhtepRbi49nrvKCidJAWz6FvxY9oB96lIjmCkvfFDZ0/INhgib
MAnj2ejUCF7ejB8neE4+ct6X+Dvf0tOxc39TKzg34Fk03FIXX7egk0M3WMr/MyypTf4DJQLHXQnf
2Loy8us8X96EKx0v4H1Xpl3l/PzfCzIQTMF0e/BmP9aE5jeMNiGvbm2g7uArMuauhTYwoy7QBDuw
rguaEwucBRDZsw+edUshBTY1uFtqwPtQc/Q6cUZfXwyNEB1ugbg7AOlJFz4fuRNEPT0jS8NThi51
wyhd33l6sydQlfibSO8RK141KLgeSDJShhul4qGSh360TYOulp9+iwLZx9C007lBSM4FOKwY4Xvt
T0gWbRX43WVKrG6NoEoorSMDeEmic48UhusmRkd1Z0GgpiwPV2vZmdj6d0D14TB1SQtHwemWBdBi
MZjP+BkVdnlFZjl8NCF6JCULgMflqdkmcTdF1JV/7Vqz52Fo9d2jpyirazPm6vSlXVA7vtJ37sc2
Wx6hlufRiLaZlr5cuX0k8Nz7sKtHvJ/muVxzBkymVKga0OQWP6JKFSdvD6V6VQBHcWLSCEPJp/97
gDxIxYm1+YLd5Mfv4F1lXGNfTxak5wuaWLlhGVI06rkZfhez2AIW0p1WApfCWIakoH040fuhWc8B
TC9QVepyibl2Di3z0/mvkWJbc0vmtkDS5g8tcGCTNhIl3J4oRaxPLkx0tsWaBiG/OOzra/cupYKR
wKSaKzmwGrit6OwgXNqZg5Zxp0LmhFX7YGS2EbBs7pbMUSJqjC3DQB2ZkSTAuKUj96axSFx4U6QA
RoldcsRN2vqy9LCyIM+8xKTJ8reKMBe0/YlHQMFJYvw7tP8wf0b1cR9fSrNYEvnkT2v901EHFujH
u8Soj64TOQw6eCYLUEDfpGEa01ywfNm2E39p+m39daWUPorqQBZcrjY8bn9Hi3uCKeDws09vICU1
v4prrNsY31IJ3J2e+oLm8t16Dfu4jGWBeqTY7ZqYtP0bKWuFNokGElPqt6N9ONmvzHlo+A9eI3ZG
ALRLh05Md6nT66KJWDayHxSF66kmMivzgtO9N3933sFeGz+oJpx/95TJ1MlxgbBV+EGv9cFGt1dn
GOYJ/HjEnGvtZK1xmf6NcW177GVugX+pKeSxESzStkASPzk7N2hBJIe9SOg/vtyqBAYJftQFHaye
9yMFVdtFTbpg2GB1m42DvnC9cNe+3I/MBid3MfOLhTNEDtcDkNUp3NBPDiNNboMk86oxgXnj7/W0
FrqI9tmlQomeQFX0UwmODm9YOlt0vZFwJJ9d4pxgQQc9kckY7pnuF4L2WP1Q674p4flRnUPP7Qup
AGbzQI5E3AXqhWGi6A1AWp/6JVoArH9qdrflcLrLVpqS5sLOlNZemV3tGWGyI7YFXLaO3SW34cBC
DWb69dk5YMgcfKlScfxVoDrj52a/DpXXNd0LftZ7041LgocykQO9u0v58hAl1Uz9436Qud3xMRKR
EvmtDB9Qw+bEvggbEjDS23KsecMxVlbArKAR7TR/HfjHe5R9Bxn2g0pLTBCX1x/wUwvbMla31mJJ
9+UIAq3CYSGWCTiYqWOBZDl96I6Qmut2zWN6x0m2X/cNYFKLjh2lIobsQhzuPp0coaV1sbMDBF4M
6NFy9HDNnlbVBrfIviv2bpGjfBQL404zg6gXtu0uNKhPq8mnAJRGD2u3KZhq1sWijOKa/Nneh7ZX
XbW/6ZVDqg8z2pStVqMdbLuzX5SYHEZSQCXBp/EDLz6h5VbSCa337kM7DokbqYviAeMcenEfV+7N
AGuabIF90qQIjnmC/0XD3vjkfvImTuXOx9IwPAno3PCkw1IhcQDxTLqHXSMTD4fCPpF7gbi9LNjH
ajTG8oHBqnmY+pdl9OaQbYW92+NO9HkNGllCOgq262RiTqIBjRpgDZUYB1zpCrbNF5MPsdLQCA1Y
8zjGD8uz39B3Hzt8m+TJjeXQbcOPWWLmWoCADRBVkQChU10conPc0tuMKRHewH00dys6HSlPxKsW
bcFzrhNzGEpQJGds7A7sw2xdz6C46ez5DLefPLTfq0UZQsgLGM+kPs01RRxO62bW0POkLjjpqSYU
RtYRKEimFhKEFIp3xjNQISDkP06waJzKBHyV0arA2PNezGnojI2imavwS142oNjMbCHCLSDGB3m8
H86k7BwT+LW4jrCKefy7u4XGrrLQ5k7kd7sp3W373l7Y/kguDao7cBrFEHyyR8doDRFIjtmuCkTd
GQTcCdzmf0Vmx7+/4YoA4xqPWWfMukq3olqEBaaYI88/QFUi9L0hmJJB42VHysI0AH/ea0YEFQb7
7FASvrOSmksOJdVmDVoHwPUtiwM2BDIu8ay8zdlzIdfBgLd3Kr4r1eOIlXGHgxPm4q0wHGcSVPuN
SJwY1VclzyYwwQbY7O9FKDlKUb+1WTe/F4DQirmW3NFm/Ut85K+yyezVP/MQVl7PrS+4Qkq9JBAj
H3dmPTJ7KJTJ/JRLhcYBSBQtdh6VmE6smIas9lLe3szsEknhgEOTpsHEc+gT8+5Uebjql/cJ0oEk
0offH/tufAf/wrtfIAcExSmFWV3jHJyGGEvHFrt3oLCU/mpeqAYcyGbXwrJrPr4RdkFP/I/ZEbxs
DWNMHfKLeWIzdJcaGtbzmOFxpjKKPzpO6HbrVxMjeBnbjdOKqTxNI04xj2FpPLzn3A2vcd+BfaZg
KyyA00gJhq0GCG0mTEdS/Z6b7zlOICWY6fxhVfOzcK7akwi+828KvelHIYIdwazBaked/P2R8syK
o1kGOQDyOL8tXPRLUkuLPqYe7zGdScZ2N0/jy+OyLFSGWLWuc850MAQ+DJ3Q5mgHBtFMs6FbxTFr
GFUm1YQr2Am7ils4Aee+LoQ+NQfOPQwx1xgiZul0OhNE9O+qBskxS6L5i70Wiw7AA7k13rystUP3
bxkJy0eNOxclY8PLEw8zEiBGixCXp+HuW3Ei2U27V8LFhpf0PNay6VJ7sZySpYeMRK5VnRATWuFs
ibbsOo7EIPE5wslhVJxX6VGlG+MBplAwI3/emZMSRhLi/I6nO1L3QU+1e+jPddTrKXEoZtXypnGr
Vlpls568EEpqzUVEr3C36V7vpwpmpgkv0p1LCw0tW+ei0j+oSbTLW7YFXXcoicJ4kzyXyeAUK+32
IrCpJ/kdqIDk6ohj85DqUoQzmbkD7aiam5q0SgxGIXSj0IJfjsh2hwShXIJ6544qx6KytZmgRbOQ
5X5woSZxi6qpNi1GwJfoUgr3hLkXo839WWrqu5zjr5o5Ryle1Uj48qg3T9WCszGXSSOW6KG4TkEq
o/wBIpL+yNhUi9Za/QpbyfDlVPIpvT7yEEi+b5/3Gl4vk0RNFrIk2as0F1CPp760l6b+hmlrFmCM
xMErqg0yxHiGw/3w3NwM5oRmUoYuveRTCi/XZRqpOGDkv8id4XTfUleW4XwUdK5uy/UeqA0UyyIo
Kspr5l94py/C7NAG+2EqYpnuNLtml5gAj+V+vUYRPPC4D/IeNEURB+7M+AbjVTauNe+9r4l3YDEt
M45pcQ2nu2wozNO3Yt+wzgP54QdQT6xCrcqDpP7uC0gs8CVAZjschv7ng7KEm1rJy83VzlB0Ktzu
77YlpV/EK3XsCaiQF4WaaGn3R9rt2E7cv83jaUOXUmiwb78U33Z85sTdTHegYQPxnIgNF5/S6HSs
Rb6wOvYjKA3RfJknDhD32ol4ZT/gq1ohfC94iRgLJXmgANLNpe13G1HGSBEAhEBfqzXQ2CDIRh0F
Bpn0CkBQNftaBaFtv+jjWlLxXlJEiKGzUXf789B6t86POhudgTc7YxDoUxTRuyiJ2jykR4Kl5Olh
lqCrTaXdXju8ZzatL3AJ18lGEpMJC+XTGW7EyL0IYblyWZaPmH/a1SO6uB01Owc6+ckjJCfTEg3O
rg6vzS88DxBZdHDNXf2KwlQW0oW8PCuUa5wxSGH5+KK3Eo09kQfUNL0L2jbALsD3qb0/cdyH2KvL
cnnLhF2UrhWqCkpBf7n5ZS9V0h7t62zZQayIg0GtKTokwfCZU/fWqwaXjUA5jQ9lXemwc2bZlO/w
WQKkBY3OheeLgEiPdUDIWbdy+PtDUFnBZs0MdMCLp4AZpjy/x7rQ7F6zhxYLux+Lhxrm2QiZ5YbK
yOKLSGFshsFsKUIno8KrGqfl8pKN1/CXHsfb2qQpxWQNuCFrpf0vnySr823uLG8Jwjw8brHugMrR
hR6ULTEeq6pZqySBYBgJ4DiOL5P8bK25HaXdxWA76mlX6JnEXwq00lkqm/+cyBPDwYca+Fiejujo
Baaztj00VOUlHYSDWZu64wgOqHoyusKtCQtStO1QXTi5Sreu1W3DWj1oKgiVsx4pjukQQeexedBf
rhtrVcNYWieZfniNlQGOpTOeJbr7iAe4d6QfhL45ACaaG2K890GwWwPzahvRrCXzvzK46eI79FqO
qxYMMpny4iMdaFN77jrMeFX0l7YMmMWcOjuF2LFeCMNCVuZs0DYA3ymgmeMV28QPIuyMObb4VgI6
3uuogS1JP0HrTe0PrcZ3Mgt29ZprhsPKI0hGYWHF/0N5dCHWLF601d8fK2XQWxmo8djArvJAqkkp
WfZPFTpZoz4q2Gu1wAxdNsyFMeFjqbln+h+hfxnLWBDx0xZ5P3TkIpt8gv49qv96yBXJKq+rOf3g
Jp1OdZ1VTYYmrx3b3rUCaElUdWbUNwppKoQV7gY5SYbdCcHfXZQwVxvxYfrWNnYl/bGCnnrWO6+o
vWHDSBgRZ9mj6Q47RbZkprno4JhxTtYFiPPzq+kPYMtTYQEXXo040R2NbMVRJItvaUBcQeBu1xIT
NLKLmiLtbnyG+hI+5HJmmWOR2vt4agciFyatHi2luWPYPeAes9DRK3Q7coyOl6EVRN6L5Q9YvsCG
RBj5+BRvxxKGLQS/WPvSsMbYZXKZb4/xPVZ5ir8rUnfjx+zl79Cru/Q45REmEA+jDn14fW4xvkRC
J0xRujYEISAzBW6MZxaTiMrwv7iiCpqrKlu15xd0XEfgpLqgWhobU+6J/01RVRfRKaidHHTmT2+a
00SFFsEcdJ2tmIhta2GR/zh9KBgKhg3xvN5Sp97fbYhOjt7T5B00KmhOTyQZQCrSLCRStmTUQjne
lSevA0ZgsiJeAGpx3Jzs/tZCcQ0Dbz8akhF2CPlhcpuW7xTmBU/e6hsLX1iuW69Lwh51Fp1P7GrC
Vw4gDjBHZdKaadDsiaIpdrrGJDBqlPtQvBQxWymOTF8XRbRgBxlEQGuyT1YIF6BoBaJqpcTe/SV2
Oixu6EEUSzQ2dH6xvyedlusVwyN8uLPgelWBftVTrn/g2iJ69Y1L6pMvPKKW9peWAsBAnXTT8rFP
CKLPGc/HkUspk/woIX5Z3sMrTN0MTuOxNx4tAk7CYBqRIEmxNriHJAJ0HNUJs+EGYh/rhH55+sWb
1eKySIEMbzsbI0NJGt6iCDXfkNUQ2JFWI/6gUODN7OmRtI/lExwCOzoJ74SYt8rEdov7Jr5X6c25
YUz5J5GOKti7edc7dVQ5vftmefqk+NKkg2IrOfKXVnjmCG/gK3ACX1jHU2n2cdh2sJwMxeJiLWf4
nRuy8XQ9Sc0ip103xKWDueslub124AvQsWPyi82F/LyjgsG5cn8TJLdhHDP6/xKWIE+Csb7UeM/Z
TtAqiFOLQeMd7paEO6bIToMj6H09Rxd4MYxM5LxqBYjiMoQxBd3EMb8Jx/atsjj185W4cwv9atu5
P4AGT89UF7wUavxyYdUcw9R8q/HB+QZLxvdXEpNHABrlMrGsSvOZkvS/xXNI03UocyICDB+60gA1
Cz++GNlxvRHUQcNwipRyYK1PVrG9XQ+VmylIGZejgDFME80CQGHhSYKTkdWHB3/sX64fU5RQnuOl
lNl6Jlv50sEEVbZ/wasY9GNagVqo7mVjL6GNjU2hTfAIFzaKQKmifqKrVacHcx5d51cffP95kBdc
+0uTfX7LgLp8RkXzwVFeqUSpMDywPmKaJqHElkmeSj3T6P1gPF4q9tWJqMsYyA7E5dZZLWyjkhbC
hD+Mcu4An6FDKkPbSwWx3OwFCUSqpoFIIlLm1QJxZkHmUiAlvuvVV6J7IvqPiBjIuetLkQnC3SVX
DhswyqNrt60eJeDjMBPJNPKxy/HvOSth2ZIO87P5tBn9B5WHWv6Z6GrkVdLpZ7iVNFdo9w0FwCye
JpNLV+2DeaM7clNk/T3yE7ghLvghw9AavsU6aM835uVKx6zpEcDK586rdN6UFlKPwD93NDnLQ4Aa
TbnSR0FIOR6+XRcxoLU/vBbfosiH5A7XH5IE5AQO/hnVI+lxU19RGnZT3bOZ3XzAZsHuJMeNXjfR
3TIZU4tLXhra5VG5aTWWKsocJg/BUiMSSCSH3JD7dREC+tWc4r3QvIVcGhNs0oP+V6yeorjkIjZo
cgwiroCg4raIM9ObGs/Niri157g4UWNY+BI4AC/YxNTG+C7oKKvt1Wz3F2fHv4W0oI/tQY3AB0BX
f3HV5+9F07UW0B94n1+LkyP5zvfUa0BXV4vjfjqk9kfNwNwXyiAVH32qyYHc1eLf0S7dzV/KPlvV
PjrnNYfm3qnp+mXxUe4339oj+jSaZHuyd0wN3P3i2UeBxhMzB/cIpv43bM37ixTIbbMbqh27CKg6
aJ9W2Xsucd9Xkc0/0dTUfoOUouPZe5EllsG0XAj9ZvKfoc8O82/Suh7r5Ze83fwbi6sIXllh7QbD
cCvEQCfydaVOhmPeMDo4OA6+PdK86kDpMT6tKaop7eIewoV7+PWqCH7A7pRanh5uCOKQm8cyVlpc
qpsPw5UEIriGlUm4otj0g1Rw20ULN8Hxu58stpr4T59oI3LmCDz+w/XOywQQBqQW+tt8QQKh42eh
YyUehWCZzqhaK5nC//sNEX4dr7+JTJ7KHMa9tP2QrSmxljx3zo2mFeD3A3u/t99FFGIRSytHUgPQ
ZteiMnOCwH/CXVe6mxSJnAJV/uH1T00ewtgPT2DVBh5AgXkghJw6/TCzo85kecAx9rtjk1G2LhZk
vKBqf3Ie2BZZEwH3gnKFeSxfUo48YwJFoIeLzTQ2ab2ri3+IbQz44iXq0nvbw1lJPQ79/jYmPO6u
UjDemGSkddyGl2h+ef2VKyWl9KqheAAOCXI3suOIWWDz0EAWCq1xho4C6dSM+hJT6eGd3mYBvd6n
addZSAru0lau+o8OE3eqHJlK5m5NrgGBKnd/whC7VVg4ZZ296cvGqKwieh+RLFjlGDYji1uMtrqh
4m7HPbAbD5BqtTD6lsbVml+oOdFH4i6jOuo5nn42Cw/uCBECXH/mun5qnWFkuYdlmQ26M/A46NB1
IBQkzU3vAT8eyAcPKMe9zMFUNfGdRMmbmUoxNqYT4wfFNu1QTTS052aWMjWRScXZLM9lUzX+NHGJ
ZK4Ivc/6iT7deBGhRWvb55Nd28aNrZhukqvJB/eUC4EdD1dYzBqgCBPYKXuHO08sAs48dXsDo3Sv
v2+E9hafCgOnoqibwa1M/4DtXX92NqpiEklxJNY9fL/P78Epfthd5/yBD+WlApbXKKy93EGed0kv
Ta6UZdKmYyT4bEhwPR96doAFH7VNOOj4BifLksL51qNjSD6YEOJq+MkzpL0Oy2RvcewOWXxrJ1oE
lvcdDKIiyTs/CQUuqd/xH4xOewE1mouHQgVfvIMz6OCa71B7ydS/lYI6ALTrJSgPHfYybT4CY0np
vH+60qslC+ks/6eLgj0mKHAgDatjKWS9WI4gHgVy1HFI+XLl1R/gT9L5M9Mdy86RqR3EsRQplDq2
MB/esENsEJn/ck6iA4QfvYqclsEeDyaiaxZiGoE3zNX4Y5l4WXoeR58XDu1U4wZ7NdtgPoPWf3+s
+XBIX6z3csue2X21tI8CiOazw4/2xZucHKp5sv/M9GygPp2JopCdfUP4KxV1vdd5bcTyQwDDhf+5
LDNs304BrGeixsL+XgRdqyjA2RogGyG/EhGMqHO+sTBytuUetpWreQ/FNs8r8nZlttW2hdTPHFct
8mZmCQIv5lB/+IcAG/vxCUvOY+r5XZdVKapbzHA3JVKXAbY41UcYRbwnzB7G7Bd3ebL4NHc6VIWi
31kp8TE+uBdyxQvr5nxyNzu7zHXVMF088+nb2q2B2Dn+rAVcbd/DH2vPPk/hfr416eiC4qQKRE8x
Lj+8atHoAFKuKUkVA9xr72zcHWMkmQMkmKgMge+4mDP9G0qjYhsiIKD5g5SZTC3jCQeScP4D41y1
UivDh07NpTNaTTEgEMZBCxUWNTveGKX1LCzU5q5JBE/+v6GGDdGViev2GjKelT9mBQUcn34ACkGR
vwqX5sATKKdQy6gZhivWK2xKbh0r8t8g/4cqZfwvS1LYcUHuYlFwryPs53+bXJQCqsQK0GhsgLJx
YpnedphHpdF3RUFk7+In6OvU0fHbm6x28BNS3H3yttmR45d9HqU5IvhdsdQb4nQCU+jY5KM4cE50
Yk+bAbsWC8y5VXXdON4E3CSRo1fOOgt8RrS3OqofkVgN4BiRZRnwszzviU0r4n+MJW9Mlzo7BXOr
wNjvPZpTcqYBGIQVxfi7hfzXu5//FHyxb2jxvgu0rpC+qtw1WeGlN9RdZ7CtgafgOzeYHHKmLUug
GSbuKI+xFMiagcQ+JUCGX7y2DRK61y8hFB00xrwH+2Aj7YsrQ5hJYTOvbkLVNojeR4FP9NgEk/ek
njPrFppO9n83sENUM75UcsuThXXxn1UE7eV1dPxSfKkmFak86ieTqQMmUdLmPJz+2I6brn6Tjg0N
D4U96ttdEjt1UFzoMZICvBj0DzQNMN/8W63q6s89ksfzPHQd1MEofZYeNXvDiJJR8/MvTVrecFHF
xNCgog1hrJqBor29jNmFsq/TdFQqQKqihQVs1IqCkuwzA1uvd7mbrBvc7rnGaIqlpwTDEPkPnA2o
QXUHYYl8L0rYF4h/AspJ+M1mr5sJ/epv9HTivjd6EuSCKmvqHVn1LRxISK+Mg2l44WCwQq4P6vnB
cdXNcxlj7wgy4eV9IzWUP3xS33yVTctdCg2ozXdAMP0CZU+9GiahlmaZVidbbuKcIfgGp9YXzC9Q
GX6JJKx3RfYfODFPq9IzjbQNmZGTl6RsbGNxPY2rur+0KGgkKjCnZTFrEFE6vqQRjPGgoXxWe/D2
JU2hTc9vNZJsRJHtJEcKkHs+5TevGNb8WidueMMkWdlni0FpEaxYcJiAfRt36524JUL81Ga+Gy14
lMSDjerI524YR11rLeB6Ug8qh7ozzvHCmzjLxuQCx744BsXBZ6WaFp/unj5a+K+xCt1PbrLPrZWy
S/0CwlwtFnhAEQn5Ae+9ylrOOglx1Xi4MDV9fqqDWPan8H7Pn8heAyAHhCItEMXB7SYp4QCzqJJ6
zSx7QZPma6+hTkCE51PXJHa6vr5rWSlG8BenpcWkJM9DhyzsqNzqbjOcjKCDwj9/pyLQZppLJAma
KnT7TLHjHrBH83p3I68pVuBhUNdq37vbb+MDM1pjfvJ0fs6R78xcP0Kr3RgyewqnO7SOjV0kj/MF
CQXXRACHicDzOMT/xd5gRVy9iT3M18onD88gWObEjmOxjWt9NhdicV7cCaCdQbNScXn625TjRxlW
/etUNVsojB7q+flr6/sg5JC6O+lcRatCrT2fyssDBg07xc5EPJar012SFG17xxQK+ZAWJMy2jO1k
TkkdegrLKpqlMM0s0PVbaJFz3tLUips8NSNcS7FA2Qrpv58sBhjS7iLRLXo2mcN7a8Qq3XXRuKkj
ca7yTnvC+3EeK/lnWcmXl5WZfOZJFT9UzXpaYHedNvH18mrzDFwszrtCR+Swx8ZQbsfVP3nc3fZN
wzGroXAw4Si6nWtQsmk9H9sOsSd2V+jFA/MT7OBoT50wk+TYLHHFX5GIIKJkzg/GckG9PnD/m88q
C8DqPvRuQq4G9AbH7/16Ji91rA00M/eyjTfpEbCiPXrcjrXyR78Fq9xnYqid6VC7wNL/1b7F8W0M
YB3TV/XaVRa8BAo2yrHOF1s0LxPODRSpMA8rwFO2XzliBDlvUmqZl9KnMeS4l262Yaq8Tnzn1nnx
PtpIx3ZH/FIUgm3A18R9GL0Mgb693i6dnY2Lv0WtR33Tth+7N5rVXdGt9ElfAwtyp+ROpqbx2qxA
Jl2lx+hgVntPK0crdn9OnNj5ZD+Dhlkb6SGV0mdF9Xu1XIDSMbms/FY0xXlr2NEAuLTMDnLjPJcL
gbiEvW3ZC06hrSDw2S+/3NiuOARIuxSOh4oV5Fb8vWxuQq+nk5Ixv3QT/upso00AkH8YBmWNZj8W
dJjILqk+xCeS4ci1oFCPe4V6/yMcweIdH0VjIXs4awcXzWnr6UTS0s3YR7X5QjBCvJD8uAGal4AV
OvRxYKrzZ7jmjBaJJ0MmVy0VYWD3fgdH5Waf2W0/2DkH7gSG4sxO0y7pCaggZ32/Bi3b4l3ky1Fm
f7hRdBMA3mfgSTCtgQvvmlbILbuNVpdnsmNg3kPbuaZDJqdyeobAPJj2+nwWeDJ3n6Hfx1xyZ5ds
XL4mP+ecHD0CRnfHzxkB38uDE7SY7CLoIjONlMTDpAIk7uHe+fDH6fjoqqmmYpYLPTu9JffcOEad
zi+va0M5LnipRDQa0MOQCX7WKZcH4/3mH00VW23hmC/z1ukahCg+EbTN8YTelCLdI0+iY1Jb+nVa
4Hveq+kEg64anM+poO8VU/L9vj2VPkVHTJVFplle8bcYjO27XjbqrVLBRutgPR6g71OOtV76iNOo
9Y8/Z4B7stdxiS5srIz6Nj7sdJDVNLtBTJcIIztw0ql783c9lqVYrGd5usYFDHNbcfWwCqUkh+eD
fTUgRqRN7eQclhuds2RALqSD7XZdiz6jVB/aph68KsBmbUeszDTHCO357xzUNKyK3s0ySuymLwHt
6vTunBygBHBYPvyDSdw2AmBfiBogbRz5VNCHfRccCGH0Zd5dDT/J+GmgelL88jlbdgUXhAdam1Yf
KX/fzgctar4Oxiu0Kj7O/B1idkSSmV+v1p8LjnTA9ZYUw9Q5NxKLgBoGgzkwIFEQ/oCVq0aEuwhd
O9watVTxZphju/yeLTkxjKyNjfeNT4BK9F2w5ZKEL7tmshO3iZS0e9CFTW8qnTSBkzoC6PcSWK1D
p0COWo0NvTvsxG5P6WHTrFmt3UXwNm5YJUIANP0kIo1rDVS89ieyuKoJcvxiSLfKzjq35kDnwjGZ
HfjJqdH9bEkYo3Goe/OfeOy0CVD5NRXbdFjUcBYKma1auG+n9+o+fWd97TLTJgsaUpX2dY69Fesq
TGUMm9J/w2YFh8zE3GA1rP8FCk2ol5zVDxvAL4E7DHcbO/O64kA7veHj36fZbkjbE6g75/JK38s8
U6obX7h1h5+oN/zqIH3J6cmuCFAr8TJUIiLqCBbqdF4UBoImQAQG9mKZyUEhyrgjwR6D4oj7Xjy+
w7lwNwgcRTVnyuqJF5ZuCMyJAn40g3G6kKTqFHiR0CjAoioatVQtYj5/Ui1i5NcSeqRT0zC7vLJ6
T7+AUXkRiEJWZgDbtxRh7pkzGYoYmVHSagHYvhgTknte/KyzOAaGBvNMD4ucyylIt6X/5ras0t27
9mZNXrnleCS/iJsxNzFLEVSrrKGHgb+t3+cc8LhDFjYiaYUv+tJk69U2ERWHfhkscLTOd4YV9cK2
XwSscjO6C9WhLBaUyRzGxZP3MWQJiOEJF9OhEG72HJaCIsaOseKvcU8BkM7sYJs9yQIMTW2nEwZn
Ch20fPeeDAjLAKqP4gDQxkW+cca76QcnHPL80rPqHRQxmcUozAvp/NfdVtyt+1CiCDdn7SOdKPk2
sgP5IlPNt3Ir0IW57oPJDq+xCyDUG4XSckZXfoB8zPYcQzx7dTgmxGjUu2SOLtJs00ZQMiKTFAqw
XTbGv6v/Nk5lxB6yFzy/xTlKTAydqG+iMAlvdy+Yhx9dJ8yHD9ih/KAKybjQkTD9D6voNG2g8XN9
QJmzajXSIAM/ZC4ZM09iwyqGqwyPc5kGhnW4bkJCxbjIyl3ZqM/Y/I91ivdoxJvZXzf6CzSy+kfF
26MF+u15VZ39zCgxjQXYH3vKQZn4I/WAHcGy4P9CCtDDvGe3yqNa7C81aftx6jKU7w6PLfIOsNyX
PAli1o9zCu08J5wNuyJn3I67BisJmmxQx5NhdEcJM1GuiBcZ7mU9vLbQgFDEijs2/QX7AZWUr4eW
xGl6Jwgo3ehVZC92NxSe3900HqlFKsYsBLdCsFrQDSUsrizyikNgGnBne+u9+6thZXhtI4MzOQ86
ZjzCUix3ULVkPk7bXUty6Jfu4mktTcGcP5Ixl+u8UpedcgsSOqYQ+uiex+QbGuA9mtuR2t8V2HOA
lz1Vq3OrVaUqsTRXppuGv+D/mldbl/n0qiSEKHmCpSaCZKnBfO3c23GFZIdNXskvvx68v2s4R/dv
xytTapo+Ng9YY8NE9Pm7WveuD74ZsTHK8NvZdNFUH3ui7ST+EKYxubnERzyT2/nY8N5I5n/HID3m
WoPUAAU2VXk2fAAiprsfP3GWvTFo7BDLm26ryQDNbHG3qWgaDBICbs8QMDSpexJBLesBAo18DC1w
ij969tQDxFZcL4nQmg6e8uy7XVDU8xYjQgtja+qlJ+bE02ClKATojaH//mt5yk6MqmfeDhtjuRsP
WfQ18kLXoNn0SbwPt9zvK8ROog/W7aNvctYOB5Ay7EkSHBwEV6o2z1jXeLVVn8js2y5xEHsWmNRz
hRr9aZKMpEHr/V2yOTe0xw6q309kvV9cGBfHZSeXdnKmJDfuddFJ4MsyuW3v2E07AU0qav93yhbg
w/g5DVMfUYfqlx3ZpeQw8NlC9zDQf24PFcGM2S/CemUXbe19PV/DAI+7OKHu8/QR/1AyyKkXImnd
5NbI4nSBetmog4UwL4AQ0kmN+shWiktNQGgOL/3WDObYQWyC8DRV4XTBSZ8tZeFBHO1kF84lXcr7
kfUl0TJEJPBiEeXXdIsBquLQ1+wrxG3A4qPngzVlKErvFZGUFHGSSdE6fFGn70jdfjM5jEGo0kSD
Lq9/ppWNKU80l5zRJ1gNQ2uTwqi0+8Vxw77oIrZb1v1bsaBeK+zv6VybhbiRIf7QzA8waY/sa2J5
Ca1zLF4EScA264CEWDiB6G32tnmfxRq+naluEjvjw8JkTVmTks/GQ7qYigyHyI2o3AFl8tVCVT/5
tLr7+rbHPeiJo0zEoxdEXcpdy/lYIjaLFiJbS24nklKss6OJoVsFyY3z7DcHjglRp4BEyEPKohcx
wWRDm0MBJerf/2wky1TEFMZLKnIiMxgqIZJpTsCweFBZVOJn34fz1J5wNfqQRwVumA3sEvtF7J1/
djQxHjZRA9XBIqlldMGrjnhFiVjamo1sTyYv5u/TO5ehWdzq9S/SX5lx33nBSKGG0aiqxWP2p8GI
b95aWs0xsAiQ4V8MGaryXTJ3uE3LqHFxPIjLs140s79TGvTWLwqK1r+fd5oTgD3SE5So4Vk6Esk9
O5V/VeDjqpM0NKhdWlqKpitCPqnkIkZrBdwBdhImBFD/CBwRnr+e7PqPLuFwR9fzHBpl+b5LXboU
AIKBZ+wJqIyIwqSoH1XXYV1mYE68o7LM+Et8DGW6JZVIJoZ/+kqzW4Bbap1J3WSbp96UcXbgc05Z
VzZHLAfo3YeS1x6KxOAz3iMaH7O4sAYQHjSRiZzOOs9C1UUxDygQYZ6ufGM55Q/0FphxfvW3CFIf
vlC7LBJiye721V4u9dOsxGx7/V9BkPTaDk2KXWhsxDFvm0P2IsRav6I22tksSlM2iWo2/qWM/cSu
KJ+HPdhdfj1OMqfu+fDXd1JpbR4Z392zYs9WUy+C6qPl214GDr1JMmHInoo9sLx9kuRhM97Dcpok
X4okDlLiMltJJC5vDyWkBkal28/wEcvlgzVUs/u0Zeq07WsWeHyD3plU803ZwEDWiLXXBuduhKIJ
XqN2ec1H94izG4cRVA7imAnjirlZzEBEDHBazfWsPifR+b2YHEayitW0ktqGLShpab5y7qEQSw10
OVKjYW40G8aE8lB++TyoAAD/dgSotGyu+RAz4g8BD+KB4wD6eEkonuLabxfWh1BvRgrj54yr7HO0
yqT7IvGSPjuLIychiEnXNgpmtxK8nxtEi2bVkhMUL5Dej+i/XJOsOwoqFKrbFOLb2vGKjOfBShTq
wyreObOcbChQRLEW9hSNLMFdqxN2yHigT32eytYeuE3HgD+0Gi9UNQtm1pc8mChWqETGheVcvmHP
p1IUELVYM2MqlrXf/L1LaM+K/tszscXr3Uq+2NpJ2SsBlLMW6hNnoABal2+lUbZHP7ELGkV6IzkJ
L7g5E701AThEjXuq8hNBNRkoi6o+rkTKFATaDH7WNB+PyY6EhXFWyz8JnMLdqJ4K79cGHu/SyQtB
YeQdEtEnELRZBjwH4VK/P4kloPz2XB+rTmm/VfxO5Z3j28I1gtI4Jk6Vi0ugcBWZA2cMWSIOqEup
BGtMppCepRlgzLu+VddlB5r0pzIR6g5snrf1caMUH0cpIp75POCFIf+i94dxfDhFz3BSqb9lyY7D
9yC02bX6GAdieJUPCcOwRTS4PR6br3DjfXhgALp6CSS8wBJlX8gIn7FNDziDSx8Hem3vKEvyjjwG
hGhEhzGLIBHso7CtwwGPiTHtZiAnM27nv49oHAm0RURRpAOxnZRctKkDMjC7rJD+ewqp4Zbqr3M/
m9LhpT8xav3GnLVq5PcpNWllWHET1ITUGjoto2iKEdtOWboXM67fjLWMoed68SfyhpJJkLq7/mP4
cKmvUXxfYxHA8UO3mSdDGWGxxXqk17SlS5YxOSv6kXeqDExOG8BPrifKFkhXod5a78WkiXLzfvFc
GFILog0tlMul+qRkVkuYdRKq01XKIWbvTXlps8fAlGHUPDTNEp4ifINqAuQWBWRjX+oNUzaQOJrp
usglo7nFCjgH2R8mkWF9iFPBBs2ZDnJwNt49ZFN9Q0n/Vqh6Ly+460e5BnNPmTWklZb0P+aGjAsJ
DAagIgmZDe/p7KlgnHGxOR0bqniZ2TKZ5pOt18COKSsE8lk+eDcjAjSZd+pc/CjSaXbgi9gRmg85
C5tB3QdlZooNxSEhOI81OQGQONVQNkQNTHpVSwvmJUR85FjvWTG8eC1Q3/eW6asMYqi4Anrt7X5y
qmWPTogpDfYrj4hu4Kk0jZKdRFS2TtTUzQ3Zwzw/th7u+B+ToYKaidouxXwjv3ORPSXDDsMjAylK
UOFhUV9EPn5feqGpDhEXUoX9DLmCZ2FWCqXv9R0our0MvhGdHhjFXwjADXosUsllxehaIPeIt3Zx
GZFBxIU0ovgTowinO5+UEzlBI2yamq5Pc1Ker2YyMsWBoXc8cLszl7itVOPXs22+dmHMj8Zm7jZR
mwMjR+luRV3WIMmWR2/ZICVxbn0EeCKTblgxK3wJFwwOy5EoMUsQFJYNvzii9p/eagisKmTIHZQ6
TfXDAa5dUBdsUjKlzwGFfDtX1gCw/3eme4VMhCkm1LyDxvdDDhh/hDGdjsf/xqMoBY04FSFisV8D
dYGw1L/BaaSowKm1dWg1P7PQnk/lHGaDGq63BqB12dwaVarU30a1FAWlntqFup2MBdTc1trJhYfY
D06ACwFBeTLZ+PlWVQ28NgUx/DyLMaprzljLTcl6q0eTi+cTQLxE6cjGiw+FPGmp31zaUdqLip9c
2RQETHwln8TX9CSTCYRe6rCi5ntAZYUVMZm4fwfoFZ4DCmBXTtgE/Cd+EL5TZ4DCULOC8169RC4D
LXjrTSLd006J6KKx18lnqOByTyYEhakv4nIGX4e3kB/tLlRlodKC5LX6XRVfKQ8lfS97qOYeflER
LrgiWx0y+hX0AIRyqhRaknfkOAwxzB5DO7GuilJveluApAqHvTbdeAMIdM9vCHkzRXgObG0rzrQ1
5U+mqZ200LzhesS9/5ni+K2jVjCNBYbcwJ16ieR2iUdg6LlHZdVMxsKh+kYy9bALYP2R0XBg8qQO
a9uoAQr419nMmhYZ/nqm0JMiH9JGBmnoRckyyFdrvju5DasRKkD144W2dw75GfuqBoj48KWukaRp
UZYvxHR5VnATz6mb2PCs6qoum0ceUvRyCFESw7nnh7lnAdvp63qBflhiAqWU5QIG0cc+ZN97lkzc
Am9bk4355beQSp2+r7/R+cYB+lkCnuz6AturCUKmHsaRnyxykdB7L9e5w4VjGvAfKnuxSCEvl7yj
UrSEOBDuOzezPBQjyHfTJEJNEUWH/KiOmMO3tNrOHy3AwUqcIOw54nK/Ox/tptc5f+gyqhyKnP9x
D3fXcImLTGGpse3laFPq/VS/rJTqQom3loIe1kaFLEmX4h+rUy13tQJE5jLWpfA3SdjhxtUZmZ4E
TeTErL08BmVkxtSpVWhPx5dxaLEunVMLtwxeVnfwJMvhigODS0uiuqW01tWV8iFc9P9COTQLWe1v
sA67QsQE+p23acdJfUIHH53v0eDZc3w1ru7crg1k5mFM/CygCPl4fCZGtXJxIp5fW+vi2M+O6HPw
emqDqa+8QyyoGhdwiHpPR+EuWsMPw6/ZbO03BCppHYLEURvXJIZFOmIgdLkl1M6phonOiLTt6x20
HMLC1XPOnMCh/BbF5ocgzHEacdLSW8eCoZkzm1OEFh4MAl1av7Cp64SxsaBt95pranzlV5D7k89l
z0qh/xFNs0J3BBD16m/P4w6BYtNXOP0fzXdwNk0RHMLO+2y/G07h/DiB0D/tELRd7I9sNFxMs/U+
Dqo2kOTCRR27gRSjyqEVUvd1FLxLskwuhsdTn6xqsiQ+KEdE1/h+uzgD2yRC5XhGokL2bA3jU6wQ
JMJSFZnQ4lnA8/q+gEcAwaFhKQX+UkKshJrAsnXD/0isX3Sfalkz5cmw+PKkLpQlsgjp7b+Iv3Ig
pwSZEsubKOOxLgEhN0Jc2WRMuxYFJtD4Xkyi38INFEupbbh+QwPafo4Uwka4RJdJR/dffZblxc+x
k4K3RsdIkJagR6RQGoUzEpJPEmvEw0v+b28qSOdiDklXms3uO90UCBosSuInzX4iJVkbddgYH7So
G21kUKtT7qRxVH77uHHkQlxTDmjuL9FDX6lCfaQYsTJWMWb2UzOT7TAIKAtXVh3bTdnIvsb21VNy
TpRhPmOph0QKq+UAXHidXdoNa2NVl7WMLfle/3THnIcP6t1c3EAyPyBUMMPhI4PNNtwTgijRulzp
LnD7a23BRx4jpxlQroR7DamBQ7Md2hEkyKfXiKjKeqyj3RrsAvB8rt1Xnh4rafmKo7D93IfsCiz7
S1gHwTuwY/nurIDJTK460EJbi+IRNxvcdP6inJ4UiQAOtLNB0Tx21pNpWA5XdBWmyfV2OE0y3oIJ
RW7AiOfjDUrnrfGoKdrPmwh9sWRiNpFOlhC02VSDQqRzqY8mRPEp/slUTKKc1A7BfIy1C3yhqneL
Aj7cQTs7QZg/9Zh1EdiGVDGSjSVzmrqA/rw+/0lUFP5Erhc5LNZ13Ns1Q3xw2ZC0S//uDBuy8CGA
FSgVF0gFr37/Q/COgBA0V7p5RQSavAZ3J8k56avdiTDurvYtTh+XGuffOc5ryycQUkLSHADhQ5JC
zo6RoocJaXoHNVf2qiSyB3NUCexbAIFZ4zbqF0Ch4CV2QTTz0X0VUNOooYY45N16l2lyMgQhOs5d
ox+2Io33DCncaby63IBmJAp2DiV5gSVsny5MdVGClePiWNrw+w42s7rpN3p86Xdrrrfvt8qiltY4
j9s5+r7Hbbi1fTjrSk4If3oa5OQ8LX1KKyQsjZEn8OsmEEnDOmQh2WbP7EVMXGBxTaslmeEcRXCU
VBk1r5y9siCZAshUVjZh9Y/fW7hFaQyU3ars+y/8qPf67ngJPBWU5hhkTHFKjx+wsKD3qhdrTD8V
fKi4uZrlymDsGbp2EZ0OFasMw9B/xMZDfu5itPwPjOKeasoJNxlTPdtTw7exoVKFDresAgC9UPHK
bhk2xnkKxBKWNUEuQz5f7NStRVIJ+Mvr1Oiv2FbEglvd3c+ednDVsMiqIC73dRPboHmJ+hgDkM/0
9SKIncuGyFTnrdt5I36FIUwUVrtQBgSCm22ZMd9iuAWmHXvN2qaz4tNTHtUMHPtFVVMx/z/ilVpk
dTtlUByXFjIRci8BwrorB8QIaS2oGZyJ6mDxn8tXs4ZGs+NkMUFVdkrTavespC8Wd9tk1aNeYFeO
7NvRHeTsvcCBR74sGlWLzVXFCgpD0u/kCE7A71x6HVBGp2l4lEWU75RntqvV4+nBdiPrizmvoh+V
joLKkpsLjmr8mKGSrkN3XoqH1uW8KQm3tfsPnVH+IuT8A2ISuuMdLWMaYF7ECXSRm1rfto0aRqNl
IGByWpuHUoLzRm2P+wvisQ1NjYNsGqD5vvD3jf+ftNLW6fZ2sbxuxMoE4n00wWnY+aem+8Yze8/Z
j7y+6XDm0v8LI46asdhzIDe7INyjmy/zqMiVwoAgKCmKugaaXIRJvSANUoLOeK/ROPO0UMgUONYV
3IrXBswAQ7+rj/aNoVz49JkNc1xOiBGAfwOrQ1PsZjACxFqKNvckNl76oPxBYVCNQ6Ku+3v7L19t
cOTIgcgUFYO6uwI0ZxUHUnsCAvjUCAR8qnuZKbgBZNhxIcmM8GBZIXDLGNa7GHpB5jZRPnihJ+z4
11lHzZzXRQd1ojJPFlsov3DyCm6yuxF01F/Hf7rAuG36pMFWmqn4CQeb9PbeY5sBEdQNAA5GuqMW
xapz7EmIwFLBr6Ao0XNKpCHFGhY77QOxRnuAtu6qn9P8RJ9A2s9NZRyl5uwqdxcq2X5Lxh3KBSQA
lPGHfQjuMMiQ24wZLBgL4NPdliIOzO9ywcp3PksCERXOI6DMJDqwvNTmLe/Dfxi04ImF+W+3s/1s
w2u2fo9Mi3SYXPcA/ZGnLH4NetY+qJrCfXaE76Rb8UYVFDRDkuzjqxlqxJ+RRubX2lIi9ZrD1CbY
FPuWgu7nNC3v2481r6YX72NFFTPFsPPYxzSIB7NQucOQLk7S+2X0vA2T36geafMGuUbXoqoLXz9f
mPWYYRIjxAQuE43twEkzddLfIWxpFlMKQdZvCrAGQX0qnC5+O9AAZM++7VsXsgUXfojjep6JcjPk
GPBmMJSb47HeNjpNWfysMrURcjvo06IdZQxMfxy4mrkOM1QDDaNSxMAI6G/Ts/cedijGhqldU8LS
iVcG/kSa2R3orlsv5HLtMGYHsXPKwUPuPUBv566qdTlpvlcxymS04wul4chcLtC3+7bVTZVdsdYv
XfyXFoK4TFsCGJdSHWYS4/7Ze3q4hotHV+dk5mCc69oy7IM2bRlYY9/otTZIfPGMrPd3KsSIQP4I
oCJkGjJKg1h60/N8hfSKlZClpkDd42NSg9xK9r+YkLtW5YrxscF2jIjdKw3Wl6Yz12Vh0iQt78B0
g93Go53NouPhfALTke5895sktsSuJFPQblJxZYO8vpDPSbYOLmWsK9Va7n4UA9GBzCURz/XyMoF4
AekIA1D9V9KjkNEfpBlO1ZOZAMvsYoW/nEJofOAin5z3fdvDmzQSHRm16IwzdLd1xnKpQKWNDE9H
qmzpovhLJC85DEhi6DiGFS8XOjkM+nEqpnI/7DtGKbn2pDyWb6NfeaSYa4wlsDrrBzKAb/Z2SZu0
YepmKFl1J/lGqLg0e1rJl4B2pVNNdpyDSrrPFJrX7qGXOmKsAiy3Wp5SJh3suFlHElZ+gABuC2ex
TpBoFBNmSGJbTn+WrOW1+Nt8avSMXdK3CjXIjpTvIpqildO0FX0ImeiiJxkEYJrA0yB7SXQLOnNu
tP6LvdBs2WjISrfi1DJQlQDOurQhzrn7DAfegC09z+sXsHUQ2k2LcSOLoECWqB/8BeDYxs1MxPeu
ClIydZy1jH8y9d9RG7PNkrRFMxNm81StLVQmyVxlYD7i+NEMkR9MFlCX7kGn5EtjyqUVZnhdg1+i
CGvEuAKaejXQZTcm/7f+MAy09opzFOo3R+127igLvo9rrgzA9ZiYiSOBdqsL9j5dOiaXCXtsphIm
vgLUWF5NN/ukWvtq0eDuelFKw+tJLRK0m8KflC/6SgnSusj79cC8r+3kHRTW8VQp1ChpDAXlmm3F
J/b1PRSoDK/P7iWuLMznhxzVRB34vFbGI0JxJSbo1x9WmNGuaDhIwcWNWIQnr3gvbLB0e7mvwqfg
ca+9RPp2OyOq5EPi+KcFfZQM2hWpSiN54wOnyQkgERbJww051L0xG4/8ROqkTsvGzUSe668cQIHV
Ka5AgfA9CRXLdmkU8yezNWtq1C0Tpbtr67V7LzmCnuRoqxhFbEixc67Agkw8oy5Zln1osDHuyjKb
tqxLkXSsIVwTVDvp+kPCvebS4J6ikjHC8xqHVGvNj3ndUT7+zBmP1OgFjIorFOmovazFjpW75FAx
OKdlEnTkI6QsQ4xMFgGTcM2oLDIkaIz5NixUHwncP73BBdEFIiLQGili0nvcL4gYxsunR+9yozGN
95hXNGpPs01NYitC/BpZO3ZJT9Dvrybui0/Wae1UC+bU2zoSwmToG3R8g+Qg+sUP0hjhlVbyfC3s
Nh6bLvrroJDN4qh9MXJTz+N6CVDpgEPp0aMDbkXiFzxHQggbxfD7lBJQPRt7nXRfunK6CTl2sZbd
u3Uo5gnIzMAz9apYwqIyFPc2uxaIVIDO1XeI6iSOXfnTDqPhLyQuDu5Mjoq5ViIcvUtgyCe6mDrP
shey8Hx9MEPKjGUYLPMQ2EIG8pOiA/0Dydy511xaMlSh5gOMwPNu9VTUU4faQXyi/U0pr5AHb9d6
a2GZv9LG0OQKxDFXuOCyZyC1AAqzQ7QVMz+lseNC4uR7ddoC0guh4IobOZgenSqfKLscW8Ybo7+o
H7Y1pZyZmX48UW3RT+gMptYDKC1Q+szUQYEhgKVRqgEt87WvQW48gMzrSyS/L2W7aSkdx5+dFP+b
O/L1yefCBiWDpv/hVhvRyJnIP+oFlNQjKHCvTQq//aXSs523FxXgos2wzeq7T2Hq4Raku7CoeIZt
gSmntwIYtM5WrOkOj0aEAYLbGKKMifwc/9BxOJ6ZNjNA2uGe4g3eC5BeGQbqGvpMBD7TIa59NFjB
7PSNAGTJLDgVc0JJb2WDJAUuJKGShIeRrMD35/45HBeDEDMjgD/mJNWySIDPh+6THcHlZNOFvQcv
JOGACCMdBvENyj9ejVOqx4szbV0aF1V/Zm2OBgOUBe2B4cS4RIzyYQG5OBvdam3OyIlfnrHhaAZ0
v37kGPDe5x6EawUvZwRmxEbv/1xwPXamwckDMAwFS/uTEVS/y7pSaucLtl8+lsbTUP3juwq6tHcZ
dXS7qNBybqV613Sx8zPxqNqe7C5CGrOsoxZ10S1nWIJN+BLdD7d013LxMUwduKnyizuVHtdJuwPu
RL0Dm/X5amXcpVMPAJz4Wo/+56wj9HI6WV5+NLOOuuSpMjrmPrwe9bKxR4/PKnd4DUDlbwhAsqub
0tT+UNpy3JoOUCF5AlBOBXPCXjv7gIF3b8WROLIyhuHjgunaBm3W90+cf2UjlPPTRvMwivaDY4d0
ZVPsdJC37hbzmk3FsnpDs8VQE3E2LOrwabr8PzQRd4gsqwBYqJsOsmDiyvnv4gZEPugawNNk5arw
yqUX3gRb29US5XhmpBRG6ZSCED28CkKPESSO1VWTCwZrgR/4WavEvEa9prZbW9BwbhjkopCZkWFT
7YY3womLLtOYyomtmXBFLXX9AN+2bPDlS3hqhyQOFD2RXIwzNZL+vhbUqDdtq3Txmufl7ew9+Ohk
9nsZqW5JG4oOckwYH6CUbX0TaLZVmJDLYjvta+8rYslXwlw5S/JCEqD1guEcinLGcgsmX4CJpLLg
eBLivwFNvEmj3v+oPLT8KWOk7dWJZX3nC5ycGWoGWQftVTSWBz3ZlPV035crw8l3IsMfONiFN+Fq
v3fi7H3DCslTQ0cxE8s+RMClCW+u8Vpp0htcDEGtRfeOUov1xFZChP5TwpqZkX8ht/LbFBHT0u4I
6p/Y9Won3poHogbYV9NEEzPtPPLaS80G4zZy4F2xRUHc8mt+vrlUKaftFINksXMWaC1PUqP+1icC
tByklOp2pdwFhUYAMpfQc27iigBYlTt7tmRs92CjpRSJg0IFdkmFjLIwekuo5A3SbxGPdGFCHpnp
J5KIEJvWWSzbQOeY1cyB/So7ShnG8E788qGV/0nYS7Jghd/CbMsQm57vZIflAnHu6XhNb4mz/qt1
0bz8/v2Za5Sr/PmC2RZz2hjzQMKNHsPAsaq+K7LseSFmDzrxrsJ6gut8N6sdcDgl/MDZo0Ane+va
4zExnam9DCKdVbm3RKP5DA9eh68Lmn1HOU78nyiGi7vNEYzDWy1F0H+/0HfDN43QvkXI5we6beeP
h5Ss5l5VZ1kuiG8aEV8YuqxUJgVDzFZPM7hX8PzOP0Iy6+a+0vzfIfeonigZrpOs9bPzcQ+WQzfT
vzcA1I57PwaxyHOwZLYDQvPWB/9ZUWM2T7gf4y+fPaYjN5Q/wp9aZ8gBAsGmvnaCxIV3fuOyDODT
nFQHkbpePzdxBOq0FDXu06wZ3hG3HtsVOLUgv65+5Glz1IZiiBkv8Y2Rom3wmrD65qxfpkvIutZX
peiJlEJ7yNmt21haYFid74mWzhR+ZTfDWjV1nsEwfdUkuP38+e2wpmbAFpOXr+FBtqkcb79wKi3E
ZGowmWpNwtT00ZcHTjQ46iEuIfK+W4aaUTbNMSnZnWIiBt3jcllf76XpOxAExw2eqY4/UGDdyj0y
e7zxaIKrr7/qAMfv0rwnI2ksyblkVAVj96XnS5WGYtBJPN8oTVwt1hjKiLocJhAf5W+Bz7os9tY5
Juk+ss+lN138/g4uxjj7bGBgO0IyVsZRIM03K8nlF7EwaGnlrwsT8TwukygQ6f9Aut6xCnrQbpYC
Wz98trmwTRihYBM2ktle3wvOlWEbcJjkBezllxH46e1dseUtWF+TfgE4N49gbebJu9FyLZdQMkhX
qz1JP79qgI76CpuQjLjmmhqwykHAUR/IkjBQ4UMbt+1RY7iOekTPmvSz2ZX+/w2e3fdyGD2V2rIP
bFIMRYxUWyd669ZGvmbeGV2JJ8kzEwG1+Fl4fI+JLDdRFRQdKDR6Ik0bfYQe0c3ybXxOxeOfXgqO
lF2vMncsf+AQlh1VMzVVv6xIkBMMYj41bA40PGkjxKVh4MIobc01hS9HSLztHcghqm3VO+HixyQ6
CQJDSfFa9CmjwD1CykcEKFi3KpD7TbWyCdGwiU9/qpzTysIzIAo9Qx8EcGxS9iHf0G4KNQUE6hJ0
lQQ8yRpd3n3ZH/05NX69S+30gfGXm693m1jklZ+mOcxPM8GK9Hn/yj7MaS3orAWZ4v8oCBjFi77Z
9QWBWqJ6ZHGm99MIMeKy5IG4vCU8jnBBD5dpVtMKGKzDCj/nNSNy5eIcGpLMclnBrO/331qVyxlN
D3J36FShKJztggEPYpnuWvVPb10LyivduE/Aw5Opv68YgJzlZ8L48KWEkfIYl+VOg5eVk6vdBOfh
tJbkn+NmJLmqGiaypqRr25UtRCkQGCCnbyf7YAxG3XkuG+m+1ZPdSLr4wD3CLuSdcj/9FUye77jV
UoVvIzAZ7mjLhFUKNbCmAsmXCGsNPoD8MmIVFH7q9I4q1fmxEAP8C8rsDbh//yLjBByyHqfgNcWO
4H6PSjl2etqdWphQobmnSTcD6wo4xKV1GUCn/6JKauPz0G0HqRFwoiCc77fvCDyGpgJbu9cElhS/
cU8OmfffKqDxsgvqFaE1NujcwbeuZBLN94jTCZtElpqNCL1VQ/4FmK6Pe9ra8ExhnO0LPqv3ml8R
VlKjBHfCHeR6WTchAlMFtNb/8aXbtaCOki3eEmOvNBeecS8P9fSy117FB2E6LLW6VIQvWyip7pIy
ScVZIuKcMsisO5Xgq/zwGQOZ140mP7EFif7K2xAS/hXGZ6IhXR5ltvBKdfIrjCMcKqESvpo44g94
n06/tDrI0gQYqJ7GlsY7kAeQUtQakWJ2ELy8JJ1lS857yv5c5bXq9IGBuOvTo/iGL1WBGo+crBFN
TEdfK0sBVXfVIOFwanvfyrGcOeK+6LSmuh4ccdXqkRL9KufTLKe1Q2Z3y/fRy5Epc/mLaxzNfHmb
Tdx6ch5QQ+W7E7iIyvNoHDTFRDNqqPnuBJJKA5BaJ/qSBDVxilKUpw0yrXD5McsqDTiG6BAHU6xN
u4i9kLrJjh9VS3k7O2b9MSUx98nBomgO4wGlVxoUoW7520ZD8ExUfS2F1qIWIKmm8yjrJz+mQ/0D
W1sBGnIomd+AyDyARioWOahfP23zZ1TPMSxh13L7C/f/AtyuoOMewq54yh9NvZ4fXt2MNSEfBF6V
3UI5djFgs/mM1MDqq8P7HU4cJTrbBKsXEfqF50UeT8vCFqrf5ZC+2zUIGK13xnafIEiJ4BRI4NkW
CFAPYtycev+A63zdSY8XFMMyntLEnI4cXf6+1vkrX5e4sAI8iatBmx4mt9ngtSmUuGrp/tu6k/iN
sHnha3rHOUEs2ADgeAJm9I69fQsmjbtFqRvP6JR/WuxvzREJTVescX1nb4JJg/wQi0QKYDqf2dq5
aY5jiIfBDOX58ANFW5GXClSFfR8J1Yge8cVbE7ySGY6uN4XWtS64COghf+xqP04uyvOzTj1c4QR1
4gJ9sfl2kmU6PFaZHZilAWQXaC0lW0eXn44kq/1vVYekxJvj7J+/QROwc5RxqKRBIrp0hOwrb7eN
QJYasHScWw+fT1teCQm5gKUvUSsMFTVlZdfqWKg9W7p8PO2mpySKiQrC8FRYdbgOARHRAfFW3Trf
XC3G4t3xSF+45mACyrntivWEyV2djdqyC5OpiTlHnZyKJzk1AbkRdZ4P6l/Fp725q+PpXTOiQEUM
npcKhBPtJAnAJcWfvgLsWYD20/KWlswA4N3n+/lZx1+eULe9gdATq5pA2atJ00+z7ggiLxRjvFJ7
t5UOlbV2Vyq8+YLE9Ky2Qb+TjXQne8+wvgjEMOFIE0LZFD5+gC7FkOuU4vktnZWHca6dXHpPwft2
DzVbSP91Tu+MicSB4poY5lciEmEsTTuQX6jPVDOYjm6UCTWluMTzpeop4CZ1dTlz8/rwOR/6ST0K
0rTVNo/6fL1aDVDn/syOrEka80Uyq7jRnVRZmE7SdCNr3gpWTYYvIFupvUVUYCLPc7F1i/Wuv/Rc
n7qqcur0qI70qqZEt/v2jJ+86tsL7vzIUWz9rgNddBDQKVaBRaKne4N/ENp2lJ7Fnwq1m7QacUUO
Nz0M/Zlwy8GFj6xfyc7pBSDxXSl+gUpQCRwfq3Uv8x1d8MLzpVcklOn3IkJVJiQjjqFxm6HZ+U2H
IDp1JQmwH2IOzugMO6HiCrriuAJoGgopx9PogMK1yAoxyi4O+7yFUi1ssgi3uOV8tTmGkqB+pMhp
yHy0wN12FHfJadaBFied++YbWL4cgfdLedIMJWxnT1kWPUb3MGw+iGdm5pa+mEg69w5gkOFsFtYO
xPXGDC2Ykz9Mb4gaPwFYsz5qGW5eN71zu81VVow9wiWg247N58uWnlRbD34/QkgKyTr//ktVPmws
sB2QL4hGUUfie99YlemF9HP2PYBF0TFL7cXyLHpVJnMrxEbuaBRImUQAZVdZcjO6Rsk9ugnvbNEb
eArKUNwkR5RlRw73+xIfu05jqAsVwVfKvL0wPvCJSlKKj8tkcvqg7bdUyMx/huzgsOW7v9zmf2vz
7EDWgf9VUo+WJxXsZSvxlafnGCkNUKaTLJfYAqvYc/uqEYs4YzPNGaNuhvLUBfpSil8o6/TFtLjz
LcnfaxLWIy4zhQ4Uf+3wffynkbIW3sj5OWhLxrX7cN9/yFlALaNgpaPvNu2z+3kSepRix/3BU+FO
oj8yEiERTNjGd0cOLNKLKpa9IjZsjZ3cGyKrwpf0m8SjwqiT5W46IwtWP7zBqCQFRGQGtPHFkcY9
5rwexipNhMR21fr29i4k01hwWG1tWitEFs69WfhQWCWkJhiNAcu8UXPBtXaH2ujIbLWxyZEbYP4U
3ixtSXkfofS7fYaIllxLpDZawu4+MS1z0+U+toGwzRsTzBYptlEo2TMULObCoOO0w8xU0Z2JbSxx
S1067mdA7FRyrIuZjlQG5N5NlMG5MyRmjk/QTlkauKIyvqiPgMRL6i4wC78TcUMPCj4F9RcGJVmO
MPvuwukh+OyfkQUdCrGYwt8SEokMwChVHSpZBx/fqTcRxSBn+82+jZ1lif6h6KGow525hR3ae8UG
cHm1+1sEhhN2Axam/SxoRXF8py9yV+7NC//nlF0Tbjj16SZ2e5CZfbp5e3J4o6gM8PByPw6J0OjU
TN182nycN/t//sGpauWLW4TJL7CgZR843VZTUdeOke7gCn2B+dsU4yoG9+WNrA5RZamIFm5vzn4l
MLpVW2X796KcU8WW4B8fxESQkNGOnslcHxzN9T15hSQ2EujnS41Y06SadnJPZ1ZZuzSYTGMQqXbF
MQU4EyVZg1cuDKI7JcOJV04ctrs6/7n7itSW3+o/iIhqffNHoW9PcPfQTsVqhPmFRKknTFkr2G7E
e/RRtJ6yrnSYSQS9GoXGlJYUkHUwFaAueXti2ksJE4fB4B+D9fBGE8RnvU04tL2xALc987anyw0w
3WIIoZuDmPMvtikgmtLYBNskUaWxQBOeKS44dqI2Nzh2xbdFsc8ihkQHd0PzWBNc5dGf4y1Axr1L
ix3g9VC8+yDwowWpiHmRx7uKzyH48OHM+v+v/gYSwM61y8AjHhG3H/gm20aEVP6e5KC+ZHfHeSm7
P9QASAccZL9DXpqRtrZmY3Ker0VzsWH/Ct8ax94J+gGYtkcjshlOxeRNdbcZ+oWNEpEG+s4Jnt3p
Qg5YMyOWTjwGDjJtjx7SNe5scjH3jkvFyHnMuOHUHSkUYOQRyziIxUKUAuyviS9+n+moFn2SV2wb
qM9F4DSqO96wZkmXSNado66Y7xR5A7mNaEggNDg+WHdPFagsQ5WxkoDPPmBxJWEPlIsLPVj3rlhh
Ygu6IjI4jrWd/ZG7BEwmXebSSdjv+E0wjE5WY4CLYSkusS2oCRCTz/m9iMQuLYPVgyOwVcZ4NINj
eS0TN082863ynpeZwK8O5/pMcKsDWxWgrQW1rw769h4g4dRMBLOizak4L1oKfhyJ8sPLE2a3U712
8VGsEJYjyJQgSNhH5IHbscQGGEg8j/RLZQXIN4ZnZKCh31BGETDG1S5r2/nVBcYwhiBxJ7zE2hFw
ZFthuunlq8lHFJFE1QsvN/a946l9ytM4cJQ3QG/4lkRtisZAbQP4DwM1OpVMCBZobVBU9N8/juzx
vZdWpfejjuRD3tEDpkybcRWZQdju7kgu5ViF8RranuLnT6fAgDI96754M/qIlX0Omi33omqSfGsf
xKJCUNCmFzZqQqvbYg99vr/Y7yquPt347lhCQLPbsj80eDggZsfjzVEqhjLKVzC5oUmhuFFEieaG
FJMB0GnWQ76rYv+ZIdY9CnKvJ7gIcB5UsRIYuA8ocyt31Z1jfg/OKYArxatyfzO8yD57NIho4UoC
3SaChI/OE/BcI+K46uU2Gpa0JbX4SNUSkOBCN6ZLUGHKWdo5VldEz4t25cep65idqtTv8tuIpUxK
1AsHfil/zT3J0UycgIvpMdcqK/UeB0AbOBFen/GrYbn9yIG30wez0IK3HIw2njJYhzDDVn9NzcjN
MYGyMHWwW6BgK4EkYAJ2mUtHuuXExJ7MKsh6lVUymIqef+EvMNtMNwVm+1zBNrRxdOHzzvRBW6ly
h7v63LFUQDGUVQsKHQMDQMQcz2ZQExn9/hqySt21irKrx8Jj6EpkpVazcf5Y5ph1IDgrUXulPEVq
TbbwPYdV9LxRvrkrltG+6/657e/LbXaWA4lTaSXxrAZzy/29YbnKeTXEXninQFBTZjUUERlsLiwC
3AeFKAaBKuRt8HViaJh+VlLjXCr18sEcx22xSDjHmoepTkEo9SjM2I+6Ac617eRkXTY+xH4XLth1
8AUBEzEklcXVVNh5uxJlTXPY2SJgCLFjZ1ttNh1dLyFKiZdX7BJkk6O4pJSF85a05I3h1u0lzx/L
WIiK3hhLr2H1ID2YmBRP5ICFklkqfEsQlgXpIcZ9mbXXRmBXyiy1NqOk9W6jZ50sjAEGFN7Ax8NP
dlBvqJET6beMUGGPE758G9uDzKA8fXhCN+wcrGagJZYzpCaBCuNhmrgsxzArE4xp/YVEBFZTvBbV
7dY888asJRIZ5/fDRC1j5aEdQsp1RrfhRYknwyTdAkUUL14wayfk+nYrlQW4lbHArwOFV9S+aa7k
rLVarF3VuaSFFZ4cHKwrg/Y8YHDLa1tymPKnjUhN9mL9Hbg+EaMilf6O/dhqNxT1/DHry4oXlWND
pxE+l+19aBRwq4OW0waXmMI5CWQk+kQng4Nz0yv5NgSnc91RYMevCmIV3X5/D20Ke8fyCTxHtVNN
cg4TLyaO5AzZFOnjkALN6JNEmlQ0w86ySq0EXUA1HJa/TcWuclJ+mPoxfROvxhn93aVxMzUAcf2P
qL7OCAgfl9/2oTUWOv1R11vMUCVNocF+caLYeRT8AkXEhO7uD9u+WAa4ZbzTsMe1D8rjriQGyZ9i
ARFjvnM2zP0LTH5UyEYkaGDzqDjVZ14ZpXYQ3+qWHF4M1P5sxGVRSLNfIn0bFy64+TglncMNOw0g
V7KJ1KSHuzQ4gd5OfLXRn95PqRKrIZCUmkdSeJp1N1184crs+LVhIN61apKpMi6guhpOzdqGY1Le
S1d9EyL/aAyupgVbFY3E1o7jfMZ93qJU+lhrYD+jjnB27JPmg67jQkA8kIQY2ly7+fSTeiop7Ssm
9XHZpHK/cDxEEJ8RKqRG/0lDok+vsv7c2Shg89rDyyHMErFuC54wd6lsvP5jexjHFxq/Nh3DQOm/
soUcyg0g3i/NtSS7hZk4yhRbM4B1C66sspG5setmSqq1Fr7oWTiSxHxd5FZKDzOjBFzNi73BmKmN
InifYGGWzsi9gfUpWn64HYKXig0e8rZ73XB14k5sOx04NSrBkzTI2t0OkSewcJxzUF/CHRPlibmR
1/9ZyboSRCxN6bAUBpBd8HA2dvEchZluI8YrkvBdHYn7KUYjEM5DnDZxFJbRJnAFxVroIMOJpH+O
Kfce7hLp0k7DPgI6yL4JN11HsYbHcJk0qYcxnRsYje7u21YJEpMZUnpLKCvh9oefWOGY51bsIYcw
EEmhiXlrtzH91A0+S8uNP+uy6550px0VqlbF7UNz+VUxDZKgRm7M9wi8ZNeihy12eq7G5b75m7xr
mT1dMKPc6i3MygsFwdVWMWSPoIku2IxGzkvZx0IWA92lHvSNpWlOUdjNjxwZsk33DkVYqI44d61b
Jb4K8cfyjBiTDEFP6isW2m7RfEBhlqZprR/uhVpiV33EuZ9OKVQwqKZK+9/auizeDRLpAcfK2yXc
PbKugvRoydKM1Op3O6skLdol+wCPVqRfnZwbJvcXVExDfCO6ObnKGQEZVqyKvxrE+bXqKBpqXIxE
lxHu79bFpyo08ZoOt02OMebiize8YpZ+jYEMAYAffBkf2UMe4hQFN3qDroDG//zqA+Xo7TRgG5gn
9/M64FFQPMzSvTzQrPe8eMpyQzPFNU6E5auQuwSbkGHfC2zpgTVPQ/S/bODAyld6DeKZTfpidvmN
eSjYEOatGfQ0YPZ83pJG6U959A+05y2E60Hp7ZMFvJvezuBixKxo/V2CHm1Shg/MzC8XzCzelqz8
9MpgTHKrd9TbU9pjohT5F06xKjWRusMcSt/pPuPj0eWiz6lBpE06pDUttZqacYTdrJT+c05IhXAD
283dj9ENm1LDjBJHRlTItClTa/em5ucxjaLeYcBsKzmiPzdrDO0fBXSJ55UOPQS98Iw8iuGR1skl
bAtDoXLnyLZ0KRoKPV6q/FuEmCTXqN13nPsE/a5kbh++3dEd2XLwBfRuVDBVLknTM50xl0oHpW37
kj/5bQ4fqZ+yH+sXtekeJDBX9g6xsZQMKvbULvKR1qbQi7gu91fDPAvlR3Uu+zTxXdAEcAj+RDyj
joTVOzCA6nbkscCWlT08fA6WgnctJ7jFqELOXl9NwmLJvgQ4RGZBULbo5PzRwEIVZ4K07r7Xdo/b
GvDwy5WA05wtunXW5lQGiRwVZUETV5GFnOo6vBUCy4UFG2N5L91H9pkPXzm3uVZfnG/feSAIMxLP
8i6z9nVMUo0q2tA1sRTVQAnIRwinBbvvT024n2xenUqgjwQh94iikwV2baxVVpauzHxJZdWhvOpS
vWYFfnD6QF2s18IAmDfR06WaT1+Graz2eAthkMfaC25QWq/eX44LSGyHkuy3d7TNCONu7g3DuYOO
vbySaGGIeDIy8cE13qohd2USWk2cprlqsjgv3VLOUzVAszRE7q24UltW7z4yHUL58pwJA85d/y8V
sN6n3uIRLg6dI+NtV5yLvtpgYRgJqOpE8B8FcGmEvw0WUFhSV/lZIG6t509maP+EWnfvNt+JCzJO
Yx2uCdCo9yt8ddmtaSpVc43U0bQRPCdGFclmcDNL1cZ5jr4B7WJBXx/7v9Ymb2L/fymQN37FyPxA
+lTaS5tgADx2H5L8U+vkOwYuNpwDZNYQVi1RRA4qm2tq8kCG+S3NaJnwTgXNovmzUnbZDEh/KVIo
yybsu7fy11nlu6FZWkPfZ4kaK9RnxQKFxQwbfBWbNjgrBAx2h9A7u/gG5/s4zsLWZx3Ok9/Zua13
9mkQXc6uDct2bO0c6ZSxHbNmXhhpjNs9KnUZFJl7+v2kARETYZDtLm/GmvHT09ugmgLXWjvfzMcB
429yzlTjgOKQsYH3Tk+cFqqLtQEO5Gln9Iqz7e9+dY6U7+0Gcu5B0IfrYpW8FIoG9ice70tBXQa2
zMSyW3Hy7leyuDNeOvkZ9NNn8D19EKhqHjFzoTd24b1dOuAZebllGznI3gIzB7iR1s2h06Mz+P8u
8a/H0LSFNCX+n2657oVhQ1LxgEpMqUGRa7B7fysytaMeEuktkepw4x6be7H7z8kGzycWfuI452O7
1uHgjVpbJfG1eHU7OmAhEBb+1S2/uOHI94/slszI54M8UHAXoYmxScMtKvL2xYA5kS3JIqhl4Lr5
ue7TLaACfAq4bh0jmLkBQR79oHUSkwez7cEmQ2FshmcFYNWdcW51HZLV6l2tKfbYFmZLY5kbaMke
Mc3Mzn3wKBL5gjRx61VfFOkPuPU61eL2bxuR2Nl4WwXGy8Z64RoIi5YI8y+ONUICayub/VrLwCep
CphsF37MZArY3wbXFqD4zaAFi19t+Q4b3kvel1i6DlK48wATholBISK6PgWuFUPZK3FKcpnyO1cg
e7CZpmrhfrgx57+x+pcjCU52AOmzcdK6quCUuYvN/Jj0CnqLWmfP1AhF/q8vgCirDqEzNTyrELUz
IJ3JzEsayWxBTAz/7/ImGImZURP2x9xSJJUkGf1Qs0KgJ59RP09GnSJ95XM2dIm5DwcJTdumoWdd
w+MlAvnbIXRc1ROnl+5ABuq3hGh0S2fClTz6N8BT2AuLSKCj4Gb3IT8fZMOPCZrNc2k75t3NieFk
gXQ5qUsmxzo7dENt0YSBFfuHCUcnIzvjid5taDyeIJNSK/xgDiJrSu09Bmp0qIuC6Kw0jMNS4h9Z
mwu/5pDopJXrYAa1V/tzXWYYRZm6gjyYnLyB5dUapQ61+koHKKqP9GrH7gIJ4KXfzY37P9dq6JO5
J/vjM2bLKRDxzoHJ7oKb0CxD4CdbImrN+Mjul3pfN7a4BRe4PCaSZ2Vdh5nrNYXjVRIm3tGLn7fs
0fjfaz7C9O332RqIw4MPBkkGt48ImDiSZdMVhLhZOmHV2kXvAG+E/9lWZqamNQQ0FMjEA6if5gBC
HDr8GmmPorniPfHmCa276/+sNr9F9SVH8+iQbbQ+pQ9As2hJZvWWQxl0b/Iwvxa+LJtptkmuVr/Z
A6rIF3aI8nx9c2yq2k6NjGpGYkfPd03G61+P/mZP95cxV0bZGmrn6Hsge3gno7f0BVNWGYa9w2a2
tNCNCeU7Q2fnd0ZjgqJs5ngLTg88MV0dP0WnKkaNjUaiYJVkrKlMYgZBsF3cFJHpXjl53ksW1sli
7YmbZGsU/DFOSZRQfSorQMyNltPGCdw8Ue6deI/4HgHhM/D3+fMTNcclk7Hqyf9ONZkSGayuzBSo
2yff7+QwOG/BHMkqCWEPTBTsXYqEZwKAMQAI/XqDAM/xPZShNFZEUcfsJmju+56jl3QqEPNCCmNs
B8ykgtMEhAYKKqHwrjAHUakjem/oQDAYZjAYeJfgmMY+LNgdF7FzTlGzIS853aoSyRs8HboEBXB1
MMa0CvxXJT5qEAb+YZFEtsfmt3PcDfvKiIaGTV6UIkj9NhdiflDRzZy1hvPLzldVkFfdj7ObI4O1
tMG4YsGVio0sVXbDahlEledK+DSaUxEwi6zcnnxvcYJMg3g7j0LF1pmJgHHYWiIJKy/p7zKqawp0
xb+RDWV1zWBjmiLGyU81yGj88OBXTrK0aiXJLj9C7RCmdye/G4iA7O6ltcpVwZp8YSA/S5lLLM7B
5NV+G/d/IIXtGhwiM6drGEdpMBSnRmXZA/8xLUATYpN4DT45N8Jwkx290XlrqClY8rlMkAOiuOY+
Klu1KjFx8vWICm9mRffrSe1JHu9OQ8wWX7c75Uh8pTao6QFhLv5uYmkoFDPRgR0Wcm6LkBlLBOyj
DhlJ6JGv0nG3jTXn1L/o3fCliH2MyAJo94yh9QGUUnbGBuwgJCCJXCNfqZsm/fqA50s+SFONduuh
yn/SoECRF8ZQtPaoVM+CO/sht7Bj5ALmUoFbha9Rb4T6xmOqMmxS/qxKR6bB9wSoG3u/JT9uG5dJ
iFVBK2Yftdl09IU/wiOHaf299uMrkOc8VJ5DqX1sL/YVr+OGQxUoR8TXm4hcbe6CZsK5hb0GRiXv
td64aOUeUyUixpMRdTskNqnZm2C8SHQGqorddpEmCwIhgxH6/tMdYDHR4QeFcz5y/KhLioc5mA5A
qQvZXhn7MUIIeLbL9CAQ1AfQ3vO75tQGlobmv88gMSrFNrOAslAQp5uDgxf72quyANMvyKZEU4dW
h5FKEgXFnE3ZuyEGJ6L12zEpbn+iM8QoCxXhyeeSSCM1YmzPmFVusbbL5Y9m3DfuAN+HqmMJFT+U
LAalBOTrX8tTOhy6neTALs3QFOsGmq8I3jVgtR2OzZS2UCY7OXqrElj5vnby3d1CXkVoVUCECsAy
Ytk/67qBUlfB3iPyOWC0EH5HA8npaLfXNpq9Xy1TKNKElDihYUwOtoJNiSxPuldQSJxHYDOdtv12
4Q1CiMuVCoEYq5HaAFuUs6AtTwJLgfnikwzMf9x9yQb+5w3643/fNqpuqS+rhm0ps5Ou6wN9JABZ
+Df0u1wq3o6O7obrSMDwyv+ghjI4eALVw4iz0MVTStcY7vJqm0HFuILOrnELcCvPVWCHlw12LRkg
Ea44V0crKdLARk9C5178m2/GtdaoZGd9s+uOvp7JlQ3/pTJoWcOQk8IbL9dCF7OFdMpcAkmDM8eb
Z11Ef8aZ62LI162OeBgxce4ukn4G6oNEYVq+i+0f1qeDOqyMjpsfH1GS3Z8IwCTesHNY6ARp60EB
hK1NsbxRmzHqnVCdsWucvqpfn1e/aCiVJoDXdnM7S0j5NUw7jNd8P3yWfcbtpQ4TWA6MvDYpra7e
dC+696yJ4MaPfBorSonpQ25fxA/3GirCwcgOJXvpLt1pJBayE9awa+7NsQz2qQqQyR+XmVYhqNfB
SXjbT14gw+txdEcelvZRoPmb9erSYHDuKO47foEYNOnQZnQ7wdEUMMCovF2DrHtroHETQk90/UOx
+Lw0RXSy6Yexew8BWRyjGmIGseZqnmg/QspqB3v5DlQEtoJ6ReCNvczG/n0Ehu4bqlb9J2rHYZtw
NOp9/t4Ihly0LiIHPNNFot5XGQBGslUkODhBbGADneZitBEnhInkmLjRGXZjlyYa6LOsn4bJu3FS
anG7q9SZ3gXal9BGMZbQ5pVmGS7Oyu2NpJrN6PajxdMJVib7+9byu/kBbTUUvKqZDQ5sJpXCMmpu
1LITTbmSesHN/pJxa6xdyTaApw5orpCpog5pwuS+P1quhGeC938jp4DHqrbFA5w7IVe/gz0lAGQn
R/uno3hbzNzzttUUAT1NeE44jtxTUXzlvL+0VuyLrsyQJAXZhubU2OgVTiyDV07p/p5B23AFC49B
l9gEYf2RF6jt9np4pZtmmyBHJi4P9m5dExTmoi1FWbahYOP1qr1S9b70Nc/ZRQe/g+LM+m4x7viB
9Z6pmYTp3kcpPPvKDfJKWpi6DSJVVbfpJXEXG3tCgajIbuau33bkkh8FsRFtTAzRJdcu+2+15ziF
IMYdUDe110psXmhuOEFAntnqkITZFs5RDM2JYNfwjhUs6UDHwVWU2jC7oHrw/LJJdXjqunNyjJpz
tGTOtugVfceYsxOu0sNuXKApujugB8jEbPxWA2kRkEHGF4PJaFOGT2qpxOi65OlmThh0H7F7GPvA
b6JDVWOnQXdBI4qbFHLPjRDdHFeNWcliEDcIm7PqjtaJ8m3LH9kDiI/uPnOOxhHKuoHARfIBPh8Y
bNtQms0WQLV09ENipbXaBsKb8GOcHG6k0JeRd3xf51/3dDJ/K3QyMGiuDTH3DNJC0UEPWKAGyXCZ
tSNKahCoYQT5uHatZLHCEWr+jG+2Z+UeIj3kHAPFR3qtBonXnJY4PFSF/l3R5B7MdrYKcYSqRTPe
aeAGs9+zEd6DLBEuGjMlU8jZzlm6dra2rfVvCr7Eqdzvr4ESJpS5tfjcPmn0iSqPPgP12gCIGPgH
JKIpzKnlfzRD/PFnooNZnADeLtThWj2+/tehx4ebsjErwBdAyZUTa086qUhA/JVyKuDzyXurKwLH
1ssDMXUsKA8y4cAnMOWse6MGkVpY6Pbq2gjR6vB6DO5KseKsbINNKpqpDbjUGupo4JoPYealpKHF
XZOQRsFxX8VtdWe1rhJKYp7QolG3XaVqfemR/TU1BYuj05c5YrtoZ2A8iCDao3uilAsTN+SfJeUM
YPYO7AN/Qd8KMlLQCpcsKMonjUyppTXuHEdCkc5LcrTBNOITqIEBEVm3jeC/dD7v49/Felcqsgbe
TEUbSlZ4dGe0+ax4Bsj5Zf142JdM+fX9a8Q7A47UkzdKI9Y7BRV91Ggrq9MMDRA8eY2+mNvVp13Y
cC8vpeMjq2x0znZth8Wx+S+B2phPR7KB5M8qgzHpwk2kuSkxZo3MJN/Cvk9BV4fVMOl58AbNaj+m
Mw5s2rwKC70LmLoopS67u7I131e1NFTrJq8tICFMVvYDdioNcBx+0MomQnNsLElqKwyv5+0KD8sS
oQmWmt3XynpwgS6R8p+znKGn7/MoREtCjdHMpbzclg+TV6Mb5IC4w1Ruhqce5cvriH9Pb6pATkCM
Gw++Cs89jztlz9oqZZgE6LOepJH9x85sKbCN5ad/w4fvA9fuNuUKObVrQw8369aIJVNrSQK4spWo
VbpD1Q9rVB030bA/AYToBHVIvQIAVBiRFB/RWQuZB3FZzxrZ6jvkou8N31vuw+fEYcgUZTvqRscD
wX7bRqdVSz1HOvWLYj/Vp0rJC4HFj4aTIB6F1abkxCpmMhrrtOh8xKk/NGbMvAXAJuoGluO3Dtum
3bG3rMZqQede8yGFQd/4x/nlLrf5del2u/9wlLgljn1V11/+APdKHmFwOS5RgQzNX68bX4E/63Ii
ObWDaok9dqdZ4tgLC8eahqHtXZU9i/QzBWgpYkWxTYOc741Qqt1RFZrdeKpjjpfWQDMeF+suhK4m
0KZ7gftu14044AHu3KO0UNdJOdyphV4Pt7tMKqIwcaZ2sZGE+TZq2Mu1zBhWTW/ziaQNnEDhOh9v
Kstsd+mVsOGxkrOcAlvSuT1waNbRJNYrnjlXvTQY/MxkEIhrsucaRKck5sCjpMAUMhEvhhFzdQHo
lpmGq1RUyA2wyVEATiCuonP9g0uHAceSIqKhqPxshAJEMemfSCOob41ZOjN89JhXaqggpDAddoZH
Zgn2hyJPA6B1RCkWL2YiwoHT7WmrhoULzhVYrWqKAoqBtzdSb0GEI9RO3xpl5rsR6f2r4BtSQUZe
ieGMujsUVBSE5uaSyV8uin4j8dICBHAHYaw/of8Rv/pcs1Sn5At/xpOCVD3AxMnxBXOSgip6fqJL
t6vXabfabmKRjk9pfwwKKkuV1yOvJmep2u8Rfhl7L9d4lFDRkYgboBjEYMBJJktQ3b6dcPLKM932
i+iuksVIB612AVh/ybA1FAcG1MQRlYxe5Zo3Z7H7U6DSHpxLS2CludozrP27qxKPlMYrrp2Fs2BN
nz9S3Yqb/0RauxLZbPKxXmTLTANEqLq+MCFbgpZldZoX1DZi5sRfNN16iMO0BKS9USXsxNZfKtNt
rvk6LFAQf1M+pv9ZD5+2hN/al1e8mNiQ8uKmuHq3Yf76Rn/IqonSpidns6aIN3fK3MjaIRaXT/cu
r+rKO8V642H8s8WeFYcOo/LE9T1kpJ2qlUcbmR44BIy4nKNDc+DJmZrtniuTTxb67/B1PAnqiTCi
PNuARJ9jobpvvzr+Ej8Ppk5/R3bhenWzBFQIX9Igk8yKzR+2qENgmgA2aO6q+IMvLHQiaeRAfZiH
nhh7IOC0jPifKavPBZvJkM5h5k0E6E8GNeSZcFFP/kHA/r9OAM336CWDM1PtCDGmrjh7fLcys00Z
EggfoDkyKENAAKlB4Twq35tI84cpygCGoclA09SXyvv3u6PcBgmZfO4X7rloIs1qth9/4Sj8bUZ4
oKTlRGzvzhVN+CyQE0V9w6BbSRRZmVGGjJR1oMMUeEo/x9pQoNF1pr1luYWhYu1Vkwhg+6aw1ASN
uK/f7bcpTDM+k6iJAos5ew46ZezeAsHRByfe5DOX/VYQc99NY7nynGMaDnCUVYFaIDyTVC+vm/Ag
NaLuOPvrR31BTIdv2SZ2hKazVMX4ct6i0AMZ0tO2YMImOjNX5r5vx9nxwWPvx4ayK6KaWbqSpjLQ
uraVbAokuZl7AipeSprV1rHQ43xUyC60ctSovjAvrhlfWhniyaJoVNeczMEnWCRF8K3eWQWnYMGz
8WIw5EoVfYao7KQarH9K6xG+GaHDynplvCRsBdFqqpB2WeUMXD87ZeOxY3zl8u4ToZa4Ctf7+ABl
DfYySfejzFjF6ed6rKuztveeq3pvTvIwuXzarqAx/QRWkcRHtzrS5Vr3PW95EiJLTRchkyYxEnSK
4tV0odslpzIB/SlOefdeLhJNGXDEUsLGsO9CXTEtawM5Szz6qoYyB9I6hq5sonfali0iaRggEft1
FKtk3bCIWd36+wDQd1PLkaWIor+2ZjrQrFOVsHHa/pB4YlLroKy1ZS/5mN5E9ms+wJtX0Fz0HsIc
0zD93MozSAcOrOBpxVQrBkiRT0VRSV9BY06rtNQ9BbRPmCG9/uh4XHbCfIB2mxEG4GmZJ4+zNIEr
OUzF/FeP1upRP4vwQZYqwJwfyAh8Fcwylhbm1NTKcR+mdF98ssAyuyTmEs3Tu8h3R4Z+STG6p5Xz
Ygs2wKLIbqjqX4YIqxiFRJKq4kAg65PydsU8jzqmu2MFBNQSP/E3Ok3mI5qNl7hQiiFm9UA/vP+E
Tg1Xjp3P9ltDIGrOse78mNfvqCt2sKkSDbHwuvdoGjzkGB2hN8csciXD+8Q9R8AWaDQ5emmqtWi5
W3nq9BLG4YeRlLejynA8+FWs87oBxyzJkAgo/AtvcJJbdGzXAXqrm1guhLi0rQTSfqOdOwga0ELV
FPl6ixP3YqtxTzVtKJlJZqRSbYW3Au+RgMi1t44SgsHkPRDDLuTu/651eBsB0cG7ZrI/IQQpe3gl
izHcz+kUih8gU9uKQhcoO+yhbxWmLcqvrnLqUs/jSDyINoDtb3lBon+HQiQK+vzl0hfrWJXSsRhk
qQgrYI3dkJyZK+n4OZtUCJU39YMVc4JteZbA5QQrNY+ToTh+m5+LQcTwoSpmI/adzEVrfhXuRXoX
vvBDmhedmxo0lsbHs8vVIkoPrTj0KiD78JffjN5I2BH7H6L54LAhHf2nDesf7QmS/u69VjHM3/WI
30LYUD7N3LmsXV+3bmy2XyQBPLumQTDsWJsc3y0TaCBwbdkkk9Jp59lCYI4WzovofrFaz/wwN1Ul
VN8IkOCJTWSiMYBZkird0s14dN48Gok4lkwx6MQ4FX2sTAJg15CORH2wTEof8oMz50AU3p4K450v
w7P9e0Qbgufoivsjr9EimHQtDVsVB+UJ4cm+tqG4dV1ReMsIS5OWzuH8cebuci6aYDMkUycFhhkP
lzMP+nxZkEzkAREta9GnS0ryXv9Q0gf0RmrqP+t8rWfY2pQMxd9u7APYdkz6Xb1k6jo1S3gTr/+g
hBInaV+A67ToAH6nlBzg/YaQWkN275oUBTgp6t2H53Grs30WiwpVGHFp+n0Ar+AcaTduhr4g7DZp
HiOB7mxCcJPCh1HsMatNf0co2CozApzudjx/wvBrdszoaL1yvkRatmVCbd+vrURJkbZCukEYBGHI
hzpISeNdyiXThewNuAOL4NH+eF1LeE67LB2xOfBMrA2Q8mcNHzCeAXrR5lX4Z+a820AAE6fNLAZ2
YrtKagJ4lrvJHPfYrfC3vYD66AbePv/vgLvWbjJibMPxcgeReJx2GlCt1VScURi99+c2IXJKkZ1w
hTMwujo46SPBcyNpd91I02HMEkK5m+A4bn59piIUw7/4Ea0qInf4Ktl8FoEBQrgbsG/lrJlOSqCJ
E5TyXyzZhp7L73FijaVdxQlqRrB4nRFrOCsNNYiqjfwz8zh+VVk1MiKdhzSqMCVjU/IrfzD+sFJw
R+7AYemEDy+4edW11L2DzFvEFetXLWhp/QcfdZ2lDEJ04eUCNSLOJiDN9fw74/HzQ/24fzssv/cQ
9vxqJzkuoWDU7l0xmZrXARpfOWA6p25P2avGj9mp7nbkEXJWfj8UGZfcF35ByI8doMwiI0wQXiCW
W07A05ykHD1TzV4KuqT/RKG7Rs2UsCfY9xzXv7z9ByfZBXUKUTh8MghkGSqBLllNVEBWtbWMO1n+
TOXiqqtbWUZoc8c7+OnpQQrDlgHBNu8AZfbM2edlxbrOn5FZOW4ywzifApg1WUADx9Ce1UIe6HKC
xlQfF1xhuyfdsWnvNeBjVpkVfmNOAuZl8K832/+XOjcKMUfcCTrKGQgyzDbZWaw53r0XYhzYQ5/o
a9Zb8J7vWutUWcxGCOR8xKJrtWWpUkZA7MP4NNJU1rMF8HvTAg7iR1+rWwYvrqhwrNkH3S2sI7NZ
4DoKX8Gq8UwOWHekT9odaCAAFJrQA9y3QgxdUQj4Frj2+WXAvpGakM/gaaQ570Eg6B17o2J0Rh6M
BkZEgmJw7Y/SzWSBmHqLpTezuKfnvusJWre0mYSMBDJPtLvyYABqHZXPm4rQSQS7HHIDcKWPclvh
VBQlX7XxDAOQhDo5/aBVXODZQ+czMu138Y0f4AMu6+7ccLSMvg7erOlQkVrz7Evhs18bOkbqulPg
1kr3EJEOIhqeYIi40zRxkN4EPz1oHI+cOh6ZVh4Yxux/F1SqMdDk8UEMq04p/DUkKseUBBdahTAN
WmwUPoniq88qBK6EFfHgM2Ftr/0vVozSyAsHLA2QvrX4MbG1xqaCOqcsTekw4q9eMv0n/3JGN9cq
mwYV/vnmFTzOvIBsuNq7+zmBq22ilEpL87IxWUtYGeeMxurWbx26ksIJD9ML/oZgGNvV3qzYga/6
Mlvg4A24GlGcJz3WG1dRarXxFm5/C9rmCKuJ951qZNNTkOkTjE9rc9RGyRnJ/d27qBxdOOjbVLoL
li7YoVZ25FnofNwViFAn+aqW2bBD7s8qvqYjmTK6KDqyfuGqDlZC4vejAycnAmssOOKgW0tkf5q3
Hz5hotkO+QyQMBt7OhWBkLFQGgXeMUFzy0R2hmvCsDqoHFJ0ZO20roQu1RAwb1p+SajXOkVoXL+8
hG3/11oVvAHJhaQzTMtcW21HdobjQXKTBS+VFM37TJ7Z8cdhKIrk+Gr918tpgRqFbbuV0g2zGBdx
2fd7V+cqU3S60JWesP9QXbxmcZfn7tQC3/HiD5kBvdPdisTisU5TFwJGr1jNWEv+16K+FuRtAZ6i
DLh3Jnzjz9/Rfgbe7buX0y8v7Rc3cLPn5iKDKfgfnohp+PGLxAbExsnsjPJX93cCB4I0v4FvKuXk
CTiJ4RUcnLcJ1G7OblRDANh5KUDYXBl5u7xY2FugTXGX7TsaIFMK5OtxmDGMFPI55/xlAYx0H/kD
OsQR4VClojB1UJy8e0GBo+bq+E6YnWK3z3b7pZIGu+hPh1gQ5OYwaFWhXA/522nOz0jnsQ2liXgH
2VUY5aNvrDcoaVgIcyrdj4MEMh2Sa7qGYsBozCwo4AI09m5geQgYj77i/i8C3se7V2rCbC5757an
bjETotSvhqYS/R8/Qd3wJ4RucAYFe8tC8wy75rmxBwLzJpmjsmuFHsgTX+UjJtvfOSF7U+2X7dv6
O+92yLzLdgQHn75OfVEU2L71aU6sB3Nt4Y4Vs0qNm2o1XGN1i2S6iif1KqkSDAmg+3zqrkuAhbLq
D7QG/NSYcLRAfQ6P5y7vnhWJd/0BuoIDIXlthVyDeu3nRLKzf7FRhQQCx8rGN/noBPIvInnmkO/v
haeRDmbxtSzWHizwxzoFHIK5ySavsGqEapkLaJGKkYu9iU0VvqGHPZjjAFl4D+hLxDbhy7kPByf1
gKkTFkgbPGOLS2gBKntmygKJrYXy9qXeuVC2aGL2HB28yVmbKPxaGNo3SFI20x/7pGFyj+bi5QKr
EsUq0SWQV08TGdz2D68vmcazBDreNQQTeaa2gsht64MZk0WBrQ7GBqGa+CWZqWQ3L0tBCwx/4rfJ
L2UyIn1LLIZEfokY47sO1eWcWNspJ37JxoSKJZCKBVYrEBnY+9BcjIp8DnWOTKLtPRzoekySTxa3
AWNk+MZvOS01ES//0SzA5mWes53qYXGqIZkH3527WEhIzfxivSu9ZIBkh6uNNVS2d8g8P07rf7Bq
wXfmT8V4u1hhSunfUy9yxERLKyboLJeHmdxzrdsmnhCeG58BDzSzD2Fds+s7+7N46+Lwgs/matMi
WpZS2qrCqKzIpzBN8bT80DN+DoozwrcH3JWFyTs1Fk+ChkBdOHOKfrVngKnOU9bnVbXZ1ZDWyYIk
Mr5iskGaoYGXzKVgRpyP1AKUAl3MOmo8mSkPmzrZsn87KdJjczbSWbtwz31kROlwkcAXTV3BqlEd
5f/1s+70dmvIsyLaHssUMqhGJiPE57aJMWF4K/vJPDffzvY3CBgf97/5IETfNU+zYNvkzhxFqMzS
SnFJLZgULYB97wzL1Z7j3+/w+Tx6gzTenh4twJRsiArDjP7rxNxWyUPTbzOA+C8ihoAh+nM/a284
m0y8fnuWb46jiC9uQPFl85acT2EILlsF6+j0ON1DRbidOdkpOj3VIF/HKtUCOHvrUFoWVU3/T6wZ
TunHAAFiaVb19LzsY5qE5f8jfR/T08nai6rbTewmclM/yiXT+eqVhhLJtVcl/v3cmfOQ9szNO+Xq
kRGLkPmHVKbtimBX8c498jaK/p0IZO4R4SrpPd3zAe8AkjKnrBb3P5IAF0vMLXXJXXbi+g1NkWKz
bhJZpahjToL/VYK4Od0+QSrF58EqFkVjSIUefGMyRviQCfEyK1m1xDRYrf66EIYcJJ5/So8CuUR2
njcX/qTzhsuiz7JFI7rStwXlLBYKP62StRJ20RzqX0IpyeGEiFyqPF5towdGOqOT4TxK5LN7wSP6
qmhDcMwfL+3DOjF2dcNkbYPD0OKyiZuVqWJ2RRS8UFHLMX32bWHnNk39KASQnWSFQSHrIe/h8kqX
7Nu6Kkk0J1hkP5bjjeWoELSpltMrgUygkb73sFXCabJnEikm90R4ogt9jZImqkG3nDB5V6n/OF4z
3ZYtvRA0Z6Kyz8LF85MeuSluPiR8nbzHWDGoZR9ZMmlkfCJfrl27CuV1QF4e4Y1NqbL4ujOpfwKh
+h/zDefw6H3dBtqzWbB3uX+cQ1FFG36KuQLEW5zCJRlibblK+TOBhGc6+3Ui/Hk8J/rINFT+/Kar
jQhnyuEE0Qtc1kef0pFMhFRn5LcPy6Um9EdWfMIJL1ueyXu33Je5UaQ3qwMWwA1FYa6qh//LTLsR
LKogJXnpk0AehG9CKx1sDWCnkSATXNvmaQNMXvqr5oOR8MKmpPBiCs0X5rT0+WACme9T+FSdfB5v
2OuzOEuXgzVgqldcq7Eer6n+wQ7nT2hffv4H/RSTc04dgpkVjwR/PPrZK3IR9CW0QQTRc2DQg/gD
XXP/mEvwI70bJ4sY4xp+DqBf78kaGlLZ2SQo48d4ZqYCtwnm7bEne6srMsNjDyxvzxQWifxEG2qk
Q1krBb/oqJa/0il19Z/xMH2FfB7Wby4YeHsVoJ4wptWUBrsu6daqu2dZUntOX4jdY+6x/2pKA0NK
8SGmJo7E83J5+84E3JykFApqWI5svFK8RR64gzRuaOXv5QB8e93fnDNUnaHMF+axS2YgFeF/lwaz
GvmxLaPCyftgQCbuOR43ac/AMh5at9BK1uufwXfUaeffITtskffoxpDtrPCCpfB9/TIKJ73QiF4s
9PjDnU/omQs/bCblTswlZ0gsHI8inAvGZZqEzrw7AWzn3fRTqVq+IeuQ7SD9MDKsv5YmQNKIv01x
iVHonx21zisUpK/SQ0SxGzPPN/y3BYr6+35LqSTzXBU9KkshicT7snKIQfdEmTCUBSUzimEvYwwj
TBO+yKHxbBaPCPjakGAYpX20nz0fugObxMxKO9d7FaXvkTKmV4JMQOMocUc00gTCebmDoR3p+y27
h+5JKtn7Yo/3l1W/IDWfQp3RSdKocsmn3Xl0sqhPlH5dvO+sUz2cudVYP6d03Tw2LUJDfFnER6i8
u0alN/9NUwb9MMLBne9Gwk2COp0FVSuryixr+1V5jVyaEORoXq/TdvWZyXJ79h7acF0JqDjj1ozG
cuFVVc1gKnFZh2yf/KQ3g1mYOV9QRrbn9jsd37Zx7PzqU1DlPRvvwJDh5BhAYQ1LKyMqTIXD7GpW
oKUk5EJSI8t2rVU20aXvn/BjmP2QcmpubWPKR5YrPN4P6P3vM69FyM6IZ09n695tB9aQQcEgW9PN
c1xnObPnhgZRv+kPf/kDwVt6FEI3GrulOKiiGLkMRRns9M+ayutW4fxbcHlcrbo5G30zhqgvWexm
2tqgBYcKG//z5JgbC1cDQ1VE52wnKUPqj9amBN/dOHjE65C0dGBvyxcBMNhKoFhfpeoKCMv5H1HV
It7jC9zejlAMaHLIgcFbyJYI4gc6SWXsXTZy60SZ4fDN7qR6aOsMyg6+itFRU06QidzS5VezLZH0
nxkUx7V9zKYY2KvfGkF6XJfJ3GIUsBsCzpuHN+55vmdqHV6ASeCqYUcqHqFgW7RFXNBO6+OagxAy
HMbRFfN74XvEKSey1gd/El1mMPdOa+UEEecYGwSWRzmuIoLTcU6MjrCaZhhqDRt4LALF4TRd2OGA
OZpKG54bssEkgigq+vwQOcgoEm62jAiBjOqDjYxAhzRHtfEexuDn9jKBhEXOZoHIpbak4MePSJoB
eiNRJNhA9ycpA9/+IaM6HNT3enPECZwsUfkCDnO/kdlen0qgq4oh/sfMDMTylIUwaSjWMQ6qgNBO
okxZBlv54lx17Rj6MhGdBa9nZidR/cNOvMd1R2y0PvA7DDUGAo5qQq3YtI8hjnPscWBGt6juIcsm
3HP/+ic6M82jLWKSp5gqKd1KDcIMlOdFnKjE9zluDRx7FigUyp/AuacJHlqmKXiI6bi6d98kB8dX
VCNogQNjRAjXVpOJM59bnTodm7cY3hzHIHvcBJoWEHYNADGZ/4AdDPiM99Nn7T/amb4hokl0gU4P
eCXjCK41406/o00W/HC/DPFm07Unxef7zn8EjfqS9KCPe2ekxhQCSD6gudvGWrYVQP+Iz8OTo9Lg
nEcsHibNgRi3iX0HieIlR0H96Y4NDqtijNwT7gyQjUvHL+fiMLKyfswTx20LmO2OhPnd9Iw1+/zF
zLSP8lufPR8arsNZxX9XzPMBSTfIkGlj0rmwGl4z0jLNWZBemLsnqnikoXL3tqgiJAuZCwoOWya9
xSKpNgf4jQH485JFHUyMmfbrzu8eBA+pvCXpdQexzugyFYzQ/gr2AJw8LSmwF5jfbdAuqC7tG62l
DZu7dM5kDko2FIyNGwX09bMen+9jD2czJSPrPIYTAMQwLvYDWsIZPGjvMWtvQzah0fHNNM+smARt
X5JEhqd/2vHvolmx1jAG8Aei6vqLw0dLsRYAAy4GZKxs7XUuo42w4voutu/I09+S+CxADn61Vwqf
ULqZP2CpO4Rxr9n9M7ly1nRM55sId+ntl55pyJP69MpbsHniT6q7ZM1jSEkvLkC8dCKLN/kJaric
t5eWeRims5qDCdRJZZJImA66JeoogQgRowenYQCHrt5c8aNuzmYKWP4MA2edjB+SYQ1Hs2yO1fYO
L67c1bwiD5jc78SEpODNtIn2U9ppC2AxVDx7AHrvsfnolBYS6+HugONyjxntcz6tQQSmRrjJy7Yl
OBd6NztgEowYeeb9IhoWAUmtAoIY7A1O2yXVAW2kILpbhcc00YBtyayFVFUmwSV0EYU7pm648q7n
gTZstMEWuEhP7f3Xdp+ubN3oBAXE47Lv76H5YQWXuERjEuQaqbeAUASDvTPR+c0OlZ170AwaoRTC
DbEjH3Az9ZbkJY0+wjS0ycPwVTmijbteUrHp5fcP/YjSVw8C9wmAM+B5SM1VSNaaJeZ4WuGm6vdX
NHVcMk0jCsDQNN75eEdiSCUb41RGpV9a9pmEqDNcKcqxMkMPik/Ohl+adpCAFOEABHng9OFsvQAz
WDDi20dlOdvfy2N9/rVTEJFQrTcFzb+OX56OivoOwbSrlLtCl7ecx/WJapHfKDC4RuQU5DULq7eG
X2qet34rxGK0dgEApLsI+qRj4yl7mrS7LF40z0VnpSnA78Y69WdHKk6CpNkjJXdXX7mWgcGjmlN7
39y9hD63/oGnnarJpBlGwNH6UjOu6LwV7Wcc3/ZGT8UTj0yl5WeoLrjyH/yVhCRkNuu5LTV0QSXM
+J1HpaZ6rXJakBY9ppeFS8bUSQbWHOLO9kry7SMJfNob9PnTEUJ1tq10e72AAdYJvvIcMVSaBeaW
yGQtLyuj9h6e8hX6+iimke2MucR0k6qqchinbNeV4uBAieSnd/hgv+8M3X2bN4nFItQveBUOCgIU
VERTm6LGzIiGzsAf9a/yFG1zzAmoDmqMXxF+2cZ1zyUafgW0QWMRWURfer6yziI/AHSGipMNkNfY
ZfUU77tOuxcM2L1TT+Qsvbpq9Kzw3NI8Xqxl1n0WDfq6yat1hvs7HbH2D4zwvDHP/DQo+CZr5oxj
oXmm+Fb4ZmBGLOQewCAUkUtLGG1f4zQcLkuJpj2HL9CQYN0nZAVvYbgrYdOcmNq95JrV38XXAc7p
xlrYYH4f0HKczQ2wTHFDC59aaEwb8kE5jqTyZ15uhFsz1l7Sotf9fsWJmdu2oNb6Pvg7bbT8U/re
jqG8PTQqxANQy7718xuPehzW+bzTS4X0aZoBvp4vdbM1mV8h4nhWZ5z/fHRl4s+RLZIaARqVEk5D
pbJTwNGSjOr2VtV6fGmZNkgSOIW35odr+ieuLCLYj0xAHnQ0vRXGSaZvUPXsWGDNwD90OkKrjnFy
darV5yqR6UP4pM0SMfgnttdCh+ZEUVlV2LNciCxJb9cVvVkh+MwrIzmQ+W2f8pz1D0M8sHsE0skJ
beEZykfdi1YuGlRkDfSrrEu0L+LmXG5qsQavVwQzrh3jSgCnkH21b11q7G6JKMkHR/v/75DE3+oE
4qAz/WuR3XTvSmCPRbJF2xWBuZgsq8pcwWHaRe/lBh58YxdyBlAKujgBHaO6Godg0iViNlGMQMEk
rnvkL28N6XLuOp21HpbypgiGX9Q4iX59krHLeooDi6QqCcMtu4F25nczudADjFkhaejBFCe9jOD9
ASQJyZ72lNR+MEtkcvDuMAGxdSlZC+6RteWkUsOavAiTjzckC7MB+EpzZXajADXH3x4QlLFRlBC+
xj+9qO2jJgq32sohQAz6oDa8OZrZ4AYJ1u2BgiAencxXJh2ZeuAxZ+SxW/Q5bdazg6EFqH7/fMTI
qzT++9M1AFFLlk3k6wTe93iyeeO1UG72ZP3iFshHzqh43+b7+v0rwhraYeBT70jcqFyAzaVpX4IL
/isDjMnvYm2AAycR5ps6jVLmxpgUzwmXmA0+OzhPZUsf/gwqDj0MoAhKZaqOMXdMSi9iEHZc6Bvh
3Wq8oSNS+xW9+lN/vKAJY1SV2QvA8mg+TdNRAfV2S7lo2xfq+nMmrUMvyQGum4107ouOxp4QlUDA
tMnyr9IhDPiqd9Z/WyeHpgLSw2Ot+pKKCca5l+6Q5SjEYB8u8PJ+cptDJTJvdzqJiri885OFf6YD
V7ONUYTuIfkC52qTxN/PDTdbuMaYnyDu3JwzYGaDEkqQPpiqhXU5AkoL7QggXIha5pbJeuLvFw5p
TohDyQhFjNrGFMCgX/ec7NmGZtvFg6svG2COvkY1gsKIeL7lffsDcYHp6hCmCTa+DEmOJHfSPBmK
PvWmEcCzJyZCIbRVakfAfe4h8rxh+SE0+QZHlhIcl9cflVQj6uZ7yqSUyVbwDiLAKvkmJtS3JBBT
KcRQNRx28D0r/Mm+3fhY5QETxqkmFyGCwN5nLw3iP9wH4UAxpai0udR/IzoXbfDOUGyHCsY/dEHS
9q3O+cRz/sjSH1kijTMEFA/wr3+p7B3AP+oDSemoe+LbECt4T9LdtCX7x4b2bO8p3eMEWlp6EJ+A
xDv16nuz2oZeNfcF3ZcVx0m1WCCcDI13SkbLXqTzya7vPawpiL9OBXLdZW+J3FFksSGMC8Fs8V3S
a53H4uuGK7mPHUv712jCg/HYTLWqXhqHTz4ekDVthus4HoRJGnQPHL4xGW4CSa2uGAPqsFf4ZiI/
alfPum9iiXcr5jNp/dSM3qnLPI2kDW9H0cBGZe79EW7v0Np1BTJStxobwRZcRt/wxVoO5nLRDD4S
q8kCv1Vm8OilAqrAgR7eShi2knbFutZApAnMPTyP4t4aWeQ1qbdR9tiqTVblwz4JDHR/aeN74Kl+
xFl7SfhAisTX2+eB0lqfYWtccBAbtmzUGzTXVaLu0s7/qhxLJul1buCC5TWMZLYJklIZO7ICeyPm
X2vwHABbRL+yfR9I2zhe/K9cAuZ4kMg0Vbnww2+o6fNl8t0pwMG7P8j/lzicnjdYfrUbnIKrY8B8
xMZgINQGRM0U+IQutI+/vprUEnxkcOSZOlnTdGAUv3VY+RWMwcinUCEkmYwEtVuEn+uFB55IgTH8
q2hCik7XItqkYKJvFwDDGBu/Awdu+dKbCmeVeGtW50B6L4TeDU8JD4gKGB16oTCVIQ42+wgHIfaW
n5Bp5ylGKKOWLrcgI7wB9iS1F/W9cNxQU18m51ZGzzawfVrZfktJ6wN+KeYx5qnvdkEbvssjYJVF
BWv1oXXXxa36Wo7UJzogG2Y32GmvkpjjAf79ljgcy3sEtYiEES757NppDnlIoa7aAe1E9OZZzwwj
1xQvJs6tU0e1tpHeBtLwJ4VTqVpbJ3ap2NcPTgWnpTE3Y6h0L7iLPC3G8mtYuW4h93CuzBT4QB/L
g0tASN5+/bHl0GfOa34BZfe1Uv0d4UZomnhtarOg542yy5SPOLD8VWZlUz/KKoyzQDj3DII5oSsE
EkRr6XimQGjTieU/sSApTi62+NsQZnQmYIw9rS+Br8C7t5sB8IQgGLlbB7llyEAvttzKB3syrJCj
1noa/JU3Prb4oox2kfuD9GwbD3vlVoq3hBk0m+kRBgClT3fKd+w3Z36eeeREEx2COXbC/LZYG4yz
VIDSmdo0heMwzCThCxEO+teazu3aOrJjR6G8UT8lAxS0A/5OM9WsyCjVZ1qA6+TA6KUrlVjvKHpK
dk21ZaFJRh8GzY8vkxVCHFKBgPP+hgFWdB330r1F0WtDi4qFC73MV2HEOO9BPbN0+jpZ+/j5WGVv
rWP3Sg6K74uJrRuyIP4nT38jFxs9dsymBhLlm8ZFQKrM9YIJSrwkjsQcKRP+L7uiqtbvDCFlOwlC
gJDayeystbb4Hadv7UiAlyHU6Zyc43o3bO/dJ0DzRcjA49L99VteYpQv2IN7VJl9SyktMeriF3Z0
Yzy6+hrJIWz/DyK9OCZ7C/7dOdCKPSUnI6PreaSue7I2GXz3NIWP0o14vBbsNNdNWm+AuDeHZibE
5xUCWAGzE6TXOrrQ1cRrFrbE99lcjgjN6WU7xCN8GKyLMps0hZ2pOH0gpeJWkHl69VC5UJl7M9f6
89gUm03p5GSAaf8OxfnqKBAZifuVjjYDGCMqI4KNIHiyPl74p/jvi0se/Fz94D44D02WcHX5BWBa
XFdOLcqy8MqPNd/heuovkU8ODWnjkQKBrbHYoXyVvEnFDdxtYo12PKjkJpOjhu4+rADk4DphHohz
PxcglLgu0xR0UZgJoqSVbXd1hTyKlGZMOYHKfxqHG95j3wvEhE13mQReezu2h9RFcxfMaMRHA9ST
0JcOsqUCgMRILAyLS1VCm22piNmDMdxAbCpusuJKdcyFqyXrhV78AFFTVYva1aglth22vF0sxJGn
jV31JDblGc/PliI2OyyImPN0mSRP44YosUi5DuMsR1Wb712DKB8bceF7DoGiMFqn+fnqB7F1RmTt
e6I4+3cYfLHqeGsIbgescfL4tbgtxLZoVGCEnYOcIVuExxXsIzJpy+UJpAkkmBpH1asxK85+FV+p
iU1/eKPP9I+V63fj4CjvJZtjtYXVMnBAtfzh/S1BT2AbPk+fOMUjMB02ygqoZ0R2Gtxxa+HZ8Psx
dPq/rAfNCVrj+RT4GLsWOAu/noRP+Vw7sjn0FjXOmX0C6Jey60iZCGQ4J/dkosMLicagw6CP5ZJ4
I6Iq9lxRODK7vlXKGuBAyr+IgZNobJOFYft3nLalX719ndsIXxZEQ96nWJodhaCcZMGOdDm18Ewn
Lbjvrl3b5N2yA1TFAaEgrzBa890S/bbD/Gy0QS/25La45wcEnDeFRWaYKrmtvEYIAl/rWMJR12Dz
jt3S8jAY7m7U//E9icfAb5oy9zabTZWxYqMGrh2zgvYNx3OBsIrfy4dfr/fJFOPNGhLNoOw0eQRL
dAuvedNcTZgIL90GXvFuxMNYlCcS/tMaHZVE2Xdgz91smOO53EwmUW26foddEJWQwWAQz1e7HWXy
+9CQFQP2GUrAPiYv7J2KtFKWja06ttiTAgHN4+teY1cQ9xIrHKK3vOkw0SY9A2oJkW/X3MlSDa44
rcrAxvn+ah7WNFF3pYOLROvFwsmBC5SQ5KXdrM16NNkqq3Yu0AcABBhGVa75Sh2hmRjd2+c2+4Hi
YWA+jCOJ6H8Jo7QvHSaphkpygCG0IaKkhUqnP+VpUrYSMI81lD078IfzETP97P0jtEM3vE4Lmr56
Vc0lk8ToGVhSu2mEL38tMerxYfLR1f6sCm53p/NDK5SixfmXC/TWbLVcPxPC8aOgDNxI2o8hWb7Q
fqTj9ceb4N5cXM/Y5MIWdgRpTz/211YgKMnzfiwyxOnQz7WApC67vhToTg+yaNaLWulw/UFYQCwG
xOkkDooZt1tpRXkaIpUtniwqK3lpK1hH5i4NM5IHiK6sn2juFP5eIBkDz8me+KgVqMoYc3OFGD5t
wcNksII5G57hZSlANGb/ewUV875iypN7v+ak8LvBqHBDpSVq+JY4TSnVkxf69xwegNTqFA0GWFmh
YNK8Nl2vlBAA9swHUv1QjKdIi+8Zj+HEhSfUiYVvJdCW2LgVHzC/CQKguW1f/rQJhoNTl14UOno7
wAGmZ4/30SNwQvzbs3i1gvIbscjncxE1S7+0xHWT+2n9Sjv9IDfT3jr+4ZHJs6jfufgt0T9eANjb
XVgmNDG2AtgulAni/T5l2O/Qr6wRyLoHqC8ZZVroFk4nxHnGKS87qLOBEaxGpUB+vC97z8jFcwrO
NumqJPT/B8UPRLJIP2277t9uxl7vGe9MsQTSZsvS2qM3x7jz/WJfAeZvUCxE+LvDIK+1WOETcgHo
2YqCFBmuNSlCb5OjgHK8oWy819KkdfRfjpl3cLWFGfV7br4E/2YAZ6bSLSE7jRyclEgrDQrdPIJP
tc5ZNz4nqgTUB8BniES/GR6oy58oqmIsLs0Nm5K0orkltLnsdbLZaaabcwEGo6waqfwu7AttLmy7
YoVCUqlLYMmQVVxwYxz70CdvDvNUc+FCwTBU+o7r+Dttfqv0TaYqcKzeuS/FjFcPKb9Jb5zMU6/A
txozknpGbXRwQ47rikHHby7iADN0nbEKHqkvM5JZH/NHzhWK06nWT3Z0TVjcCATOT9yYdBSz1wg6
XL+VRuZ5POZXBjxxbw/AzT1/MNk/DzLcd5uHiQBBFaewhAJempcvZnRY+upshYX8VDacqdMUwOz4
FoH/mswNzhg/BJWZtGpIPfbsPY+ygV2veCgACmdde+N/O63Bwx2ONEwwNvyjwda18ssEktl4FHRu
r7tCm74z6rehUiEcnBQbm9TtJGM/Qzeyc+s8uAfys9tWc5HprZiMcv89AjS3LGYALjNs8stX91Oi
HMWb+wlWbDc13ot5jL4D346rrUxJFKZnda6A14KShMKmNo9eNQe86VL8NeIJu2S+BzvGvG3Cw1ZW
vlqtrcCvv04JcCZ3zKC4e/Xl184nwD7BKTzDX99cIaFX2DJl+hMbR5yu2SntOre/A3tQfI21lY3q
SYBG1TNgkPcmn0Rh+ydcBFEV4jFSsdDMcV7RRGqv5nwOaqedPG7SlQA/Z5P461mNutThQV5Bh2Yv
KnhLURvsweyw4X674NbQ9SgI3wT+4cjjNYBurnaSRsur2uwQJ0m0qrGI26a1bzOjTr55XhlVdkPZ
R/Jkcr1De4uH7kWlYLSRPW4nVSt8FG+VK9gsQfbXYhYrDp3uo+BGhpugNkP7k3F05+pi2N/VNWFM
ewSZjHYBncmugmQYl1jdNbtOe9vMRNQCfFaFJGST0MgPM97Noaj9Pd7cD8/clacGSP5VkRhDAEAi
bj3Gk18rkh24XWLS7XDLXlrrGQv5Yg+5q1sZa25BRycvSn59CW4SN6BWAgF6mMPdxT27+YNYki/a
oD4h0ZNkF888vhckvwHLlfOWp5JSX5fC0I1YSyedchT9CSZ77KVONOshmZFr7Sic96ZSFoxJgBWj
uTQAx+qTB5ECM+W5xlYwQ3YFfyIr8PcwDr9nSMqHV9lPahSZfUYW4dM1ieRrUOpFECg+GynJSdqa
Dpjkv1pGEo97VQsPHYUWyBKaGUZq8jne4VWbIAYRv8rW+gyHZMGFzAZubyKo2Kfs7Ct5+M6La6ha
wLeJg465bf32fyBfDzER75psWyI4yHp5D7LzRBsoQTX6+VPop42D3nNPigsr8qjK2ww7IDKSyF1D
+x80e5z7iwzwfB51f6+hqBI0H2Jxd+65hVcJbumSeprBoGcq3bcMMG6fOJqWyzedqvBl2Q1TkuxA
eu9G+HueTGd4dcGg9/k/18ud94EakxE5VDVt185n5K6MTQt0Y/ch55T/Isxsi5C3duRBdcuDvrUU
9eiZFKmfCf78G5aR8Upebe9Tb8SgiokzaON+U8imqR4SmKJzs4dJF1KLevP2mPeFF+KuxQlheW/T
JX7hAOrAKa3f+cFlOGWo/zaTo+vdb0tjZ0JCcEd5ybVF/jMQmmRfDL9DOcSysExWxMsd18TxrNjb
4VMZsPkgH7qQLxcebiYwZ4njigMZ8MOxbM1GdzA0VVfvtfQ2y3TvyC1tzHtvZC18ZgvTsLwUE0Yx
p3U3gUkqn/cB//rsESQJlrVf6I7IjujVGwIbnjzKJNERGNkfq48CPCSCaBBx05R3zDJLhj9fOhM8
CPPTNkJUgCyaqra3kOzll4DrzTEfadv9gb9fJBm7e5aUqG1UXwrUQB1mhJGvROz2xLT/bC8x1JuE
izKmK/SOanF5e07JAexIWUtOLlE4vQM+Rwvz7p3Pv0lO0ct8hAkoiDroScAEgK5N7cioYmdmIkvL
T9Wq8VjMk5NVI0lgmbE4i5V5/moqxOKPd/8VAkqhe5s6B9dRUt8Yxywc9kDNzTuuSUcR2Ivulr5v
lttRTCt3Hmv7eXDmekHa1J4R/T9lWYADxWxZMfD/IMgH8JTOLrVKt0HaXyj10EaOz/n6PjWbBh+y
Rf7TujcRNVfWO/g7asFlyPBtlkResj/deHXasFYQYjF77Gu5u0SdO9FtaU8np8cHZF03B0RdGFBK
doN/st+je2ngttu6zPUWZvIM2i2gXS7/yq6VwYQGo6+5ASkzohym7+xMh935PPyjcYbDVcG0XfAm
MGz53H4gcbqMzU34W6pGdEyOh4gz1Ma4ad/BJXqr4c7jPfwwaAkI2ga+lxTiKsuurNHnFixFXiHp
iYatnrzPLT3QRTm97dsvpPtaIkax8b8W35ANGmgdGTZKxfd7Fu7qocRR3DNPuhQaKpGt55hoFrOH
nWocGZHeqHk2kq8D/yU4cR71Gx0rffvrjS6WArpsZaLz3KKYafpk5PJAD+hVTMlvxlRRzXNPIkXq
N7EJ2S1PIQzmwSn1GP85fuYXIagPOkozwHyM0nsR+VDL6tnefs24taAOcs9bE45srOYU/9SCf0xt
QsREX70PV1We7BsymGofuwlhy91bBmB5/mqdYvR8pQG4WeT4ZwklnlwcIJb2nMwszJbV9lhuRlpK
cjYbRP0iy/ETQvTmdpMEdmjBZ1HLO6TOx9n3YtlImt0SFpuftuhOCwWPVST0YoMegt1iOt6Jzqba
3/VOiXWdS7h6JMyLr6OUNBqD6C9L/Oz5wpbvVlUBCip7m7pzLqdlLNuVIQGP8psgCXvBleCHJSP9
t0PxPnj6juFUR1KOJ//iVSPAgju4ou4oRwtQMq+rQwrObX1/ciZOpGZPN6Rb1kVR1MK7Kgh/B/5e
WwQOs/WOKH7FdyZTkvE+Lpg4bhfaZoUR4SfBKUONsM1Xz8UxydYWu5OAeEfO+5PcqWg7md9sKeG9
OTl633CqA3jaGnVMjRD6cxMWscftk3aegwxBzC0bB6ghGKyJLoA1n1/m546NxQUvFIWkm0+wxrfb
aRLRibsE2zXDfrL+kjgzU6kF6GR/fMIhGkOPREXF6Bkat2cmKiv0O9EnNTh8Nh9mGUMYymmEpM83
a6hmvSqzGl97hzOuKJ5XTDRsdaL6R02DaMwQyp/wGbBRyHd7GjEkgLjqoDOlt4uuIRox7ajDi8iG
yThLVGLnqsnGuhH1fOcKCss/V6jlg1SK2wKxJLLmRTUiJ0lc70wgv1hnglnF6+a5A6Jele8Be3py
cUCl2unEOYGijrhaRPO42s51FfSH1mlg1rk+3Er75tjbIhuUIAG+wPWVEnsZkqLTEgHWGofrGmT2
e8LdzhV3n48A30qERvpbjMjQqlCHXZOhjBVMge5gXvqWUDYYz8EdZQOHUGRobQIjMZwc14AGrcBD
OUz/qBY34qo7kVQq/y3oWx/W09uBtzMYxDWn+KyawaxblNE5U522wfpOgzjztx+vrTvsv2mgymE3
35vxxYttpDTM/Ca6hMgeUkpYeUlUVjRtyf/rlX4Zd3siVGp52eO1bWd0BSag4bShaLlU66WN13/S
csrgRehBxXMGLhD0lP7glKDgmBykODrZXabO2XbmC/khdKNExRemvl19g6a7TDM9kmMHpJv6PMfG
tPF7dsmZ4SbUcDIYrMgWolKUWAg8SM/y+5DNkCQaEnSDmYC70gWJwkNI5FgHmmDDM0B82tU44udn
V+5LkVW0Oqz509B06Dt5iHxvhPVTsbrJzhKyz7V6HlRGEcTyF/SAtnzg78odgZ01QdSogCFoo/on
BBkhVA58pemH/K1qFZMFviamuiwqBaXDjk2VojXjfWvXIaT9OjpyaXbGUALxRNf0b+njtfocl4q5
kryvYpivwam9vUc2XFjqzhXZ6JmrrSxTvMIfDJXZJtbLIZaJ99een3Ny4sdI0Rl7mJCsQqaezvOx
LrN8g0w+FMGYJ7Hr23ouRPbJELIBaPsR4EDOSg9Fy8jDd8uG0J8290eIwQsmSiAUmyjRxr1h/8Dd
NRMIgqDgNRtVyfAhmmrzqOfJ5nwTwgtWqdRvhldmXNPlzXIUdeDHZjhR54GNaoVVfmvgWvOqUjAT
BrAGOLUCja0uRnT4+VmY5nWhqkAQkOea2qYOYq8EYubHR9wAOxqlP9PkMJHhUhS+GKuaRdYRq/pp
HJCssL9708BgQkhjrqzfaq4jcXAoKDH965UWDXdAW+v1u8Ol4kh/bhpfzi6vDiA2BrgmxlRDFUd/
RorEewsUmknROvUO6ds8U5w5O/6dIHPHGfUYq5j1OOkVv8LcSHRTjFoM9iBDOEXHBxkEJaSxsQmp
lyIkfFPxOpM6++gh6dtTZY3UZIYFaizfQlfG7vcbyl5VeT0YOkEyysqItEyS4vvjt9ARo2akm6o6
ZKu7m2bWLSACpDF9M0HrPKRRLCqD4SjjpBHD5UlzTreXI4jpGuYtuZf1DFkuP7HeCDkHOvsjNXSQ
NIuhXrDxvVQ08l0Vmrsq+O68Lbk8wWo9U9pCc5QxTfb9LkahLrCrA/67YW3LXD/3p+q7YkjtpzEb
9lz03dzniB5OGwGneSqJ8U/5CZGdn7XImNiI7OnUoRPEI7UJv4p8xobohrri6iuSC74NvXoNRtGN
AQk56snWj1jBsb972428YmfsMloYgZcWZziSri0Ijz/VMrSs0nBuMBwbl97dLGhz+YQzyXXPAxnq
VtawJmdz/5r+aozVZrlof7pt9WPUXTHZvwMVTKm+KlB1DsGg8zemoruaTWOesCO8rw+dItLfCfdH
IlzKS2CxWV7fdcZKRFujk7BqzoP20wJNyf+ubsuHnOJ52qo3P6a48xYngfrMMupPW/I/Z0pnMcqx
YQX94o3ZT1X3EopoMp9a3JDJzjk4PrIBOxuGfEjiaUwWd1CeX3bTR+dofw20U7RYSkpFBu1G7k6V
mp1ZIuF//655TssyWlOhF/mvtX/tzAphsvF5/MsKyivikB/QN8sgvEvjOeCKDB8tAcNoOdwDVShG
Vpc3UDsgEhk4WMiRZqBGxogMcunA05jvRes4YtLH/Qb3G1XZP0Q2CtxPUtLK38y/Fnbe7LfkjGLQ
Ryaohn4nlgs7DHfCb8D1qcti2IUc4rNtvFNB+RILSQliQWG0pbo85CdGEO9yReljoBKjZmB+ZffV
QMo/aNJzoTe7Aw85W256fOybPEN2eMzNJ5M/JhqZOauT02pASyM2Gu/ti8iIod60NTmOEgqBp/ba
4Qvdf//ib9DCfZPMP2OfHRU8q809tFZ68JNndwsQy21Oxh2VGtRtu40KFWTeCP8pLipCbMwRZMq2
yYgLF39QmQWgpMb3lFGbSs/zw2ngC5hp4PeH1baqVfX8kuFtmXeMw4eXJaHh3WBjBclZubywj6oh
rU+cjPZQXgwkUwueQSGq5UjlYRmwPZBGoqD32oadY8BI8gHht3/mWmqgBziCiN0rVGWILmvqDTMF
nYiHeuRF/LXwOf0yvHqYusGRE4FQPt4S3FiVqdggm5fk878yiih3FXS2Bj4kRwcapDwfqla3x+n3
4u9wRnINKDl7ceLOhJdncbrPLqidQlicA0Pq0KwiVRRPpnPPyXgok69/hsg2v+1gA2rIQ63S1vhD
GYAFHLcB8QEaOjINBXq+vP8fy/QBiUHXvRseSwXuVC+pIqo3aW5rgRBk9UjeWYjCrTO9i/qbDN5x
c8Y/9wha/NgtpEslPEDkjHngQFArsZr4HzEEt6ruWQgU9WsLTohPTYbLboXvyDCMuS66mI5cVisY
gQp2Clx2NlZy+UgOXPYH7S3F3uPd2ViXteRuq671v46V/cCxdU+A+1SfgjPWDEdtRRFWpNDDDNvh
TxdzS0Yx8rWLnVYaexlFgE6dBkNcs6BzLokfNBGkwlCE329BPk+qHXsu/6hnNMfYtztddqQesu/g
GJaHVKGcMrtup91V0EGUgKPuK7qYlCDC7vPfYJHAZJtaFFc+nPe09CBtOCoQvUSYBuvF9H19IiBm
JuO94qcfZTcj4+4pKweEgUxZBZiWUbWtyZneL11+wsPEsEpUAkpb1rc47g5VzxLylt4k3Z9ORbNZ
f2r5c8zYizJKCfMVKay0eZRj/I1p7L1kXjhY5oFU2KqeXOWx1DpNgn1DjrFsWD0b1lrQEsWgB3M0
pXYhT6gO1MgF2lUhwseV03YLmLJZ1U82YI7t/PlvvTtmJx8Kw+i8j2klJ9Tetp8J38rTjWz9h69M
p0IXBqS+H3eYTXBiwcQGqEwPNKcg5KVZbPyS9xELjmP8T1FBcr9ZpuuxR4HaERM1c9+3goYjxMVS
FrkK1amefmJhnm/kZEj0O+9LNl55CLduNvk2xpncpniKqA/pVSsRvWtCeQu07A3GGQRTxirWgJq5
0EEqVH5NOGB+8nv4NOZirLqnDOB2sv+/z6e4rOeg0BWWZPo2y9zTQnt5g0LCSkIdHGTSHw8Ddh0t
52lJgSVSLPiZeYW7NXLgD6RF7q0lIB67YK6vPMI64mjWYzC9/RceJthl0L7N8O0Qrdm2+NFnLL9G
4OGxnPErc+AvBj0maUMJbbahfAJNXxNgRgR+Xli8D1bGp2mUMhQQQaxwj2fQnh6waJtH4fJAzCDM
9c8j6FTGbR/jUQ4r9HYzHYiNVURcVhCkDiezkzUqB0tjAaSihW2+uNA7++3Eb0BvR2XdmH9KZ4vq
PJ5tgMvdIv3Rizdb5yLjNDU2GHgCMYC+3ekgx6HPBtJuunBZsR8wAeCpjRIscyseujQk2RZAlea/
t0hXjJzNqaxTgBK9T0jrNjGqxMmQVCBu7fuEtXDuG3k6c+CRyV/D7p8V2pD2FnoAPWF0RtyQWrBm
Nx0Jbup6eY/FKwalMpVcQDZ30WaEb9GP45CP9GbDvyR+CGBaspCqI2mMQ1MEJpNomPmMx8VSHb4X
X2dpEs6t1SyKvyqI0M5Bp4Y6uVXIQ9EIfp7rYJtRSou5MGXOXVOTyMmrJHIVShG3C845L//jkOCx
KfmTgr6Cjh8bsvLF/Pii0PTiFSOepr+0nXpCvru7gHDtuyQQg2do0UQIFFrqQ07G7brMcGRYC7w8
MSUF71gVmZoN2xS6gogPcXV7tqx0I4txh7ByqtpvSWmpHhfnQgUjkT86otOPU5NMPM6qv714hhfd
sDSyi5Zi+SbY4q6tCvWKkKdvM4acRWlAL34Q9CrvZrYJ3Moybu2Fg3Ifh3M+ffjVFuGTDaUPznvZ
aeKPlTyHCngLcNlDf4E0MDIYAu3dM8R0eEzrvNhnhutQxVrwXIgYfkbMLGdqsvOpJGy7Jn3SZBM1
NEIMkxn1CB19hs7UvdWiH2pMT+tMN6PqTt2Oyv90tknmQ6xnCwXk2IDR2tZhRf8wcAnLJNUYXt6F
byy/ycw2hy/YRiok6bRAkYPjPg/s+VMUK9tBZKA5JzySRe5k096xcX9rv8WOFyAiLSizKZgRnyHD
gdiHMBFAzWF0SG+W4mQ73vjWJwztuY9Dlk+qtbQZqe1Gig5hUsmZjNLsfwLZ0Cb/wwUJhV/Jn/E1
tDPDll+JUSw0OIY7O3J32io3HkdO4TZRrzo9gErSdhZZ0N2W7DYhko2GSQJxzccIIeMeSsAQ1sep
vMiVFzoslwCPfgURcfVd091+QoV0xhnA9sqvD3KlM+gf3RbQh02ba+j/rH/tkgZIq1aUl6DAAFkL
LxvNW/n7vaiupOdS/V3YoyQn8L1HwR0Yr9SHJ0ni0/dGnkyp8099OcQ5Vd2URutZvGKll5fpG7xU
gvKrFg/Urb4zxOp/kOpAS4fwFqwd+bGS0BxM7FuMRrvIl2JyUbDen68maypoYTMJLc86kOU9xgZm
z2g/Pjjm0tX6kYJz28tJfzIZ01uPCflKPqMhBOPf+iKOv1jfGlVvEKjRH4O9hp3N5Uj7iFp3WCpv
ROm/03EQulMoz97/k9is5UJrnT9gg/+cioCGJtgAFu7JshWmAm/rslE+cRzHYmamt53vh7o9klw7
5bE9ha1yabR+I86nlV2e4pOuIOosKQREYqdnoF+uUt8DOyhOgDA9gT6iAf3MznOu496WA2KcLBQE
HJYBk89LmqNmqkUwsOsAmMjkgKeK/2xjc9psZd506C8/ZEUyaesSsUDh3yRMnIGile9hLrLEjVZS
48X8G8MBlzCNOxtHgJAnZ07mpv87sLZzRju6BYiaQdUKh3yD85LB9+v7wRKJDGZ3rhfhzRp7Ulwi
wUTFKMkYJCTirBdebXtwLhXtT2Ry6usgY+sxVxpb1MmKfnaiJJVs2J8iKoDSDfKc08rsp3hNceEX
I+iKLjY++XEronJRO2VhktiHVbkp2SlDPG+yd4swWg4h6Bi1D0ek0DN7vAtMRjGQdWhmv8EpQf97
HYf32neghOQqPsRUFaJBj5rZMMDwmEY0qN4Ky9GB2e4IblIMk+ha2EVj+FAp+XfsLUagXQr/rvym
6TKjtfBjqHWbYshliiyqlhgvy1Ik7BEV3A6rz4eXiAMm+QV88irgK+OryEalIrOf5D7fgWltfcTg
Zi7FV3egFJ2+CtS7WG5Ei9/mryTUXD4vAHittMVHSMe2pykFRpgJBL5bvTZ88Pzd29iOKyRcBx8J
sjtodL1pBAUt108qwsEODkwFmuCUWwGaGCTBm8Q+GNZN3zyhp0LY6Su/8DmW+RnpBVLjJPlk0cGv
2sAjtHwh/wYRTzLSh3V+7UtQWETb/l8gDzGYipYeiShKrJdg/njKD/3AtvApcL+gjPqwpnjvltKO
o7dkO+lgGusI1WZPsCMYDk6vChUkr55f9AUac6XXRrFTr2IHdL8ZzOCX2sWPmq1hMjRSHaIEk7L+
QtbXXQJ52+f64U4wQs01Wl647Z1FXboKG5f6j6s5AOya9y6MxnduyfC02pY8rMi12GV1io2EzwSZ
UUlfQZyWrpdG5fUJkEHOyxkM8xpk8twfbnBRjPuZly57c6NvneSrp/9klco7sTNLc9Qfaa8DERqm
lXG+gNiaavuQLWEwAMPuunYnNX2QceaPNM9NHUTLN7CThmEfJRcrjXf+mHji4I+sofcU/2G36aN8
mWPrZzmkC+rMzpRl30yi00QhDpXh0cPHGRclfmyhgu2bk9imh4JjIPzJoRcF9iZiWmdDuZpbkBvx
Qifjt4lkv73KQvn5C9HpSwc7ql233/nvbemH5r0porFQwEf0I+UY17A2ul/0vtM+v5EGjI4cSdmm
8Y1r1Yb3xtIPO2aMR8bt1plqmpvpxHQ8davZO98y+Ml48xeAIGaCxDDIFmYYB/jCu5Dpm5/qFomb
wAJ9wjoB46JMv5mHyNa2ILGLctKtIwQlHNYvo5Cjebwamu/XJKb21bFAdTfiG8lafQeCYcuAD1Gr
km21WGEpmlFmoemQXgCL6X+veubE3ieDa9+akvcFd2XwTRuoKyFVu7nIO59vnVdRqXUMwANXTKBB
YMeo6Enx3fo28quq9caZk7aojIk4GQZaBtn9/S6soSCG5wyikLbbz06IilN2iPxDd0i5SW7Pu+t2
I/p5r0WgN0L3D5dzj65x+akeNq5mFuT29Qr9lFnkLrC7TKquRqoR3r6t95SfewinLdqjUyIxdP2Z
1dD9QWI4FyPBe92Rxu9XM2/hmVYfNhkyqIpPHCm2uJNXzZtZqDgbOMqs7FEWqPVd6EFxSKBo3z1U
k2tHvhQzc8LAcCvjNzsLRLU7xgU/bbyB/NDpEOYGQMveCcrminb2u9X8m/0rHUKNdRjnlf2MgX70
3PogkreMjq81MBnbTgDiolpVNO0raTmPugQYuUwl7HeZyK62m7a0xMPthDx30WEEJmnPeYHnxGT5
TpqRONwEfRAT972mxfUZbaAwkujjn3icB5pSmgu4yHiRA/IxgFL6EemFX5zATTV8+ggDvCq8B6Xy
moAmpP29mCjopoS4IvTIWcAUMKqHdPuvN9YFFS/8VwG+LgMS193AUaQxEFcyzpoX/oPNa2pyG934
ufD35uQA5VNz5LnStQHOam6YfSOksTsNmJq8TSeJsanIrvtIOO44u0YmOolUlq9KM2GuKDpEghEE
hX0q8V37YtC64aVWsCCdhdinX6n4RG1wXtj/Uu7DgzKNCN12EWW4d/Ux/nZwbDF5jbyMaA/o8s6J
AxA2b6XN4Q3rfAp2uX7P2/7isu0lOo33Y56XQhAO1GWLN6mKoBYWabotCPDI78zEj1V+ltK+8mua
9AEKuUZ+gVUxLq51a+5jkiiVRh8xOAqz8kgfrEhzQ+3TiZp9Ks+0ujrqufIk7iP9LUNCHNrPEN1V
BXvv0yTZTfhOVsHOExkBU9LI1rlWQ0tVMavFxO2ZBG0cKYrBxvgYUX33vCu6YwqcVWVJ4MICwcgx
/e1c5Cre6yvSjuSDVau/HsA2xbe9cynjGhAJYgD6K7Z/TCARJUFPUT3HYxJzypAOhjxkcg72oiv4
z2WkeCdncyQDOPpIprUeB0A0dzkPWRv5QeuM5GOcsaRXFIaniK1DQhoz9oOupr5KjKbzpDS6bBUv
quapXRvkVt5yuvlzZ+LXJ8YNJs9jE1ufXplc8kz+qC2OWQ7sZlnnaxXSZIrdiX/4vc9z5t9yjMKI
axOeN52LtYwN8Qgqp+6G4ShUcf68FlLRJAqS6fdrpDucBI07vtOEt+kTnibxMNJ6S5Mxeqs9GiZl
IAeohQ2kGfS1IVtxMezCYBaBjTio4oCbvI9amdW+MN2kGJMxjLdGJIuHKzDgxDynZhP6qcnWJkCk
z8xPKIm7CafH+yqeGLmfCktQr9kpiENHriAcvC+IxIppjwaKRzPjQd4P+8n5kJmapGXQ0VH4AYrS
7uMXy9EDoH7Liu1crQ81DMwlb6p3jhnL2Q+LCu8OuctCdMeH9Pkj6JVYaP6+CTPzE4V1rUw8wO9W
HyqZMMdXPxoU0e8WywnW4V3iOeXJgyYRDB7HyBDD4YpJnAEr69fVsiASDPazXnPIidQ/EbNIMWLN
TGRAqqREJfhZkgrcV/734ageK4APfVM/D4Rk8EpN9z9/1HqDqRJ3L9Xv2Y7WM2PE9nDisBs8Czdp
0Z9GZnAhUw7gxuszXXjbrwrxmmxpVETyAqCspQ1OFTmJL3lEjq8Ioa4lPRK5uiGYLSu+QuoL36zh
0Lgc1FDxEXHLhCMbEE/Oio9Nkj31oC2/erI/1CDQUHbBN1VRjDDpBe2bncWz9gzTqSvTfNr/REye
QGDF5vijD2rCzAiXJDrVq8PCYdCSPCEQq2RpRZhT20hbT6HIIlbiwPBl6yBmePwn4pf7gGcESTug
mwnLEzsecWh7LCnvCPKWyEY5wccDMMi1ndgY3IaLDUqDJNHtbTGkYNBT/eL1DYG1AQKsNgenDDzX
7Pmcyw+tYW97enLluoLwOqdFHdVspcrJrtVZZhdPtJiP+BukmYLm1QYWzOFIkB0R4G4wOxg1d97W
tNnH1NIIf78HLe2k8e8kxiA82fJ+JTLh/UYRrZfB3pINI6VyWmuPtCbm9jnwxPyWj9yRHWqdSdUA
vCpq3bfNm4XSD/4dcsljyCK4OaS8qaV9xXa4JH4RMmR96ExhubBzP3vyfWWB75f/dlvkkRW+KThN
JHcR5zjHGpsWuEN2RkTmoWROYESClpYaDbk6OeMXWYXhMH3W/BWhuORaDm19gRDZUMEoayR8ltHF
X/hYYxu/hxPvIVPNC3eJ+4huSS5oXyyvhrLywU+4srGJ79qIAIFyQFyx5WWznhUeT/79lt+B+tGO
xjvgsYV/07zIXa17dB4eYUlCKbzLXa9/8zoFH++OKNIIo7IKmA6S1d0XeBBxA+l6OH2UFJPqx2EF
zJZr5dDgoOfXcRdSROOHJC9ucRiOdhlzJY3gKLqNcs/yLHmXitt7VIHC5ryM5VgWr0JmjXEM5eqm
26PwohTrpV0NKoXaiK6vb8xUknpiXJipIGwqFuF9RqLvICNJilBE/EWZ2zE/So0wbuV4qBiLl2vN
TJ8OpKwonaLkvVgSDjve0/+5lOxXTjA6I8h63NcfdwPR1SrQW+4xYk+CpaM54S+7peQKv7/C1VYo
Ym+rC79+8cNdoualsNHpnOY753P1C43x92RA1c8g8JP+hAXT07cH+NzvleSbPemcOhj3ThMhRffw
UlGZd8dHuJ01+U0mj/zIEcXoPuHERqPJYzHIPhucf8oHHjsZIEKEiTxaku8VEnBtpSWbXf1/C852
aJPoh79vseWDd8/bE47YgU4YUbSXckKKqr5BMWPI0Pto8x/x5uz/pzTwDrK+3k4sEcoifrC5sun2
ISTPKhvSHcGqHS3yjFo7K7G5dA8ylG4wMrepr+aaahsIVEdmhnNB0482AU/W43utjYGOWtNASJxP
QcKrwgux99FtyXJxuytNHpr2SFzwTxk9ENBRHCkA4K09ayPYzBv5fJRGW8bhziG3E2YdACIZtZiN
L8yEEGJ4Ge5kJQ2jX0N5PpdZ4DKZKsOIThrhuarok/nLGCx/VsGUn2Sewt7FKYsXfME7F+E5kGYu
PlnBFKNV5SyshTMF8d6cSVXQhYfxUmXNDvjJ+6TKZVNcfUNChN3gjtOkCWQwykwuNxw+iUUOcsU4
mbdE6/2biP1Zf4xzdH+zVsZnZ+K5OoPoEMCRTJF5P+GWzy56ggH2b8UEnp43P7xclFvbNtNa1ZW5
PDXtQp16LNNlEtCv6FVhPo8Z1iwTSbcyd9GrJFAK/R2Xzrh+wscRt95+DrNzek5ZTe17YWvA3k1L
oi7SPPQucZb+youd0Jw0mW3cHMY/XEIJNUhTNFvftwdfEIy1E4tG5I5F4Go+Fx2JXPS4PO8Angfz
itEXD2xSHhsRjhXP88SsRRDsd0JbQdpLgBOSLCwckuUsxDJQ7w6cEkC0ZPr0aeuIGXfS97fpe6WH
48DScdLWiQEG30rcTO64m4T08p2rLzAJRwjw9+KjUx6TIv4Oa7T+gYiS8d9bKBqUWENMcomHwPaq
woAAkdFPp60RBoLPbIfuu56FtpxONHyC4biOQ9Q8SXxMX0K1Vm3BJxg9spNqNifL8VE+gmmYax0i
wtdsZW5oEfn1tNzr096c6lUqXINeVb3iz/A1qEi8Gar1HhyqvSRHPopxPNw9FHnSxurcofyKPx/L
Aiz0Z90p8vbzgZeUzLaohLbyyVDt3tDutNEzR7jrD3CYFCpEb+p4oOaYLx2IVEI/BctgLPI/XJg1
JvxTukubKpWYzy2VOl1EUB4ZSfutAKMHI/NprlFl2L/Jt+WO2nN+22rT5dsmnHknazWwv92DXyI7
L3zbr6Mg9y3CxM2ULpvsI/W6buDfAUGwRjaA7WQzWurKIAZZ1dUSz8nzm2OLMX7/dEs8X/ThRK4r
ivfGZk6SLEwJbfY8T8Ye/cs7iSUnyBcp1zdgSYNuUm1pXjkwUNtsUXoxMj6dXkMRYXu45ebFRUDw
O60+1ADo2Xktx1oxch9HBB1gnXg7t1djvhgFaCYzbzDLQjIR1+WQjQSHstSkWqkJE8FQFuUtehq4
v/24TcjHGfF8mtRF9xubOubbNOqHES+p0WKMmT62Qh+KfqzRwdp8tYW8Z5dowkyOqhZ1qkJ1kqeJ
WjQ5ESBvFRppdfzBhRcaSOjDaXlsufFXBgxGQX/zbgpeJ6chR3Pu9JrCdWjEaeYrAf1cZqfuLd6T
z5HCHAx0btqARvpYDmgN0hAD9Donkvsve/AAovtmaHwhZvTnnwCk/1+qHsD8tq/rFUMYfZiyyTxh
xmfjxocDQKJIxlYQIHBM6tQ4jrdW0twetQgbsg3TBHN6rUxxiLwbAhrd0TX157O3JQchnuZxuuZS
OHCYN1/CvERpV9Q0r4JVvxkEl4nSbNpIq2QdfGKMGilrRCNfrihmKDpJUUa2nws5KucFWAXjkq89
Vgm6VZHDrZA5o1C/JC2ln414t2okehO0yb338wCHLU7NLxRRmUPgHZlSFGKpi2OAjmxMNxAi55E+
j7N23iJBIwxPWRlDjY3l8rL4OG9FAOC7KqD3Sl+Qy3jffubZcW5WOTPqF4aaMgqeS95sWHlclF/a
m20gcuQg2jskWGRtYMJxi963Tb1LeZmIZ31zXjCWWMbuGxVLBaMSDU9rX/FFY2OW386ACKAp/vXS
4Sask7GRVXmvs+JjTaSkn4FhWjcMw/COodlrigy4jL6aoPwbXoyXKlgMxQMf4LT5BaoyX/+Tn+jP
PeYbeVzZESVg5Z37SgJIO0Utqi0TQzzbuQPejLKsyp3JhY4+57M+WY5vmYiL+5CXWr6PS9GmesQT
/GGc2wF0qHpMp55eTP/9IMaAZx/6J1KrFONAS3W/qd/s0H4zBl9E4cwqJaycjQh7HvXOjEljhAGQ
purQGHVSiVTsKLhcYSRQFE5y4hKnZIvKO6VX6qIEOnr+ijqdu2wiWst+tdXJjiuIfNROmtVakriA
KgdCIMN+GqK5PaAdbbO63tEjnc0rdtBq6fgYiNNQmfo6qVhPy/qwNwC/fCznj+M/wohpHZBAsI1k
CcVmvZXor06H+9jQPPC4+YGyQal3wNEW1apL3X9p5/eKWbRyk6ORQhMaxwBSbVkS+rApsZWrF7St
1n7tdmFo0IOQ7YFc+R/06Cc+b4ph+8wtaWSJH/JK+KCPDBFUkQ98Yrx6jBHt5z6bujI0DIXhIlbZ
qnCrU2w6/hN/9qvZLfW/5W9RSbs+rHfERC2jqUIysLlNvDyOYERfsLD4GIMJji6eOoSUNGiFNlMF
vdQIwoj7AMxM9k5GZa/17087018L4lsRRbOvViuReM1I+9/z/PtoBbZjCq1ozVYRwJnbscsWw3YU
IwUuoTpaqKQChs97urs1fdaZdu17PUL1G1KLChBAc9kTmAksvqNgRuOBjm8Zyc/WyvWPtj2bPcVX
uKYQFjEqtBABATr+Cf9gE18UIU/JmjS1T9e011sPon5pyXJtHHWitzrbBJvdw19xbc5CZrqA9uaZ
IjbyxfMjyUgonGljGyAuS73D+aB82LCe8/Zp5oMOvl43aporBwhlwDyW4/ggGYPiIUXx0YQwlDSp
yYxNBJMSalkchgjshIRlfoSxyGmubGyWrH+4i3bEN7FNV8FvB/TbwDbwIrJAUMIDmyW7g1joixie
xggRrVZzq9TnP0+EPKB9fCxf81G6g4s3BXg4QzpEo2ixSl1FDPu9CS8cA3FEwe3LDJlWnNY+kBPQ
uf9+rLlgF1yzftKSNpolIP6by9Bot5NXN5D6X+B3J1tBfTY6AMsen7uXS7pO0NGcqdpw1q2OU9CS
fEorD4ZOC+h6sQaqImn7njZChMV8ixN828TxWM6LKACaYO3JKDW9d+klK58Gdg1Krxo0CeLxPELo
1WQXhT2jdHcbYjNeg3YvmWySvGeuL1q4jPIg7D/xdFSHEdmFXpMEAXdGvA/r+XKm3WwHRTYJH0Ol
rEAEnBpS+IKmNMs8f/eo0KjWwvSOeTsoCM/6SaLZCSv5uUeDFKUa6Hx/ZDk639D9dP5W0epK2v/a
lrGPr7YcP9CdLycMxAYtCF/0cN3G75nyPzb8Wrn0E7MpfZ4DF6Cn2KCcdzGFggwqyypfoDYdHCdt
uPyH6OJ4YhS88ehoUSSlLGrvaWftQ/XEhPxVKTlgjpEZZkQFYkpKl9W0KTb2FGBYAkn8sv9tGkcA
Kh65EO1eFjKjoNkMHEOPYAg0fHpc26N6aM5sbFq4vasTkD+Tl+MHNkWxGfIg/MxJBYSbcnJWlWmp
VVr4lZuoybqM4a8bRdzzsk96Hr0xuXwfDcq5dU7Mw/Sk/5HEQlj+vX91hk7ztSCBoi4YBK3C7n9a
yGxzdssycyKrsIWrY/ESsR6GOjhGVSvtqqzAFqWSKe6wURGUQ5CBRwIdbS816HyOjeq0XUDc/Iph
7xpJUgLRzqgi0erl6D3O04AGczq8YWhn/XlIOj9dl+NhXq6GM7c3TnTKWRlmFRADoadVX95VgESl
gn/wtvZpImUe2DJ6atJ3dp3yOWtUmvendne8C2BFjcvSuULWKLMpxIMdWOqSf87zjj12aIMsvl0G
J+Q//cAn1ZCxCPsy9HE06+bg9xfHLYoz8yYcBMgXwFasGajUD7MwCxk35ofy8gcbG1eCAeQSv03r
T+eT6/xlhw6Q8gFVDJ9Y2GD+bzOXuhPDF1O031ZF6ImeybO1IA8sO8buCdj62cnEIcdNtMub/EC1
hR2udaDMsk6eCJFfu8t7RvenonWzoSk6rQbmpbF56wU53DnOV8wDxl8xtU89O0xFuKF60j2ZKLxb
t1cjLiCNb9YoVdhT3PpVRjdsFWhSXYY2TJCAZ8E1eFtUUDUpzYAEfTZKLEDLUIO+i/k8lXuQswzh
3bJDH4Tk6pWV10ueP/4uG89yR8KDPWsBqSPbKaNObdSVjISndU0dT+akwLyEI74qny3iVRkRGgkf
Y395wG+2XAL1aYiOEwBZhBz7msq4IBC+fEyrTsb1ciunq5AFwGbP5n8Hd/7Ar8qfjxacu7ffHXYV
bn2KVdho29Vqf+kn2eR0Q6QWJbBWkF+yYmO5rUPimQqHZGemkM2NaVjm5PohAK8PwR9n1okUKQZb
5KPGIKSf2tAydibrrO0bZGMYGbNS7PlzBo2U9SWlky9sSp0/fSbbHKwRRc0GDfHvS/w5sQaXVbxK
USj+ZMJcHmFv9OtUqXzDZ+WZ5UKTjOg6P/FfrFCRe84nKV5ctcYIbYZXeirmalSKkNmwmyWepmkc
B5m3Khd/hgc9dxrj8xViJgmGzrjfak4/M5aSUb5GVAvVOJKBkF4XSDQbKXfQY8aTDTl/StBUguE6
zQQl6aFQafHihlAbrrwCGDErt6NeIKEZiHoFCWK0si8Z2mSZiQdGtOnDAQGRFDC1Qwn7r/vu3VvO
qyFilei6uxLJ+v7jGx0G6RLFNjxkd9jweQHiWe3RytEOgM9jLoHCmVDUIxNJT0ALksb/SSkYc+PX
5+g3ZJL4g35WxGdblAi31KsmRSYap2ZNllgnyT+iArUspfqOJ/JHjJ9NRH5RjW4PLWW0vQ/L+U6k
vABTrOTOuuX/OUVGfWhXxXIW0hsdCZIO5L1PN8Rt5xZEGuXP+e6ET2s1AK4OtC3yTOK5WvxoWo9A
JeN1LDrgN6tzSmWuWzCJe/RyZeLwBUuuK92XWv3zWKYAfH0Hy9mdOOFJP246c9iym3NfO8gYMBvf
iXkfNElWCHWDRcPtr0pS+yXPwv5BEQDiZbi36a0oNKfFrn8O4FPQ03SWwIzXJIQT7b7qNf8TRgyJ
y7uVqSKy9r7TgjRz7FlIwiWznXqiQ+liYcwHsBOqlGb7SDvIxHI59Of7CfXhTCi/nPtQ3EVR6lvt
VAHFQjBJvwdPsLXnsgofwCkMYzNxIv1Xn43acMvILRqEKPVeWCLZSoDLP7jux6ae4Y6M40HrUrer
iqqSnjYjMXPt3JDe68fBq9lak8xIr4QTmM++kkLBtqKlJf9aU+nQ8teBeoseF2FPRIC6JWlQ8Dzh
tX3g4cXKPT1qDlFxU0XGvwmvyFmPwTIySOZzBCUzYa7u8MT+Et5cJfNJx17/ocDD9LXXpSSv+gH4
NxNYo9hOWPkXCLU4BeX/7InKQQ51KzKX4j80Y9GpHYevAN/N/vTAXurnoi1gkYAmrnGEzpLQt0pt
bGXJ7K/PRtxxBRCjmPLkrS6td8piaraY+2y3N0HmU6+LBzajWwABKUaLZzX5FXtQBYL2IplMkk4D
VrybyVzX5SVJkkEwJQFXj+n+832Ii4482NRVkXh1awD101GJaq6uJ2ekAHJC2vGVy6tCfRnkVDWx
D3wDAh4S++t4MO3K6CZTmTSBTqieRQwT7jiuZ3SYAleT9XjiC7dKbtuoDauY0h5AIZ9YzA2Uilkr
GZBC40+VQjKzdHKE05iugnUx99DwExwokicjShHnNJcM9K2RKhJgWxLStQOVp1H06RLyFL41K2a1
fSDsPJ353SjE0lbsj62yVVHGiaZHhFnU+BOXG1SBf5ZKa8LfnJFQEF7SQH8z+YZuoGixmbGQgibZ
y9o+5yf8kKEwRQVYVJfN+spJWxnp7g9MAsd68O18BLLajZykpwN99Gk9fGuhu4KT+GPYTHog1tIJ
oBpRejwySVSvSjY/jIBFrwIpwePJf2+g0MaazGLNpFbA7hP+4jssiVxtoJdjFjn1Qs3qes+FB1ZJ
Ar9ONqRkZ+wQlSgQns397RyI1y6/aHLOF8zm4SypZE0ael1qZID40yEjXZ9/OvrTpoC1nPSL5Tfn
vQ9/N/w+kQ1GdllIEEm0BOkcIGjTLeC8WXxWFH0m7kEVD6UumlR//KVDgafPru8g8xTqUJsdDwPq
7aqCO9tzRnOj+Bn9r//LoO8CrKl02gLdFBS+n1dFJnxVJdxOBr0XuDAd7yVDmXD1Ihio5N2nE14n
9VfnJDlgEXbjopWmvWNi+ptRi1vJ++glrKCcHzjXkCRtyHufJrqlWP+VaNc7tXxYoTgkgNOBjcyn
D9xISp3hnXtrPVQPI5aC8FFutQLPiXIzCHpQCyvE26AoIMXifRsPbx11FFTIyedb1ZCF/mrpEIKf
RWiZ2vDF8gQrz8LdHabLtyoY5RkRmC56+/9vseD4RAquyfehCrvQmBFnpA0K+rSutRsTfgxGpHOe
4iU6GMh5Z2aUdqeRfJ2T1wZLkDuZBweZlTnDXgwjTEhuYaxXYViP6Ar1l770UfQGjNZ7s0xqk4fE
NVqyBUn+rOpO4wIR7+vZZUipUtGJ+R6Llx5JzLjMC+ycwULcy2hSxrgZ6qzS//mKrkOGd0Ot5hg3
fr1vbiVCZZWMBrx1Xj2V0x3oOFr90zZKcicKtEpvcnF8sWPI2Sv2EA3tUCDgx9dP5hLJ6d3F5V4z
IIwWSP7yvmBPpEftxXhtfQUbFZxU/wYCtUCjtHU6aiJly6wyvwkGF9IO4/+rwh7r3yJCQKiDfLRo
3X+UuQMluBdNF0QwimHHex6WGuDJCq3eSdsL0XelkNR85SAhbyqi43AqKEKLHb6BdMec6LS9arbd
X1f6QX21REvrdWeRVjP9sm+VGDehB14Ye5a8qk/XgCzjWdZpqAMZ8YNetdcmxNwA67TczIOImK99
883kxZzMRCrrenrwzl/Q/WhstkWDoGViAIGvbSl2TU4QwAuSpLm+7M2gWyVKmmK3Btl4iHP3mbhF
iRb0VPnAvDELBvBv/USCZ2jDk7/EhIOQDbB9VHqAOZg4k+HZSfXKS3n+K8GY9WqfKN8dp4puboZy
iVh6uD1EQcyA5HBP8HBHk4rjvuGo8KDQRP4SkX3Uj3IMkYNKWUAbPwp4PObSPBrwfmTgniMUU7+k
KY2oLXjfkZmLInZoSl1LKP6EIHN6mzxSlASXzAWV+DSveK95jFTuT/8vsjBP7cIFWS+QIHO+ruer
MaxO+Ss4lQmN5iyTeY2GVGzBLoKbxhexVih1EwRyxItpYvXXnCVXuEIUujjOnbGbTjEH51BOdaWr
LuHh8H27gu2roUr5i/PTIQXMQzhxc9ifqBA/3eDLgC2+KKcogsdah9uodFk8okUl5lhI5gyqifuZ
ACuRhjiWH+BSD61lV0msBzjKVCIIk4p8MWhQYISZx/iDkgXE4grk8xmxZGgLfOWvbgw+elHh9zgI
AHkTpuo3JuhsgxoSKTu+WmG3kTo3yq0sVlGJfVZJmbHojlDgFlMHsaxQ52ILHtBs73xiiKAwe5sX
crCeGWp2QpGaEvoVMeWjWhDBZlEU+4z3/K0/jtSThw1wonOluRP/fuTdGXVxCSazj1IP6HWO5/o5
gzO5EFjWrRElLsYjn9uuu+JDxOCB7hMHNYTVHuA615W5kM2CfeNqcEV7hK7euSTUXc8apmxdb8t1
WR7xAT0Y9Zdu+CuY6RN6LOdQnfaRFto03Poxtz2ULMqgU7Sllv6svqVNI7fywYFAMi2Fv+J6ZbZ0
VCompmMRtEW/JIZPPioOUPV/DTpr213w+/J69NaPDcAtqeVjZaEeOwFiKTx808NnEpfQcpKf4CKq
7H6OfObovTYheeI8uv4FNERSQTRyuGIG3BFgf/WNTqa3moqxFNITiEjWj6lSPFKvlD8EcUeljlnY
ZeFexWPizrI5vxF8ksS7hrRpj7qfgb6y4Tlmwge+dy/9tCsos6N7nG60EcypnaGJHf302v5Ty0Zg
Kmm4otwHKOO9vSfj4rpR4GMuxy+g3IaMSVGkgNWmlfs7aGsPF6YyfPFBkvbOaaKtBj5S9whFmRMC
kLXMaQGRAi3Gc0ngs7WVWS56sKDQLEyYoDkOkeP+0rinJ2LTCSy2Ub79NOgV2rf1fuuzKeHEz/Mr
v1TH3+kiaIVIaOKx9v8LlU1v7P5nqmOzYnc9QSF8M9l6uGFjwWnzN2OGsu9AMaD9mCrremlwEiZe
zdM3AiD8SGX10Peb3hXT/RmJmEAoMLwoni4w0VMyi0puQDbZRhX/KlBy6D7tlSi4CW9hLCgCzds9
tlVMWBR1wsZUGbRWM+EhhVYjSMzaKLZsdKal8Yl4wIOJpupGJ05IW2cbMeMIpYsrDI86BHX+cv6O
PeH7xl1ZIiiSqdc92tHvr1tZwug06n+uymrUYHOUpVGsUSFcxuT6p4KG9DWdKsNjqJSAa8m2OPq+
Edq7yvSkpYv49avRh74RKRJxdAZlOwPGjqYRkM98W1q60sZIxmrbnzG0zCOkOXmdCFdJ1MDR5ts2
/nsZIBAGcCml34tPmv2Hmf3attc6t87sHgCTGTQue/aRXe39IV2kseLy6+EsWYzLb9DQ3uVkNWY9
49n0BplTUtPEj5Vz3wokgDc7iFj1tx4KqahzMKT1SoqW7ZgmucLLJ3eeqkzR6ctVdWygHUYHHZfm
xCPUromUjSKrkADPoj4iAoRxHisRl1zJSFZc2v3itsIxu306C1HDesu6yzTGB+EpPLHcs6AIAcSy
7dLxk/ODk/nK/cGg2B9Xfdf4WJozVrRGBBej5G5mCsRKqoSVIe6IRf4+VZ08r+Jnn8xqy+eQljfL
pG6nfx6qFYhPcnWFWOeDog+wpH2dy5YAeoVN4jpTH4P5WpzJtU6/HYdP3n9DKL2BEL364Gp5vJjv
sD0TTv0CWl6njGOyMIVJtl053fihziaHzMeVy+ruiy/hvM65rD8w2ZDsV4zjFVoILQHvYRiJ/gUo
KlSa18mtWCfsfA19HBQl9FLiR6raMa9cpNM5boFfcknhA7kxDaNKtkptWRgUymTrLTX86QlXmk4a
So09y5igdB8f3fzkjfurtLs9Se6ZpT4ln0SAtmqTn6PwG4n5FBs3tlx61016fLV8mwL+ASVXFE1q
4zx7/iSvneWYbC2mU/ZVY3zSyLIbIWSAVp3riqUPswZeEttnIGAooDSBbgeI628Agt7ilXGwXjBO
0UBcdm2PAt2NaXeEuO7WsRrC8C3hMx4VhpA8eIG7MPRwN8tBz6Q0s5d28A2Cb+R7KQWsRqOJC8KZ
OmUQTselqbmlRCNMU7AvYRnv6TJ1QDQeWHjIF50KBlFuQTginbdJco4l9hCHQQA/ZWzGmc5Dewvj
SgH8vrfF3sB7ucImgEpR/dIKigTcyBuwkAPv/rYJQ+ILeUbw5xmjzRh8KwkbTDmAGtlNf5EatHEa
jrXdPTBcgyECouQ1s9+tAJRBlfCGvPJ0as8WVANxThkRiPBjvMxR3yvXOvze2ijEu5QylgOLbd2B
tR5FW3Mjn9319S2dl4Dpx3Gx4e/QaSjMQjK5tEm43cbkEWidloQrTvtfa88O+To8yZTLv9Q3bwru
Q209hXnJpRkydtFM4OxNQ9JP/7x69QbHayHPUk4z5nL9BE3lFik6D63Tav9vJHp3ACJxcuJfs28p
a/hVmF/53WvlgcFTIc61t1AqnsfheW0uR/xCuyuM/S+8lqkkLZDN7jBvjVKur0p8a4/gZcjVm52M
goPguWzpA3utaY9tUhDdKuHLZEKezU9LwqtY2tOhGosRMOQ6w0V0NDGuOoU+pA31gf9kQG0U6Lm1
ymVPcWEgLS9nSMbsTyZsZEMS488gpKowQnHcwXKqdKAuaqYFGOHy1iZ+JPW796p8UajnOZIanSql
XuU2FseiGZCh8lXnDSLu9alJBOWqAM+R1MXsjQEbkf8XojUV9U1rtJet1QkS60+D59uyvvgt2ugN
ybJHLpany8b9pg1PzwjUHRq8fAiAio79TYbpnKm8W+OT0x8FvF37fGNzUs7HImX80oZ0bOy70Puw
M+qio6vu7HI8NEuj5HLu1VQ24OPkhCChRLeGJYDAvKBW8dwKZZc+vcyqz0dHU55g3z3WbS1/Q6Ej
8Z+HZ13v8Cm2MIJSRqXMhWNsmvzYr9jCJAc2A6SApNmkexcEIlkSc/m7gZK1R6UbufYjjq/Ok7JS
hJSuGfqTtEOc6/+j0fiP1FWvuQYJS5FRKUd1TiGYqFND8mE2aAhRBN3OeLtcoLR1IBn1vNUn4j+u
WEMnyrGNBdkGRC7+3RQVuxUbW2sT9xjOFja24nm8xz5JPDZvoP0LBzZJF9DTI+npq84JpnwDxhsK
V/1wIyYtFq2vXXgLyaunai7sPR8v80w8NXIp39btvYPr/EN6Mj1uPpEMdqaC+Foq81Lj84fcCSO7
LfZJBM63mcjLaVXB66uCfoWV/iZVGHib9issgmVN4EIu+Mf6gKrJV6PmBeWjIE7sqDyRzNDlfDmn
BZInXVXhRDzuNZE3Y7ndJbYO/lhYiyej2qj4vdoDPnFGHRL/SmvQmagskhja3I/k8UGxzmW+xluS
OaNJ2k36zUFLfd6MUMmgW0SERpOnkvjrvfwPTJWxzu4L1ILim8/2r61uWrhDxb/qOdOa1nlvITlw
iV8LhTycZ7nBu9s3q6LI/XuuinFeiAu+H7b7k79a8hhnWKBe8xthBw1WYW0yudPv2j+qmdpw5WGY
BrH8c8WWMJWZzhLA5XVZY2dkn3roBAXcaXJgucimc5NVhGC21G6lSyf5Lm+GY8YhgwFmk38KxWlg
Vd+L6iIIYL43aOQrl1eq/jl7RTmC5OqGMTgt6Iw1zd9hjcTPp+sbEu8LvadHsUoPWZkmLv2SB8VF
hSf8JAil23+PDAl2NsdD2YJ4gcktmfGoPqW/Lgi253Jv0Mqx8QVoFB7an7wa6T0nNuzdxV43KfDy
jYxIRtcuBljNSN8ppVlrOGTKk201LoUNbxfzABLPcaCu5LV4Ju/foh/0Bacc+0Zd2zCjYaBiFZQS
WOb+yD95K27S7IsHo8qg8y/0K7RU7nzy8a6iDMhOiiZJz0A3fqnfKzRiqsRtDL0NALoEVFCoC1Lr
wHrpQCf9WKgDrynQJQ3064RlFznPpdLeCRsoyk1YDL/HTtXtqMYm5APFiJKxC4CqdS9xdaez9kNs
dm8+1vCf35zceUPqvTYIumgk/51cXW5dubHXDRCVxWkpnFnVp7jcfUhRRoXRjt6eYSGa1tIP8PMm
Ym6TAGHy579i8gvEJV6te1Mien/ufqLO7RI4rVq/O0GjG4lpdoCDRcR0Wv/4F3MVX8Z0HfOQ7eTh
Cg+rW6JlCaVdfr2lc2aqkGNfNJOLOnVkAZQJo1IxPkIPQI5o6eBBpwXXJMctqiAEJ5tFPDa0CsWH
6FvcQEku02ZJdQk3EIsJQxjEs1ite78GR9Dn262OxvqpZW4zuxMl7LqMU6qN2AZeWmrDaiFPnSbY
EXjOYNU2X3kQWCnS/OmiINVW3bgBOCngvUYy2b+dcy/ZoHWsOPQ0Fb3x5qsgHTbt/sjy4iO2jB8U
KyIY5jyuwcbPT9SIVQXbQN8l35bJAthGohLvcWTmyEUXzSWdfpZzV/MtkixRGMpNtWUCTNVyXkP4
Hk7lmsxLChAlgE+zajiQcL0As73Kz14JiDZOi4sSQXqSpxq6qhuuhjz63xdKbUtfMoG2uYLM4kBb
nCksOweZJ1a3+gzXomC4XYPBqf4gw+LTu3bP5dvOo1fvmE0/PbTBLXHIAKq9AhUr9mSwY62AD8t1
reKcvx/qddzbsOlxTFfYE8JrAJjY/0AnuFN3o0lSTuPwB/mN6oTTeYO/LlhugyS3m5yan0I/ovAe
h72EHuLcvqd5gslG88BhrG3nDFgyArIQZ2q7I1FDw4KBsWd2hTzMJ9Xv2pl+YtgpDya2NfDH5Gyd
/jgRKy3cCMmbrvOBrYBU3uGnGOlYtyXd8Yy0PNyWyGW/n1Ads5CfPSX7yLP8upYvCz6TeLWey5J6
Q19Slt53ABXgjl5G5HEv/+Awcela++eQwpUV6N6qxmMOhHMPfvSRSwL0nsdu4ZvFwoIrBMn0NX7y
rBbZQpnAuAERP08sB15ZjgGwFcrspY3m2UUh6B5+FjcsSR67SrAgv/KoMKhE+vDvHEvkOUoqCEJ3
UI3f0wLHscGHPpmnnX5a6wyvFF7sRyQvVMp+/UDt71HoU97/ADoNz+xCz5dZisOs6+jJsPDxih/X
4LFPF0za3wXHqVeWg8CNgKEfxzgepVjy6r7JaCzKZIM6HgkqsXfLnPf/JBpE5Tx6SHv7ZzBS8dTt
n1rv+ffQ+zr9mjyd4QuIxdfc7R3CUSxuD3+pbULIWWNEv9a6OBGJHD5ASmRrZb35dpJ8LmL86L3E
DOdp2NGOVfZDKtGxNe7BHx4OGkE95Jvmd/o+632+KfBqHJbrZeBIU8Vl5ELbaKy4SmKO3yc6Pcg1
lq6fdIlibp8OC9PmMTHnxo4QwEJu/lS1uLPloKwDtDPbTw8xNNJvb1+gp13hRk/IFxH5VriTUtnj
gms6aNn2py9DzgjFc4StG0aYb2W4K3vMU7gvIVDMqKS0Ao1YEVqCfgbUVbzjACECk3dXWWasE2Er
z/MdES8TXljwjLB3nuspJAz1pNRGXO7nqdKR5jeom0x0H4+JVHoTsoRABizlZ03k8sh1fLl13NG7
0MQ1T/BMUc4L+ho1TiM99xg8cH6O41Qzm+YP3zvb3hVL9WYWI/mMU2XSKihkRPHfHBGGKUg6yrH/
a0C34lGf6rNV1xzGnROauZq49kPATSDsd/EFsz+MhtcoTfNs9MEkv5/J0EaWcv7Knbuq7shmn+8V
XJMtEraLoNzODCVlX2/PFWURovgGzc+cbYPB5a9cn2WSzLPRzIebrqq5R0VqRPCrZwrd/9SXbBBR
7af8G+1hoT8JuPZ+DIJUu7xZGN9i+cFmfS3TlA3NP2diSNKYIoRJmYdoPeFWsCrHvHuj5kj55660
lxyaC7c/8CScYotX9lDXITrgE41H3QcwcdkssupfON999LxJHmNt4p2Qi5xoeFSyQnz28K24yFPb
VkncQuqNTQFMXBhwHryOk8TlWUeDkgQ90R6Vf5gJctMC5KU5SIvkB2Avzefo+Hak1LCKCsea6O0m
pM5+EUCyyKkqpCqNVqxUOLxqYWY9ZRBoMdHpUxNLvRsp12z7onpuzZhnMpBoQQVNHPvBlzG4Z4iP
hoseM/X2zFkarADw5wQI6Lw+6Y2nastdE7CtNImMXS59t8xk9ZypAWtJdaauKtWLRd+vRKFxNuFp
fTlGqUgEBpnqIN+6tBnKX+g+URpMKlqyVSv0G/A3InaKJewdoTy+LPk67x1FcXy9RG8BiAHUxAoE
aqwwX3F+eL7FXF8E2+frXJr6b9l6ReeHNCRDA+wdRqHjqX3mfvbppviUJBspI8liF59P5YvaXqvf
dEE/fcJTvVYRTjZvcSGH8e3cxF+aDPJXZf3YFHKRv+SpDPD/2PTVyVFYyBzcUszR5n8OEHkVKqoM
Wb9aAWxJR8HE8p2RkG1bM6DmVQwMWXwalqt6TZB4G/Gsm5JpjEZ3c3l1kfPsQVMNpjqEN5G7q5ld
QMsDXUhbz6K+8VBXgW0dTC+lE7+5fLoTa4OL156R94XHPN3jdxwwQEj8/gP5tul1dQ7c9aZDs9fW
jsTNzYFtLX1rOXakikZ8F6Nu6sGOxau7iDm0br90C5AZbqmlPxotjYadkhlGpjtJpjVBWJfR5MUt
iPg4xpCIT2OTnncb3km962HIphi7SADgFFwWCzQ+IkXwWX2PIlkBbgq7KgBR1KoLAjb5k1G4g6ck
HsguL8k8MtlbsBlfJjnSAeJ4iftf+P3+mZndoQon/mX246eSQhfPZtVjawqasb/pss5UaFS/KkSh
4VJ8aGxNx07ujiVbY2ALufn3Sy8B/uW7MijBJuQn2KE/c0nU3p0w3S3JLzY+i/lp1mPkIEsZKGoj
hBg8tCIw+rQ9UQHEP8Wd5nfIiuC/mJYMn+l/wea/vZbFOXxe/kVFeYjy7wChnBVejn1ILobQ1wgf
Y27nBpIAr4hZDnouIPR7Kh4Sivn6oWVNZqJNyPRe/8uPikkbQV4FZWcKj4G6SnUC9DNOiHbW0ACV
aIlA4L6OU1y2GDCvoKnmu7YxE7/lBWexgPlUir3nxL5rp/DScWzEXKkK5qeb/So6Q4O5myqfzeUu
6Zc2aKY0kbce0Y3xM5hCK5H+OJ3GC2Fb7KscNVuLqyWEYuDZCKQ1LqYeliUQLNJ1ShGAe4KNOtKW
wtf/Q2H0JRettkazOD6KXvaZvhv29R+h385weK6Gz2EckK03m/aPyr+E7tvg2wpBvW4yKzy+Eqwu
RvUXdoCbRoYwzVKaJxq5kFG8Xqdk5r5kXtjwnrC4HiFMsUD2rvk95i02eOQYmdgwxZeK2vXXW7Sv
byoCTS6iFaI4gzYxPLQKXeq7mBNIodBGi7+eipvUp/Jrdvprk4dP/volS7/0S/0opLQP6VkFVRdc
41r6gkMRkGgclfQaAmxAc5nn6fBzYU620dPoUM5I6LU4kWgI2AiThLyJXdxS5vCNG4Pjuwat8QxB
IjLMi5IqHcYUCsp3edKgUa8oky5XSdlvbyDbftmetOiw2xIaf+msVnjYotwDCT+Pnxh8eVRuGFgP
Ds7oatYRwAC98zqdH+/FnaEpP6L6c3QybHuvnh7jrQLskCAUk1O4frIRMqjXnrHCUvHviZW0QLNP
CTkX4JK+BcdztD9vQXr9RQF1QHMe+NAzfUXLnhkwhqqz6IErKGjAu8JH/l9onVdk3x9PLp+gDm2g
WlKb2nUP+hJGgdVZj7hf/t5tB/6SBOJJW1ajLlW/+cqPcadt+DucKheRpYs/HzNSA9oIqUrjMsI2
rrgmwxs3sN+xtP07ARv9YNh851AhtWaAlxZt2DXvQHsSW4zfI5CfcpgzY1xi9pFiOo7E+2U33o9J
wY/og9Va3jgQ34jZ/NJ36gRK1/QY7PGQlOLo4FVUWUvP06MsWU4X9r2YCKjtMfoKPW5209pF0ZJ0
ySiL+VOA6Nz1sPD32/+35z8oHB26IyyUAAbqxOccIzcObMKB/gLqJribH8Qu0D5e61ZIH9TBFfO8
oqA+wzIgjpshaSGjaK3+tey8HWFRRZBE5cWnFyIbkDXhPz5DM0r5zZifG1SMDliudbWfFA9lJe8F
WMaSMxttnZiVx3PCqDRgFExG6PMkeABPWhms4p82jW+nXlWW44m4F34KCX08jH2xfYKeZyaS8WAX
TVkKEJxxGrA9+mohtmvi4/gpL+sc2q4H4zMYyQOIP4IhboM2sP9PzyA8PqarYk9/PejmRfJ2DTWY
cSw6iSP1U+TO1NJytuP0WHnDozElxwRBtV3r6g+Stge2LdRUECSK9OBQckjJfovRQnHl/Uj6/Y38
+4B3ITrOAFFaEMyiypKO2ZANlhC97dnZS4xtg+BdH5yF4lynyVlMTziIXKVZZkMy7X85UtMZvSL1
u6vaYcYKMoH8yxBH4M/WIz3KaSzDCbYosl2m1GjhAv4tNDrFlaE8FvLrTg0H0n++zukRz7fYSqmC
YPEJ/cpWpG/taIXdkkd5dXLmH7EbllTrP4YISDseDKDN/33eWmWjUbNcEX4Q7bMZ5+zjEKwAlSC0
JsQmfUmLpp3v2+BB8uemY0PaaOhnMhLwM+Zxk230y14bj9hX8KngnAULsoL+nDYSe9UpP7dg+Mvs
H4nfQZAfiv3F17IBhxfNJ5GVcCc8T1Nf8NQN/zQBDJRtIrclrIjlG1sTJpUirpSoSFuIB9UIkzl9
R1NK6t1TY5t6XGBAoqaAt9AxaHwJHi8ioc303YMewFTvm7w7OymlrkRlfPTFUBry4voSFS4zyFy+
Fl26A5o3S443/Hw1CAEgDFNQ5YifAbRnUQpZHOSq/MwAMbTt3+/ZKAtEprX2WbshvHToQHIQPc48
0MAogp1N7gm4YBoVNNzmEaE30F73RBhdEBAs/DgZdX3hb7ZAlulrxzz+fDUo7ELmV1jkzFPX45aY
93LqEL6xb68Z7NQAVHRWzTxcRhqclvRB9DNlYONZcZ7b454D45+V4DwpsbmzoeE7EFeQ64CgCDt1
1jJCTtQZNYlC0CPmGgeqgjSYEFpFUKknyB1lkS4elaH8D4j9bYsXUpSILWGwmY3r4ECEZeTeQwxK
XAS/N51D9BnTBCbg4eR/T6KpW83OTTF1iro6t5IAVJpuJNSTdvf5f4j4nujcQ5b7xkEv7B4nNAGj
UcG3XrBTjPMCH5d5oT7hZtH0+2M8j1rrtv6dmZUhO6jUTrJD5qnWu/cPcUDsjaV+QxvBpN6yrd8v
dtYEZOpZqMYC7Ekd/VV3buM1zXfdAldEm8hKXMeysntacvTj+sxK1mLcIA6Q0xdvMU+8AYzUcDgE
2xl8zfHnCF6qFrm5JIP4Tq+4pRf4ccFO2ueXaBv99lvI/3FQr78meug1o16ZjB9SSBhWxO1B9qxI
a06SG1vKNMLVIsC3/u0+FpcyEh/DVPFkTsPtJMCHg18vag88gqyiSXtVmGDPaKV0pPq/wVuAU7YW
WPXYAg/LnYJOAPHPO5eZtdXLELiRq32/ApH5QnRF/dHckKjdYzAbr1/WkT+djC7XB7hR3an5r/Al
UW4oeoM6n8B53wLjykUv3eQXEv/XUyoekiqRMU6zbwHjguFH1ef76QctZ8ewBX1nf81IrWtxgzwe
fJQhnpoCgS2XgIwYu6Rrlm7QaUoMcU0/iEApOvNTOKEtn9s6JBjFubFrtApwDw8NLBmQms99SND0
Ot9R5Np43a3Q1lECUw2P0WpCmcw8dBd6YN9OpRYBKO4Q6yzRKJVvBTtscU0c3TZ/CacPeraGCpcO
hstGW/QVzSV/q42kmh0kN3PM8Pa+RWTywtA0lDWl5E6XvGke1q+yt2xnBC8YRy4AxAyP0yl1B/97
IwsXW0wCsDS9L97Qt5+gyYuEn6AcbOlEABh2+cudHurN7nfL3amdpIeG2AqLL/iSPFoUzq0ts5D/
6kEmj6IbyQemk2ecx9yin/ENSnd2Xw3dB4OaRjhBVt4yCvHx/fpJ8xsNQf7BfMb2yLJdv5Te3rXf
WYdJsl540fuHCRtFKaV2Ti8SCF1M0JuLq08RKgS1fseaKXuivk3u+/5Tf4jiYec7ZMvjYKMdyTvE
BHahycfoKE3DwdXqJdVvIFWbizp8HJ1/NcJVmWFDgGu7SLVj40pfhAuX8HsaQLD61ISfziSp2gBj
q+5obpSRdbRnTdRzINFhKYZHlIrkaKWJp2s6IxhX9/OBAM11fpkOkVUF6ZluwjJMzSvlJjUraIMx
toncB6pL4I/Qjhc2JrcEeKDaVc8IStIwSj5FWyjDx8z3Wy0csIl5pNjL5zMT7taaEDkSxr9LvjQa
52Xjj5SvJcYHDmWCbEjXySvj27AMQDxhPSfwnmiD2YtP0ugvjha3l1TQ2Ky9++GouvdsMXocJKW1
R5NkyLFrRJ/xaeUTLyNvzoN8/HLlLO6z1FjA32HsW28nLQx5eVbrRcI4UtGEzTV5S7FIvi21qQzK
NgGhw0gjr4cWi4BwUueYcLsmdemphGDcJ5EQnu5dfUHTzmr5kL8QT8JA1O13OZSCKbXSAlvkdcEh
DUzJBZ38Q2KgsMCSvpo0apXbNC43U+Fh80kWXy/sSTSP45hkWEfYAWC02QeHIv8hcZuWsBAgXS0E
u+s+91tanGNRvPtExWIJDsMFIZFciw8T44IicaySoKMS2YgVTqt938VDQL1gIKVfvBkoDTILmb+O
kQBRlxiaIL05+BCSuhYX5c6oaRBAa1/ERu38umHhjqO+RhERxII2MSX8PICR92LGaQEyidSL7F1p
5Olw7FFYXcjxUdVoP2/tg3Yhx4kYPa6wEIdR+i/KcoxBxwNHsmK/twd851W8Vet8yBPvk4AA2B+D
+EOmeO/V/vU8gsC0GR96yq13YHIoWStpwoeEtkGqwckcj5UyUqiI4Jn3G8RB5RBKP/T8h3jN6pN9
NMb7h0re3nJaSQvpq/BDAc0a8rfxOBF1w8JttUoqIW20H+NAbKfQQUMSvpMcPUCXe+O1Oj7zxW+R
qKhPUO6w0wLYBX9aElKNFclqo/CIR/zDkWVIO11wXYVpNFVu3Rqv4Cse22k1AMJjZGPPZyov+QwZ
f0YYu9BfkxtPdCwGL37bUmRHqAcgPHNhhm5LUZLlfxZnVGDeg2guZR2oDN/p3ngX3eSy8KKP1zNj
CAFJm1up7dhKGhY4Za54p43QkdFAjJGgkJtGRDx1UdKXpxcSZ/ym4CbnvnNZ3lmVHy4VFrN8D4L8
WuP0Pk3oBoDQkb5ytvS1nsBtLUhWDhsciTfyEj38vJEhOX9nwKTlFAO8F/a+plVUIcAkZa+dl/KU
OJv7uUk8ZpSUic9eZVTsnqI7ZNHLkGnuX6dKklEpSbkaoL4bU0NQ6ygni6ip+iGlWtVERtLFLTen
IhPsqzZWhoRm4h4Tz274cuOC6kphyeq1Y/S7OiOtKF//taWuM6m8P+STCh7xaAp3IOMjNBFni1Yd
TzScT8wfV/YlTdxPekbazXbaydiE9j1ALFhFhuRsTZXiR88Ka6sE+Mr3lHEjRRRXhFJ0CBhFUiZr
qsGFmYMKl007r1bNLdGdAxwMoM+JZQF8lQMd13EqgE3ODFvOKzLmZVht8QK7Rh9d0L1YPR/PKjlR
x5+mvkSXX+hqXdQyRLZa1xGC+RWD4mNuGdHGwMMtAXqVZhAGSVSazgYsXOCLaYzIJnInPYquGaJq
QDykuyCS455W+lUngw5j1yf0eel/ABYsKMBZxEc6j3r5ag8bMJJTaAsy322Nrw8liRP4Hyb/GNZC
aMeJP8OSgE/0LQcHmHJyK9ekH9f2cOAuiiswWcVjvCHt8+ZDSJx7zhOP3wWaJf4AD36rYF3E2L/Y
bO2gi1eXQ5P/6BKWN9ID6/k0DlKiC0GCLJ8L3hEKEQadtiTQw4URdDQfqhkgNe0B4MVaAGSLdzu6
X3ioNcQRRqJFrduxcsR/ADQKmxppV1pUoKpSSgzBjkHMLHqornsX3Y5OzAHHn8QP822rxH4DngP1
kzM5T9FnkGR4jdaOzuf0SpN+FHeOTp3G2X/hlOXjdzZ9YFhoOdVaeaDanJJctgt1hzWk2oO8WeXQ
l2zuUfvdjFuielbA88rrk5xd+qPFHmdE7S+UChZm0K6JyHtunOgIEK+t7q+sxWc0q7qP91+Ofe8d
ZyDqJ3I2xqgqQ3T2a7Ptd7Ml6ugIo7rUGpA+5qNWREPsLFilX7W0m4xsikLpU7im5FV+mxoqrm2X
ncl4CZaAW1xwo9GBRya1HmSnU56K7S4j/1/BNfhhGhaNgXYkooLkf0qCeZ3twbmrer9TQ1lqiG92
huWvyG0AFuQ7szhtnjIC/WYbwaIP1Vl1y590YS+ZaYL7J7rvcZJp5B8GTBFOH9yABj9ObhhcEeLK
uOtlBI6THaMZRqP4hatr8EA83UstenqJMZt7dZVIQa1lbd66eqU8Be53JhBe/fwPunF6kyfP8KBY
zp53Vq79/RKSUuKmr5Zq2kcMwxPSPk1QLattmxO8bvvB2K/g6EvjLNXjLMm/Y6A8zKEQBOBluT7J
Qok59X5Gv1fTabkyufeRBzaG3p/l/K7EiagNn1iaL61UjnnjFBbH84DDNXNdXQMZsv0tI3jyEjpq
uTnUHcd0cmI5U3ddvqPaqfMN3MgvxWB6I/1U5IEkgdpgc789DwhOxCeP7gFguKiUBFg+5DNSO/rD
dd/gXyrPLu6oypGW7RwOCNS9AUzAgZhY+uvmXRi5lhUZl7I9XpdTcQ0S7yI2T4r+vSxp4l22qfo8
uQXWAnrLTnK1qHC8W3Z28NANvX+7NicC0C7G6VDliInfPVIJ6sECR5ybJK78VADhC5GvZyicojPa
lVpGGpmZoKg5rA7peaU0bqrutBmkNGzepQ+e8kBhSvQQJ6wAXBFkC9Bx09Q2Pg2IXJnRO/xWGf6h
+L1Oy8q0Eq5QtGV6J1md3kE+aK8wtnztvgsT1605c2xk1oXut+QJ6MF378MvAjkRc+hxWhSdf+k6
naORQ9PkMNbpBzvjqsMwAL51v1PnieJeQdM+w3RGPVPPjuXmPjMSIwW44rPK3qbm0JnscDQ8p/+T
Y0+cTl5EMZ1aEZMbZKHBCu/W28q8t0ArBWRIWvQwqbN1BaN6CTycrbVdg3Fv/EpPXV8+v9fdiOmJ
5USla9rE9i/jZ616LQCVGjJk0S3Ajb7v0ZXvzvjgYKFd0Er+6VRes8prXyXiWh145GPvfkS0C+9+
qxgqWoQxGOz/2MAWk30yqVv0GkfodPQ+FiD4dyvWWnP4tiMrq9vaWlK1+ojUMBnOdbN5Dvw03Sch
xgp/19lUQq+2Xtk6dMbFqF8gcOR5Wdrte8MdnUXJclSfD998pc72NI3MNBWwkXhEnfRLBIj4+HMx
MbEcdeYkRBq1kFqVEljrTqtsCD7EdS9/CPpvTJ0CLp242AhSswOPNEW+JrMsKvi2jfgu45cPvwW1
y3+CJKAgR1kKd4cgHBL4ynCOnBGPJgp0D433D2GfhCi4CeYXUcm/rEsnW0OnOtNfOrXaXkO4Ldp+
2mphDnKWYi7VpAYQbU4ICZWte76g5U7BrKCaR5iYE2WiWUvHWdycb1mo9wK5f+uWyszWA3VN0PPO
UZyffPKqKEdiq0zb4ilCB7ACNayifLwwiPXVxFNaur6UjjYyRo2nTQE0Ov70Qj9PZec89pYPX8jy
VOLbhRuakKgVmsiduvPZmz1b9q7DK+LEmlUfQBUU8sWDouy00g4YeQ33+EA6WMHIZjsrREBEMyfF
+TdBfR+Pc74tigbCbf9hDeJTdjHjkwaY4MGMVGOEGS1XQb3SZttOSYlw/GJc81pb3yxBuNZ0bkWK
oqHOKwE8zbNNbEIt2vlLU8YzKbQ6RoKC5CfdWZ2AGLSqEfaUpTX8DbW3KPcJXLpVcFgegf4kSTmN
GrMtuKWZ8xTsHTyEGA8bhacUONBCjRrrQYbYr0Gmc5hp/bzjhnsccWoVLi4W2SBBVG3wYHORf0SW
cNvIT+sfX5t8bXQ8PfHk/kqZoc1DE+AUvdZS/BwdxhH9BhL64rEbJtpENXiPXdCzsURrCtn5KZCZ
mqoPzTeJOtgN+j6AtULojvN3EdYWbu6MaDrGw/q+3moG5bku8h+dRBtDzdqLlbiZ2fgV5hcPPP7x
jbZgR53o942F3bDExrRh5L3eCoFbXV0QMb3VOpENoHMpSiP0k9zLcdeyiv9R0JrUFhT9lf4HB9Rm
fAVpp8vLH2WtKb450iNW5AQdcYv+aR+PNNfYbwZJER0FyUugYMoPMetK7hXIuUTUrCTyRXico/nU
II7uclgVj7Ps5G6wGDeD9stY4OlFORmKe74/G7LBcMxXR7gR3MqdwndY+qyMrI0L3iY6lSVxscCP
zUb6QmekU8J3N4i2IB8vKXcJUolxTeT6wrr+sSkHMA2QEPFixVEVV7WHb3FmkNJX8eP8tWFSXFcc
aw6HIySWcjy8NyGOtzt6TsA0H/01HSvRn1Au/ETxjQDozNUjaNpU+jh28jFHUupG8bB4Mft3D6C5
TkPKv9ey1cEhnGGQr9LuwhWG3mK+6MekTzuMxrHBwIQn4ymIgzkR3cVGfGidtUlPxm2zsEKtFSjN
VcItwulAlPq4jP4k4aiXQIw8LMPFovOEE9hOaVQZ6x34LJbChBwvgbjWtxmeNmnEZI+1EGSHqdok
sVG/YcbpzQy9EQ6leEdVBifKcfJDIKUZwSe+2NXWozPBLYooIt6zbFYA4f28RhlbhJBiLTzSSQRm
FeL4+4dB1Ev4uk+as0IeD51ls1S9IgpA99ESUq6FvOP1tvmQ+UzUmLHZ0JMnHYw5NzH3j3q/WExq
SoPsWzgqwCvuDzzMsE4GEdCet1CDt9s0WpohBYxHseY9bhYyifpjwZCuxd9IejRYU5ZbKzJsGex2
A5QiaXuxseGzHFWSthAnuDZJNXPJdot97wAYhhm9/Qpk0mwWsG85K2TlVyx49Dz+KAvHxmLlCEeh
zj8UlvLLEnySOZyQOCILu/el78GvAlJ5ZVIN3kjs7M64MfGWHZWyyVAUVdY7Ycrp3SthlEEllmMh
Irgl4x2TnttaqkikY/87jkJAIm8GV53UmZyFI1T7BKTbuwSxgUoTFt/qR2iNUl73GVoy02kvlHw2
fOTrD1lglFw3+bjvRVnNrobL2lmOo7cZnjVWh8wiY/aQZ36JpBm4lPnrOlR/QV0BGcTwRpX7as5X
gFIM7JzMeTYGGFlCJ65aFNuJqvDAoHTe3CIo3hw6ZM/99HAr2VAVE2lF9zIve10UoNNDwqFJla9p
E7jDa3AwbWmEHZnTCnsfw/eM9rysSO119BYzjdMdciwXrdGNgpjAXlKNJeU1FgvpMz11MF42QNIo
FL3O2K68dnNFCeoLTAgzy3ljCcMWe2cVel2UFyM8aw5fdAlzFa86FEOLIlIHRWdNn1YnK2hvV3ga
3uL/refUtqH092bCuOnfbTAZzlCCDFeXPdV0kq+k5uMFomWoGMWYRdr9lzptvxclh6YfCFlsnTK3
g4+IxY0M9/n4MK0bbuAPtXc9EpCJh4klw82fFcQo3X0OlgDTyIHRK0TXpuyWG3LTuP9FJR8hJJq5
WDM7/7nvEocfYHbOrmxJnn+jFEFOZAJb87IUcazHZQTuCZunV6IWbVJqzrtXIVuVeGpkq6USsH2U
2Fw+t+oUh0hnCx1hFsOdtzr6SoaAdhMnXQV/0jMMmMAOu6fruuJFy+F86X/vosvOE0D4DdDZvo7w
97ulYNqjRO7ilWdz8emTE2xx8sgAdI8f0uKkxKbLFYDkN+WC4cE192MW/3++ZOXY22RQ6k0Vivco
FZVgLhFU7GZcaw7MIKIbz5f2EzIij8v6klLxUkzoU9nL+44Ua3f0gEMoNvolrOuE9Imz/a5et6eD
8RvkkKs0MtM6bVCFdmgnMIivf1sgZc9duan1ih7hgT/qYXAEMe/StVFfpPdYrPbB+9MYEqXwd+qp
zgTUZd4TzFoKmd4CWBsSJnA5rq8ITjh0i6boRuPmBRLNZjacaV9Yyxl3JhqT+DQS8pT/Tzk4HApf
PILJ9gXjaqrSBK0LLLZ1fUthhhbd2fvIR21fyGPobJGV7bJt930hDLO+E0iQcVk7gmNGWCSMGb2X
wD8DFynH0jLtS7MF7oP1wGzSsE+lna5VIA8pb0dPtn+C8m3xr+maC+MsCvJttq6YJutLL9rqRcuq
MtiMLDfx6wb8fyixQGBKI/mzkme2A0SrUA8qwq7ifVD+LmT+4wcFSjebvKr05zCFHyLAnRMXVN3H
if9u8HGbuiTZ8m3RRhSwO1oeIn4qv0M/CTkm2M+eR+D97wHuhzRIz3iRVfsDoYGc34LSD6+jcprv
MzA9tITDy9QAWvCJ1xTn0JfrDT+gk3DFB6ZPG0p4q4XM7Jy9Wq6HlScsUNiVd0nWCNPRqoRM0wVR
eRsGExTLVEqT/d9QJWyabzT+dB8Jg46uQqWIS1un04iNCmo51AjbT2ILYykqfchzrxyAZ2e0l7o1
/sjFd4lotZBl1XLf3tbZTyuxdYlJQFbw50w42uKsOFMtualo+Wkplrq3jMsfS0ELF8DOVP17onvq
TqRc/Bv5oFqonblIEmG6OzmUPf1EcA6vB5JzPoA6te7ROj+Sl4IDiBf6zgdoB/cEIIPaeOW392yz
TCzkGD/bzohji5GBTMCTScT8sQ7/CAB7BNryWo9CFfSls/LuFjbc4RhxrK5gz5TO1k78SB879WJk
XsnmWmrO4LwaDLxx7fwkWak6kFlPOHNR+cuckXuYnjWmTQB7FkTF4O4ev2MUy+vs+wVwMsosUvdC
9JpXDJW3FHnlt14mbU05g9kwtXtsqqp9B+JxioJuPV3oUXIIn3WTo51+HpBy6yNaulu0atCGATLc
JCwOm1gBREP6sawbdJNW6fupxafPTXc2Nju1YnHhVMOufPtsVTqvW5CNwQQQ2qqCytuXVX/pWmRm
PnuBiBZAQVYazrsSzl/dc48GB+OCGuAoVX1dusP7O7e49oojEKvN4kDRBkVnm44dAGwMa0QE2hI5
XElYVpg9+Unr1hMOnil+jFPBylGGy1lS0FjwRhePy2TmXk6FSKOEWiDz65jDcF6b9XhCiCFDNrkP
LPZoiaAdbCbwKP+0WJICyfhwyJk2Xx8rP+opVh35uoLGSnaWc4yYBMwMrmO0k0ZNrgiVR7ldSGj2
7kPvJQ7Nbm/6iYyCYNnH2LFbJTfyFebffrnun0Umx/p8t/qHmXxil4qnp56bN8ipKGnV2riKlPDX
dklcejLrR8EUA3+O8jQSeNf8ikmQ81Oh2xIzaNVmQ2DltJxDMlB1CGelcI4xHzshQn8MkUHh9jsp
fA9FkyWoD7rE/YrSlfAqYtX3VY/DKJ3QcTxFpfQmlWU9E6yLP/R31hordFQzNzJvmChX8YQL40y7
+Q+5Ijkna6PLgqw9KelSQdsAUM8nPYJzB3ruvfwQ3ojQt7zf43QGZt9PQ6VbnQId7Ky70VP0Xke/
yaliXl0fsDupWew9RVXHnVm2oNLNSCXj/aMh+4q1CG/1NHDd833TFppqnkzwdxvfqoSz2e2GQp+X
dZq3Fzpsy54sraoBTBmuZuMWeks+8ExlmCTYbrQ4+xLfNEz7PWaKB2u7rHD1c9SEYvYOWrw4lUVt
F40sFBOIetp1tUb0JQGBo1CUiWnqM7DHNiaZs4gaveMs2LEzsHdsY7yCi+U5PQfsk1WF1TmEpq4b
0Xqs+hgQg+6JADVVGl07mOIaNp716WjEIchpL1zETtUSx8pe8BR0kbGzI8n9BXS/6gZR5SYTLPbZ
DG6RWvwX+geXRETS3Z8L6SbRgHNoPjuulsGgqJyJqOXGOlZdpolFqgp+8z1Grpa0xilA6qdfLI2J
IiibWpU0INnMHHG/guWqxvyp70Fa62/YI/qBayeiNQLPNqH5dyTp4JZWXsFBja16AsKeBhx6T1rd
GuL7sUMCUjKaBViiyrmK25E7jtOoJ04wml0u0EdKamDcPbLi7ch+WRQuqk0mOXnZQX0/lIMCNeu7
CDzc+GFnnWiAdofyMBhF79fQPPzDPvkP0tU6guwZLzn7VcICNytvOjtcYJgIfDM7ejljSXdNi09j
N4ilhr0KZp+Qf0xs7mwc1jL0jr83V6OnN53QkpuLDYMBUp8Mr0sG4iL8XShcFnkoWyr7RILwWwa7
zs1FZaU6Axnp3hmp/1Cd7Qh5tczwiu4/Oost3Nh2pwYPMiE6v++ezqn/MjZNByLRjARAQDVVAiJf
NJKgoKwUwUGKWp6labrVENb+0E1KpaP88fci2G1Mwoxe5l3yW7Pc5ZKFrcjKzgTs7ifQsMBIc40H
pCu4M6HPTQ6XwNJLzAFkngpwTrnTWSBCGWrBDACQWXPxSjzgJaoCtwXjYEUaLEnQcyaj+LXeha5N
DYuxE2Xd8TK/CJbo4qCiQG1Hx5BcZ9dx4jv6cfAAYYqwD3aASzFj3Ww36gMioKqiprgeOPck0qZ6
8CS44SQrqBrQkwmrUy+QqlhL4tNeBL+cDSaeT3/4/ymVlsK2RMKGw+9kZpbXLfU33yXrE6m+AMyd
o/HlKFRss6EuuTp6E+ZNc9mNpJ/7iKCzZJ24h83LPscvY+xBOb/99DlhkOjAYDusKdvZgSLHp8kV
i85uo1H5MujJITPBVYnMCE1k3a5b68NxWUF5NTuxoiuJPhb2HeOxkAbbzL6wsEWdb8CA5Q1s+hj+
Wb9bD1ZaRvo1FGAm5NiLUKEbpFc73LxmKz1dwe93UNo/yCzwebKQf1fQa2iA1M9+pKzwb/klHpzY
7PYeKnG6jwKaek09uQDu3TJ+a3zpFLCxZyb0UxslCZscvJK+1FxX7w7loOFtYs+ZQIVD2X1pMEDA
9mCk3I8R7zKU9Orum7muXGB8XQvvH5KDXFRkZxzDycAgTUvNmEs9lcpiYv0Etvc2wbRj8OoKuQdB
DchrSqPzP/X9n6AnSnTRLl46AEMwihW2ZQZjbZgRYE230aVcG4u9r2hXkl1miXBcS04ueX7sDLrG
r5gtNY9EHpXeyZ4CW7QsYLJbuwh5SfkTOt7rCdIkZVDwsdxhlnseMb0FZFivFxhdqvOx4yd4muak
CecPS6kPOOqDKHtzYzR0T2c61dGoq0cX/x8aDveAP/BJjK4fgkHcBXkE08/GKuiIgezoq2TVlLT8
EZdKc4DpTp/NaSf9c6UU+zqOw1D0IFq5aX+1sBHUaAwfS3Ap0UeLisy4ytamu/Yk5DwqLHfjkHnk
44MHArw1kTCW9LqGGHmeCLhOhYbCoIL2lUED3H2gaO69MLjT0E+2hXeF2uv1rkV035HQXexvgmG9
G+FpC3LqLpirm00X0YrPTigs4bJy4OFTxJVguYliDCwf1ei8g5Vw5HIwa11ADbH9JfuBjtwTBAMH
B9xXWFrTb9c9TDwSiBKPSgUb6qWQzyoJ7yQYqSQwkRQo0BKFvsl8DooFBBIPuQE0WSqwotPHmK6Z
SZfU6IuN0oFkcg2L79VmjU3FiMVv3KaAV61z3/3kdIS/+dTcw255CRYznoWPoqRopsZo4RZv7MvX
P8FtkDOcRLq/+FAKlz0Xebd8M/haU+q2nAXT7UsyxKIuNbslVg/x7vzdwdubhIKaA4EaF4XnIvpp
rRjs6/MlitKNJelmZ90YhuRSwDTGP0+UJmXnUoUGvGJVnLosXM3xpjJHnwCSQN5Ftyt+x+GgIdpc
CSnQt9RikFp6Pt6vQraqblOP06ZLjiB1wZ9Yd/WlmLPCAHwFXUec2hBHikEL9KWNwPZW20HvseBM
iDXS4XWdW6Y9ZNdniE/hnDYxgJ8m6ITUoIApEQy2XShm9HR6lhGkv4PDCmLYlHU1pmHLs4qdTdnl
svTGigTBl5yfesyZ0jXQss62Z4jVEfhRJ0DVxJ7bkIYFoDc8MDAJxcCQzf6oja86mX6aILy0sNWH
YQPLKlvSD09PoLE1dM85MjSV2Ll4RDzYol968OLol51CiLWqhMGaLMtF/oq1Y+2YHenoI7u1OKi3
504yACTLZtOHoEi7Ei5v7Q2eyjWTvKhoIfzMeEsREirgRilOGGvNdj591OtR1oUwVRFnUG9/f8eZ
HVuh4wpzHtMC0gLlAN30kIg9Ssct24QdBtxeIgIyLUnhaMKiOV944N1SaWfmE/H7G08iSEOSgDTo
Vu6cgsskRzhoCQaFmcbzZ+Hc1U1qupC2NwKK+2cxFWMZFqoS0YhHgN2nufWOy6yXGSIaE+gOFwQN
jmQhv6h2fURM8Hcr4cypjfOexrS36RGCcLDhennSfIBWwuvIahQ9L6q2WFRV1J6W2UDji5yWQKPJ
UtlVAjUiiIH0bJFrXv4IToTMunJTUZYDbI9T6EpLv2m7qJVT8uZSTmUVmW1BddjsE8xzuMlYGlXr
0gFPsUCzQF3W92s73/37yYLUCI9IvK8DswHO8M58Hi9W765EOyRYcLRuLBuQQ9VXsZE97knC+58o
BDPlxXqTyrz2Gt6TNKg8W9sGnyZNKw44n8gbqrR5Qmk31CCbs3v7QVUYmxEZ9lRwzGszYKsDLXJA
/ONCwAnnc/zeY4be8KqKxUICNrJaV/nrR3QaubPoM++snrea1NwCPV4IyvTLs3wT+IR59Dn5NMVu
F6LlgXXebK0LKCFqe6Adaxxl2Gvwb7uH+y0YdRBRbKuUdOhjSyOJ2lTq5OY/SEXk+v420qbBtmDK
ptoATC6K4c9gUia/3hCbf0ggPZabKX7Prf35HXUjKOeDKvt4qfJNxr36zMCwiJqU/NhIcOmyMzTo
2r3YaHBDNKv1BuPU6uM/dpdaDV074AtIHsr7q23X5oxqLwjCbSz8AIblpgcMrVgBUUM66XP8/VJ7
dhTJXMSK6AD27yN3hD/QdTDOy8BEoP23Zr41cucTiRZ5vW3Gced6CMPbdmyecgAb86//aRzygtjM
gw1uDss1tgtRtm/r+M8H6/hBp7q95R8nSURW11ttIOYbqwPx5sFtrE82Ncbh795YlCIoQEfMiA77
GsB7MQ09/H/RL44+zXK5s8lvljsvldecijwZM28l1vLe7v7zy+eefqTMkcSiltN2qEZQGSFzWjiT
b+5JLpi9L80QITR3WYXMj9l4fllhYyqf7DOD+1DizlDKVLI5Evz6/Pe18gB3eUUC+u2yc18ay4ph
vFOYQy5azXEUYxuqaH48XlTTqrK5sqUqznCqEVtm85vqMDjcMzrbIG2g0oteQvhBgaaFFf3y+0Ih
LUnXx1koItzFaku3EPFam8ecvBI1qr1dw7apOakITPbhMDHOc9YaKB5Kalp1ApIZGdw+9/m2GT3t
m1IutVOBUPQKhmUZNk1We0I3CjcKwL0bkVRL6hKhDjP8BtUQoz0Uv0S/wRkqUtGoK3Va2G4K27Yf
5TDVAG/anFed84V4s/2xy5YFSLkQutCfGUFgE6zRIQnU/OZxHLo6jKIgw2DldgA41WYcfW4+6xSc
svebu/h3nTnaiJAvK2vURXWFzWbEzEBudg31XuWAgpRqgOsz6qEAjeOZDrnUsXxJUob66Fo1Gye5
hoFEJI+rzMkOT4dSeYDfCkBmP8vEmxg9Kl39fIK8DUdYC4OSmpBIRjz1e9H1JHYI7Ekcirol91fC
aX3GLs/CYqFlaqGJRQrfiwtre+PmD5Krl5c1/dJngTry0ym10D0Osfw4rNMn1gGbKlOV4Afa2fO3
pMspQgmXa5/QzQU2aTc8KQXUYcR2wGsqfh4X80Mj7kNSDUuvKOTcvNbWtkDEI5acGYyBnO6YVqCe
rXgl6T06f72wez4CRDnZal1prcRlGQljaE922mleEcSF+R0wMAIj1zuY6+48Z422cZ39WZzdaw/Y
roRZMcL22X3ZHyRzrNRumwJ8NDfqpORs7VHk71w5bsefyFR6Q8FYAtZPGEF0Galn+ZF9grC9Np74
swsuCxfWFQlrOKVV7S8xKcpGRYo6iFYF4WbVONdgsKT5/ogalZCUgxFQAgQztS/lQmn80qQekjlD
aamOoTxDDsPO/YyI0wfGCNFwBTEvTAZ0qMa2zzK2ksPZqgbV5nzqfJPvxxQoBucgwb+3aCalGZeP
5R8DeGANFv3UCUwWt0ONVmB8PSXM6rC5M3/rxUR7wJAumJz2pRzeiyFHFElz2DGSNu1kTpp/aw4K
NpfW61XKZcTa6Qw5jAmZp8e5tZXEmzmbeAyqTZuxLePdqRAFl/9NfT5zNnONMke6BaWCcO94XyFt
w5rnLBbNh9QrLcYMIbwbT03EE2s6wiMmo0ZoNOTLI9eKdgElngy0KQ/ToAHk01mOfwTBMvbiVG0o
pzBChDktPRQ7ufNgf71hpzmXzdEX6yKmoPVC9FZDKw1wU87CBmYTaRx7TYLUwAjbvhdcL36aWMKI
0PL9y1o6TH+l63Al3PBdMndQQrsfuw9gZlVL34EYyYempz+lvspjppNeAq+kUVNhquyS12W421pE
mMlNbmxNhCRc945v7Ahv/M9VDMz25ap16FlqUOlMvHwMgIltEKDXpLktPDSb+kLNz/c3l7EdRgYV
zb46qb2C/jUMKKNl83BoxFKOYYQg1vBTe8kC+/X3APULYQxBWQOlkB/I4gmlnMp49F3prP0z17OZ
+VtnyntteadCfuALVWqnUzK4aWmxlhTHMkWByqyiua1YNdPutvSxaVOHCGtedTdsHAT4RM2zt9rv
4g6AILKCk7lKDnFmy20yM5SUbfelOsJyCnGhP9dDuVxNAz3503SgF+DN4kn6hFNSVawkcNNbYyO4
XdWXSIbiFn3Iko8W1OHiqQT7ygEXOwJLEITd4QKSn0Ly94iNE+H+/Y0bJEGioM5FXPXq7LASrRlv
TFEVFiTIn3n7pbK7/65rIUc4MfxT+M4mcvfJkJz4p7JOA9APhyLE0wa+E2zTJB+oWppHQvsk3eux
+Tp/gspRkB2cnfHlAkHVpPT3uUEvmOheDsgpvo7p+WvQBinMIN1N+ccc+HAWkMbR9IU2K+Y3JRF8
DRx9h6pDjUHfXMfpDUt69m3gLrck8cvVka2YVWUx477pTNEmSWpH8JhApCiK4T9cqfuoYbd2NRNU
MNbq4Ap5g0uPs/8odCLMQRRlk87aP3DivrSyhICf7pd0yTjzTPOTi1+0HWxfRw1fUqlBag27ySe/
FRR3xnFu9cyqQmCdtegIELujnYP4/ieJe+wXfO/zMJLJ3arIVXScid25Ev23MrVD9TeCdNESpWGU
oUJjFc/vKVoeQqbm5gDmj8Xecq6leBO5t6bnPM50rQSNJZ+cvP4Mv1HGWDCC8yc3K0GzIVZFxoQF
2JYXvKSgIrH04FSYM29rhdWKMbDax5Zu1hm0PpLM/Eyila8H/UQ4ONbTaXesF1rbd+vuhKMVVOYH
rKITJZTb7MNicRmbHINS1wgwsfbq6KssXwV8up7AkpwasyoLXFRxx5zmKPAPuw2Zcl3DmOjpMaZo
14tHYLzvQvELeox59UN9Jvh92jwwilGViBIIuWVc5D6qLwZ59UyOfMPs8r84yIqE6++JFrrOYClq
Gu7t1arUreI69yPGYHRdVbrczdaxG+LvKGhZbWf9xYRoe5TJ3wjGuSiGqXtnLrqNGq2ittuch7L/
9ORb6J34I6grx3zf2bC7PbdlQyUR2pjKarUmowaUTarYlG96wuHL/T6mc3h4E7Gq3YBbyxeLx1Cw
QFtiSn4F0aPZJ90ka+65iIPosspU4aBbJkjRwur3MuDSClvwbjmTNGb/wRUHD1nupQuNpEfBRkEi
rdbF0NLH9RHpTcCUZ0jJQE8TIzdAvCnJ47tor2V7Z7gc92WkWFx01Yi39Xijh/OQNcb3m6pY4rvY
6tl/70oNaDCwIPIcV106SQY9LtD9GSoEVsT59xcQO0MUx8xgZvUQz6vbgS+fTL5NnHdeDG0UK5Du
3I7OeXCXjKEu48N5cCE6Ifo9MZ8xbOFauYC84YweGhR5S02RiUVvwD10cmFFUAEUAFS2bqAgHyNZ
THfiSvBsj30IpA17gZWupqBPx0pVhdHKpdH3RwwQ/Zoo+dfdfDebHUwS4XJ+5CkFDwfIBLDrnZnd
KmwB063BU2lneYdKW10WLGBhU2SmzhzbV6e+x6ZHCT3LaX66jpi4rkX2LQdncpdGZLLkFAAVr1+d
/VCXOcVIvoZ9NgrHgQHZuJcSy6uNW8S4n4M+Jie/LySz/kjMRx+6Jsz/XSHGyq5e4k37HjwLv++/
dI4nfe0NzoyIDPW2LVqSfLHszr6iugIeUJVFagQzWLzuISCivGu2ZMdudP7KF34H48fmqVlEdWPx
F/OEtLkjFnD/bG9jFGCqa91Ilnus3DpGbYRWPHIP/lFNCQOXDQzLPPZNBj5jaAbO7asAcQ437m1V
akXXuQ2TOTAY/g/uW929ECNw0andoiYh+1riKme5BSf5vTIU3lPUNG7EVkhqZm0MmOGS44kHffu4
aWbyv2BwvBk6SBRhHWiFjv+D7odaq6ZB40iPQuP3P5LAtvMLev2+1zymI5MpXZOm7/qvjIGk1HKC
SzmbRUd1qDhlo8jmHPhdZX/XhUJPahXEkDQfgBditCmXG34bATZNXMkv1Zjp+Lq1A6ZSB908zm0N
39n6RQ9umrAUig7R13TgG4YNNFHbygSFGeUimcl1chMxEZbU+RRyMe5PxhVhJFcROgOs9g/Ai3vw
5qcga9Vc+pa1lC3hS3gWV9Bj7LM+DMAuNZXP0XKBR+VcBRJiHR3pNgn6sJ5IFeV3OLj6f6IXIftT
GWrRVOd0SXFwnHPWfQZba/BtGJWpdRbbZI4g3Nwn0nHNoC79iJiF6IVDBITYyWJNEtUe3aLcCiIh
ufYqbFaSm8DTZFqsLo7btjii29LVZW9dpzy7VX3fleGAPfrtpq1eG1urEwu5rsrS6z2ChEgFYElf
K1pNjouj9cDITNE0iObXiZvDaaQqZlXIdIRdjQgmiJhCWJTVyKEI0S58tRdGQpxsFUZud/1NvytN
WOgmg9oDcwY6NAJbnJ4SdW35EKmYpp91IC7HzT5cj28vzr2tjwW9i0NcNWxS2TyJOnPfKXf14+7c
aPWiBoP0VkE1pdORwCbrYqct8zv8vHtlubwov7+zIWqYQlV5cifVFV2cjMeY/J5yjP/VktBvyCdj
ecdVK6KZiFzD592kxA1BWdC1Xb7vcC958LLygTga60GwhmBc/gGYFpVufSGKWL4bLhRFjhwjwTN6
vsoIqr9V7DCvg2f+YT/EeJRdo1MLgBv/ZZz6F9Stlw02KRzvlvkMUso3bGZtvZtlUQs7bioHdkJ/
5UuunjsEgYsQgJqIYFJ3xUABWIEWLNYWj6Q6efA7Yu5mOp/B60GF7UIWhrJSC8o3V8avd4mBhYl8
7/93tJgPwSQq5vMBlDVpI8qcP2AY++QtB6MVoVMmDMU2ACwLntEPBl8wH7HQoD9M0guFeqdbMXjg
aYQ4rRPAEocquPwIn9W44Uic8pzxyPyYdaXA1FOuAvEGFErbWagXs952jHc0Ro9DFiICQsdsMmav
MSbiie/x0L5ijie/hwwuj6eMJb/HxnducLLePOainhRwd4+RVzfjHl4CtzdqWW7OpqkqAbGqYtmI
eN+2Y14KXkyboNYnXoTzqtnrKHC+z/dc6l1AeVyja5VmG7KQuVak+LJwmrlFHz1rC8k0XzLntSVv
F1UvCTFfTAR5Zz7wIaAGCtyNqnyaNmt30lSum2/b6bTO1xkAHyY1vunlWCX1v11KL6ZEf5nmN3+S
79n973AH0M56K4W9RqZRy0S56mYSzG+xv+lZtkR22bI1wuYixIU8vgO0UdTP1ZE/sdG7E4RB8rDA
M8Yg6Mg9e57t1rUJ2ieJNlueDuJUWQaDaNACNE3SIcvLtU2AF4ozaClHOs8wWUJ4RIjKjSl7xtAF
Xqem63ZNGNeIcxp0mD6IkerUTOJV+de/Dmd5hTGqCz6aNDHiAB7eRgb5QjT8GyupTTPv4CsamgTE
kZlbhq+4OStvqEOO1Vyx4E2vGnKCgdxdbXXpMta7A8Oj1KOmdXDpqIs4BKcPwbBBWAM3516qHOPK
DvbVRWBvwnE2q6HXMOreOzwe3BdX20kZplflbf3MGYB+2/bRcRZIYmktba3WWRgYZJlmvFDNtpNX
Ay/rgUURmcKYvRc1YD7GSvU5XmmccNrdDCRKECYDl2kYxr0RDF8ib/yK9RI1vtdXR1qhYEtX9PEm
2zXYBYMcQNl7RlaS8R3myFisQasBecyJqPoYF0mcwuzrXQJZqzEgGO+MMgxL35GGma3sQGefy4/L
ui+vKPqgLd0ALANAjLGXV2LPLrdIwFKEgeDnt/bTQfFlFyDwxwqmnx6TS/JI0IlbZRWVQTz9JTlc
obKFjIToWvc8uIWgc398w8sQ5JglkQyxy7nOLDwX7UjExU01b8fHxsFtRyhW0JopdSwDILwynD/p
FM+g2lbpOkNoHnFELoOtfWcDck1TDehKym4BVu/cUOWclplnrluAfDzFUZECBwWLX8yRTz6ymNRc
XVo/miZ+o+Ws4KE/ITZg9KAyv87jf78wvjIIxDsSIeHieu7kaUm0PCGLmCEpk7CRU32UirANmens
EqJincawxvvfCdxrz/b1de/BMPSNJejH7i8m7ey2p94T/GgMQbsxVLhKfXyNxbLzHHaRD2jbbDUx
/LOMThi8QbQAFiVgje/72Oom0RJHvQ/U5Y8YTd/WV21mZiVwYiL+PGllLzo51Nwr9Pq+wt8XEobd
1f/jSzZBzws9f3+pXVM8NHnC8JVbX+QJm8GmsQsiJTxkIJbPsKd2maTZiR8bFy9P1D9eMAlpllI5
+ya3bkZ9y4zhOl/3SfBmrliy64+4cYhUlnxVkcf0Ygb2zx+YMH14xsrQjSShZEdX6mkOH465y3mw
cliAm12UOatE4cKTc5YFDaC+NOm9NBtA7O7j9a14ni3inApom4ven3f39eYIb+NXDu0YBdXBEYOF
vmtZtLIovlmHjwyLDoar7ZJYXgJA+F/U+6u14rsshsydcqtX/blb7opPxplANVn7gf43ctrRRvZm
xDJQ79MRU/qIOryDGIMPNQ8MUGWcoDDpgtfU6cSWGMAwXdpp3eU/dlh1fCUJ829zpjfySOE+yBcs
D8AxET4kfmx6b8jKKX1yX9vUDLQ7HnFdrWrg5/MfoD96y1yKmx822nmydh4pNXHMVZoQRy30xUWA
UwB6UTL4jpi0ejQXgtlzz0p4821AOLdoycje5IXTXqoWsSO/Vb22D6kA/o4I37R1u8fXlB+BqD4a
oNoXUjWhbCj72OrSRwzdmPChz0bRNMLusG85FWdOn3Wu+pXe7Zh7MctXlR8VGQuxtsoEGhpMnKx1
MGtzIf0esF5hMxUpRKz2Aj3eXlqINHqiH9BcQsbfljTkITFsHjvxsoMrVgThfV8Ni3bZFiVM49de
fBdRgFHGMaPqHvy6iV8G21uNYb09VjkmLk1OaQ6Lpqdw/orbiBEcPorqv3EI9s8ZvvIV3ATpG8Jp
2TV18FZ/SKHnlt8/Vn9E6Nn9Y/fLL5yFjroCkG6qHXHhlq2fuKGL4AXBnydf+ZUehjnHHS581Svz
zcX+yIzbIYmtIDpHipqEriAiPeyt3pS9Bwmg/2ePmYyF1k+IppeIIgm1nqbU7OWMKNo7T8e84+Nm
mRuaNLVcH8ggafCu/hY/Ux6z8srY96eP+RDAjV4X0KYKdSY1kExOXoiTv8XMxZDYgnUVouJ4bPQn
ng6PJt4hnOkAeHxbd1wvexmWge0qgPjPSYgX1X273cOEmG1etZb+6KkyUIFwHSyOFRej4vG0PnpR
B5i11c+LVeli8A5tqF4C7CuhIWCIKbvGaR7aQjsW03q2imyGuozXv+xIhGH5oUeJEkJnc5p4+65f
2pLZZ15rKENg3gSnoQ9mzpCkObZKswFHmf4NT/E5MQ+vH7XKFeAKO8gYOjCkxbMnWHSqTIf46PCf
JDiLTyjaqVxeTbw1SmzGzmQPWQlXyAPdH/KWTikkWjRGQ2upj6MMpiCK4HXMaNIg4z9B4bTbHqwv
YqyBKIkHFCZUumcaWkH6vsNd1SP5uZG0s3755iFEiIjGiVYfTmqu73GMwXjpounK5nrFztweZ7O8
w68eh94JS0q0jRrm7zbS5yvY8CzbdqurRFvQFLqq0wMBhT8Eey+wS8b8HwISGUtucRyXOYblzACw
9i64QGRvsGS1vVqJtshj9eThwKuXdCBShSD8RFCGjyZtKWmUlKO1DVyiDFrlVbxwKPeaJqzphvPj
0Sh56egWOI+LQRV6KhxLyqBTW+ln12y2BWWNsNtJSAQrk5uuQQdxER7AgdXLnwY0zeCNT6Vpakrh
RGSJpd63fccLP/41w9aWxWHVek3hutgHNbLfg3LI4MYzFPyY6Z95ymYX7hfvWDy8M+PzGpne7WPn
bcPH5G0jbbNzk7tVy0dgjkJWR6yXjr9jlHoTD5EzVL1LpOv1lzbrzppnY3y7A/bQyLyh+Ci9zCkg
4AEBHhxBOcR4i9lG/HS126xgmJIb/AlyeRncNElpHdb9gAPriV5qdfQpQrbu+T3X6b1iKn52E94Y
bGDrAXR5SyR+m/ffNciVh45n7L5XOCRyFA5zA/bUEc6FfdJ2yy+ookYYRNgoW4VariP+fCTMf0ob
AnTZWp9CV1C2twwVYwtLK6F4pBPj43JVugN8QCo3d1WTJsQ9pJ/xbt49mlN0yPetaeOIl9P1yo0W
T/BxMi/I1hjdEETD4e0zj6RdECjbX1Z4Nw8stnki+chia21Q+iooJ3P3/L/Po1jdWLFCmM3qK1sP
ytJMXrXRiStYQk1BSJDdWd/nvABC1aR06uB/RwjEcMgzZ7HV/FcNlawc47n9ENUtkzo0b32hOunH
Vn0CQIZvXGKJF987o19J7uJD4Lk6VufxIig04TxkwefyAktgkVccrR9/f6iLoyEIjdUtRjoBbxU7
RFqOSD7SN0Q/RqjC9mNx3WNBJMrVuzkHVOLNAyiX12FVg1R1mtFWxDiJqRNmPemre7dl1M10MdGo
fhuGlO9u46VmFLcgnzl7Y555DvfPhLxZTAmcRSQA/7K4gvxUPzN4dIu51OepwIpvotHJz6jdc379
Ww6Oi0N0PyoBPGOBNGyu1msfVKWKALFOQTGYnIIRPKUhKszc/5EYrVZv7TOuPlAvcKYiwJv8sfcR
Cd82B99xODnTdg4BgJo1VpQB9JuYzUMUYZ8qmWN4cHc78nUrEqy3kLBKPGX9sxbXegemfqQ/zHJM
7j9IxOjmeI1RR9GZhSFmhyTUiy9xc9PKcc0/0yNmd852TLosi+PZEp/kDabHp5350l15+P5Mdmb5
++4rB+0e0XQLXyoqbTy+yZAfeL9J3+aMFaGeG7GmpLo9s4e/WMtP4BBnPZPXnI3NWF0OMREYNDsl
nZxu9bB+LWR7cT4bAg4GVBjp2lxGX/cP9suOHleNjBgTIx7sBF5nECLwommQpWAnR0ST3fKls+wu
SJDFhANWLkjmfaq1pmpI1KWzyhGmUjgSvLno6q7+lYXdilzTEuOwwD9ReTcL8bJ0q4Qp0AulK+rn
AENMHFPhvT17y34UsUixyJydofyEo81Z/UpMVpH21MFASmq5NaNFVhnvz0rY+Ma60KB9J3IBn89a
dTHqA6jgfE3+6g97AwXbE95yuSvK4Yg3PVnueao50pb2D6+58ORmlez3ejQ6P6j3xmuVlE4F2HoQ
cohNmpWOVgErAv67S2ATJs58Ys59OY6JCNp2dAuTdrXyqg60qNBHLPH8hU/7xsVPAOZEuVt3YIlN
fX8zlPSerOsfh8biqpSaU/CLCjcP3I9Cv+jGdhK02dql4g3+Aejq1u9bDYOOLzJ7NPg1SPQoZSV1
2AGhf+4PgcmKhkRpgWC4q92vT6L9TBKw/+NqVw8a+2AWgvOflTzF2tcLrPXx9K2AS61xqRvt1p7t
4BjZXrRACwrUC0aoYQuvaU4rgnkssEBhlUqaP6iXgzKsZslkyUbLAl2RGJbGBseyo2Jo433skIJT
6Y4S6dBBb+g45KRP+KAld9r+8jnvxnakmhVC4+93QqQrqfLwPwg3kYYUgCnFP+2XgsrsIXcGpyFk
Vb3kBSFRKK25xX9L6+XxrN0Fy6rn0ifgwoSS98Jvki9sXdgEbG7924yXA+diCN7GeuT+Jfd8msel
y+2uCGWmMQPDZmQljacEG17eFSy3cxJnvsIOoJaJc24rCAqB/fT3mU6F43DrMcMC8uVqygWrTajv
OTW8eqjkNeQtdcXrVDJicw/d6IRi5sELdV+4hAV029Ky9okMsgvfHmdysl9WBUJsYvEsys+WdurC
bVfRB3t5OWKyi67XJgYr9oS1Es49pI6mT9X+gNdLVn7oCK9NyyiOBkZANBQU5jC/OsI5TI8dKqYY
giq1zhX5dMHyUgnfKDB24oH2XL5a1oyqE0KLbniTAjGDAlQGBBAe9WM66Kv3xV/dkjjLqAdq/SuI
9q+x5YtnNMzHP7UAfeTmSokK9q2YUtlF/puPIQHLxQWdR5g/FvJqdXyDrVZFPV5+1IvzZa3KGwJh
NwHjfv7nwp95X1jXYVdeH2XWRDpPRAqavFxCbHvRfALhEcNvMjCRhDY9Np6VByp9UULBC2VMyOZf
E3ziTio66XoDG0Q+rMP8QCWaua/Ed7yTVxQvh84F7T2AJI5AtgWcTdBF4OZRYPXZkJzt0zk562Tg
nizYuokNIalZkrNyay+zdoU64Gjq1Juxk2UijA7myGYXGWUoMbIbBvJNra279E5cWwhFwReXzjYV
/MTXHrBIo4qGUrEpNRGLi+jqB1Zlu1ygv8UjpD3hpb8jruN7y2/hJ4L7FBIrOLqVBS3UUVrHs4PU
Vf2M8ZexbusMNovM+swgJApn6epgMnARLpz+Z4ZsY3ckBMgpp0ybbiPoZBIdg92EtOp6ZhHd/6Kw
lEOleoTcGCovu/YC4MMLNQZioHxy4cq/pKz6mFM2KxNc4IxOw1TegjwkR9JJeB3lmnEtUevgU/N9
lUnYwGRvQPnCAv6yng+ThXfrts9hTAgtkuHnnextqoK1kYXO9gWo5J44wl+ApVm4iHmoP2ip3cwB
S2eqdjEnqaIixXhLYGwg0cT3UGdfLvS2p02cQf2TQoUOzSlFQwzwYooGGsUZ4FFLej7BvZgx8cOh
ni4k5vlJgdxgxOcKPfLnrrtWqonJ7OFLWE+g37ei8p3XQM4waBdeiJ0jEcQ8Ga0E8k5IrJX6tgjG
7TN7fA0jRzElOafnDErEC7J2bSC/a+RnBWtG7zR7+HVXR61TSuEa/+znAzwlwTg3B8tR8O60s1Z1
+kx85KaEKjNqLyUI4t1rdnKJLHXzuMJ1QSwgiKk8T7jwwPH2+gedBKXX7teT090+C3Qai+h1wExB
UESlLRCCsorZarzPnpvA5VtH6Ar4kMoXZ9GZdIG+sr6oiUdrieQJH0RHUVBHC2LVmGlhJAd9qvRI
HEVZ0AAmsjKRn0/1IsmVN5TdA/lWrXLUUoxSmX4hP0beoQ7WwPo+Azp68A9FZckAWFoi8yk1yxJ/
5dyZ47+qLaDy3x4k4iqC92kHZCWn5O/k69fCXHU5jsC9U4182yPXkg18W22enCqhaplFm4SRjUe3
5fTHYYg5NHO9b6TVAtm+j/GeBnON9ONbYDQfYqMw072to1nyNaj9Gyt31zcnNj2uluhZdr7IhaXQ
KgSOfb/rlaJCY/YaM3p4dSMhORsRa9BaVqolath9Ba7W1gpfm2sZ/6MXXAUyGspyBNHRkhX3t01+
VxUOb/+4pgxtEI8G/HX5B9cAxxvr+rIgBi6n0mi8YiRfqtZzLolpN7nqxofzIILE2HI11LodgbZE
jODZBgWlwBIYxqOPzERb6nGmkkehlmnqbdC/NjMfltl0wCE4rks/Vzlggxs2eIvuSfGWHRDPikUg
76sQdGxt7LR2ITYvYsKV8zpMioji0ncqjZ1T0zcMR3rid6xqSfo1OThH8Ycfcf/fQAAk56zRLVxg
8TBVPlpgIYJr60GaR51ZAal0FYs4dknEoA4p8KIW73NG+ce3zi38FJybSibQFllYGmzamhmpR200
zgQ+l8xRUGZe1rOWoUkhB4vH9Uof8J3sSYY9HVHjvybHvithipBYyjjxaC4islJBZ2giILxIjJBu
7ZZk3+s1QiFfZwdfYCXNt0eydkoP6wxdPXJRP/fanhkqBqZ6FaqDTSyRPeZlWhVCrXhXuxnWvx24
SJnIknMJBHM099BWIY/R1n8h/crrLgYs04Z4xcAoSf0/KNZoAAMN0rNDrga4X/Qvx/TN9V0j1+98
vQ2RPDFecp5pJB7TrtEmvlC1KAiF7Q+NXLbZ6yvAMC8h5RK9PE7i+xMmYl6etS8haOxNBaiH1R31
en4hU/XM8uP3G4KsNvvtmS369uoZTQV+SgDMcWyRVGJwQPkcjikBQX8VnIii6qk+Bl16mEfnN2xk
0/m1UW7EpdeD5i6MNn2faGoY3FXlS6+4vRb3oW8j869LwmEDQyVulz65pYakA5GVQlqubr9dXGM8
nX3ajh0HY+sTXtiPCkh+wWEcJ86i5epPrN5m9XG+7/xq/HtLRyuJ4RM15OgP7yP3IU/WcEvP/MzF
he1QmNHiT10sgKNz+Bld+SJZoeYewQt0PM0txVJG0p9wj0nmLSId/JhyrBnQkQH575qLrtDFUvnQ
DOWHn9kYyf+CFZMxENGl8bFSd0NvkiFEUgeCSlSEmR6OwBuf23/4oGmclw5vw5DwhyZL3FflFPYD
0fButK8gZV0HGCshnx9ev4nVewzCu9qJvGoU9sckyTog0wB7SLnfAsKfpdzW+32noD4lZ85F+3rf
N2GVH7kCOnrb1Fb58+sQwbVKoycmcZjPne75aSV+0EBbRMFMY7s8W1+ZDGZ4zLzMPZsMaBM8Ui2W
9SyZ3zu/RuCN8OzbJWuiA4uKll5i7CUDjHyME3lqfvIdGsnsgEJ58Hqtxo7PyBeVXdYVJe14bjXG
Oj8zD8KI5u+8uMghgEPWF+7Vra9UAPjbX0AwEbRhV+61Mzju4HjwqvEIQY/wm97JP7Yn7JCDC+o2
SJoe9NSuHLckEnn48q1lrkbOTV9sVWL6yVO1dARviVbX8f3lh2U0aX+nuSqS3u3V7PAbqn/FASn2
ywXXyBzD9hBiIBgzUIQHDFT8HAPL+6paznFQtX0oseepPYv6TCfQgHLI9OZfJ1499f+56y5i7W7Q
H05ueu330qWDaMkN6cFrvEY5wBVVl03sc8y7VzPXv32+3TIDQwJNwyyEHdtSMIpBTOidJkqZG4md
8WSaOGPHcEPxRm6th6TmvA49Q+/NkRNwuMiHQeyvRPbjspkAt2L7Xh686oURukvvq0At+iPS8tMo
QCllpH/FINBaWfha7UwRXnp7HQyiMX2ZP6ciwBJZeNV/OiRL7sHyQfUhV3cV9Rw6VOsCIUU/7qTX
agi3y32lrZRKgvIowCKaMbrtwmLOWuo+Hrj9kRmactzz/RU7N6kWrLrxzdlvNglTv5pSWBCp0JgM
zvsQjPk+25XqQgcnYnIMNqDXqX6ArJpRxvUllnU3aoYbWsLwfyPOBVNkzodspdcYC+3LlxsF0khr
JFEEQ0VxKS5uVs6R+fobjOQZCTIYcaIWRdWBEuwwiGUNIqEYjOtAK8wP48fM+C6k5/pPsXLag473
H9zq6slQtHJ8TeIl6Dsj3dCmd6BcVIbPfSQq62l7X/eC//nKAKuf963u9rOJT8zF98UKFYqa810k
/pVap8dY/1hgax5g3tkuJW7Jrxb1CfhBkVOlEw+JwrzK6Xr25H69fAkcFBFu63Di854Ahgx8exvc
P6bGc8MmgPVR2ME3GibREai4RAzwC7cKEF/w2ssa/YCzh790n19LPGejeY+svCDSCO5Z14G1e5wD
6dnzPYG1uIeZrYcKcDOSShV37jMbfCG/lI9GM9XWDSCpwnDJlez3GEM3h/PqUWfF1yLIMHm4wKqr
EMXybPFy8+fFo0IR5P7FT40ZEw8DOSyKKTX5HKR1nD/+blHEKFyBd+FN4IsS75B2p8heA3TTIuRJ
6uvRJeDs8PriE2s9S7qS2/OrqBN15rUaIvMegom6EWKDyeMetcE/HnuOD/aYzKIjDwLpcI9sd7Cn
JU6tplaPoocdOv0e4A9sbk8n8k3TZHsJkO4GjT2g4e0+Mp+AbTkjyt1KHhlic1qx07Sj/CFWpOQ3
PdhRiIZtvo/jNufy8fns7+Z+iQnSLLGaEQQRcohv3LZy6TKJpjCEv68gPBY6JokUIZGkoYjgVf0U
nBTPneh9KkVSk46ONKRXPfTV1qnmvnPuxoehDvfxxzoKSeMet0sOAksFLiYDJRhS9sr1oi0VI7gK
57uHqILrnIQ7eiNUSVo1iRVLJzTzjg8mJGa04jiu4D1+WYyUMbf9A8qKYM+VjnyNBAh6z/xU8UP7
4QkjACpKC1ecSfLkmkX4AI1kgdqz1Ui7pkLQgjmNSIxQYBc29vlkqa0kCysaQqXnmphluMXrYTTP
4hyhYl+F3Q4rlHFd+di+0Fx8lUjSNnUdlxd8Po/FUYiOfv6bDD1xxcY9IWQN7YIGdQI/5o83lgCm
HNQ4UACDzECIoB5bjHUTjqsw70MKoNKwRGb16zyVsBtQhLGcBQ+JJaRu8zWX/37PwiSSDJKcc9C6
OWeCN5s8qNx+EQHgHb4/y/PvKycs82NOstTeOiiOovmcEf6ySidSgQ2zOpQOBwzjtQY1fSUKSPWj
hE5rKMrL5BLPuuH8Vet5bBu95r9hGdrRdPD3CShBRtRG8J1zgJ2c4oR8Chj4aLa9GWjx2Gz6+tgn
az48YuRY/D0XkG/cpfCbqD2mSYqYr1xTP7cLsSmm2tJh69s8U1U6PvY+GHjvb+9bbcchcLfmGDfL
RT8UMq/4hBSSBbEuZADX+jYQMEhVAGpiEio5Xu0ImwxziRzSlKFx3kIB0ZqnJPx/c/Jqh4zqa06v
zPIHzFyZRqSJa7QZ0AdtefGjxVRyvgFm14h5g62AQdLDnmrn91vGSOi1HeSTu5ylfCnKlim52our
RQptHXN02k76Uzk99I1BT1Wh/6CtMUd23gc/pF2cmtL18wVpOXQrYNShgGs9CmN03T+K5zMLuCvu
/s+BL7IU2W0c9GEi9AlgAf8DRkHI78atjmluZuivCiSOJo724DzgRbKztJrOoxat5/E9nHgGMr8/
0lmfmVfGMMJMmQKEV9RM7r3eXBSGDHO9xkhllRi64ZDL8EFQPM7UEZjLfonF0ani8RuFs00QQxYC
uMIg94YTtPUUQqEqZ2XDXxVQt2HsurqSJXwF2dat61o/hi5ZXdy8UsnX1yBR02jQCzzKa9WkAglt
ZAtY+CRCHFaTHFn4s9XbRxsWvrXGhRXL0LnmAY+1axQvT0X5F+2D3+6MdJXynW+hO99oxStOH6y/
8yUzpA7BVf4Hcj0FbXDVHK3wZsExfyjkLI95Cj/7v98RXhBG5h4rydqKVO1ms3n/Dp8mVthTVCPW
fv5KVEvD6XCzAl5uvULUrP9iz/ncXIx37vg/W749+i+mUvn2A8tMRdIBjASCLlnsdVsacLQBMKmT
+YomH7GAP/KcVBeSzpJdlMnNSfdgXfzEPiCoVOi6ADvRYzkN/mc6ZMh41NjK8NQWaoXoBq8YxKrM
/3kRQe4xD94VMWuJlZ4tJ7zfqodpln/JMgb0H+sMlmFfpKG0FWhbnTnQacLnwHr0iod2RJo2C9sk
m2Cp57DDncSU56XDbJVqO3yn8jA3+O3keQpdE8jWCEqaiPPyGcJStK6qw+OvmkLMKfsEz/dbmY7f
visqAgi9YIvdQqmI+8xYoymfYgl4IlR7ej9JzjyLeE9LbMzyjLFrnDHw7oafUYdhLIEG/AbIE0Ae
WtyFtEitz1mmbxOCM3ctvTxv5tnfyZIdMwhiy+Al9ySNzbDGLgqINDaX6lK2VPkEhhoQ0HtyAH7z
Zjh7bbFY4ujuMTK+bJcbXmxLUixLcCjlTSFi5kB5hROlghH2xL/peZwb1c5Sugo/cr90wisTjaWD
oMTYtXyAMN2tjPVn0cevsN0cl6SxiqHBDfdA9bv3Sr7rlsW43Flnum81c6en7EGNHhTQD4tJaq5e
XzPgGa8wkcEnxnb5NvlyKcpGjpYa8thMyh/rGqwJNFFwTT5oAmAc/4HAOjIMKDKFyjVbENKo8uYA
WuTe+D1dt4BzmLM+T3JUG7MDJ9z6kUb+/fgUSxUIuysEOVH0bAiBwmQT/uVLyRZyPKvp3q4Q9XX9
BsesnFIgoFp0Vb8voanlRUvhRgdQmEA5D9F7056tGeX0wX56e40eDTGEBCJQuaVKjjJ05X78QHPi
T9icEYTADjgTwzYDsh48+O2RCs2Corf75QMzIOzUr1DGSFnicy6g12qkioWw+7DGVYu6EJfrzLn1
x9nzrb8g9omF48Niui37x3HUTmICcdHMsqnIHBwpudHSTB+poBIULH49pxsxSxL5e8GB3DrlMe71
2g5gocvt/43hUEpXg2NaOZjmwI/HGM8c/3zMfeKhqk/JHzWdpricB+1MHvBVYwo9Ca+M0kjuXIGX
BTEn39Yj/aFzB/ybCROgcv4jpu7hgAxdRgIvykf7tA8kQlPCN1we5E7RU3DAhDdQKNdNTiiQE178
jsO5+Jebkggi98BGGwfTIvhi0lZCy5tqSx0C1RPIbH6DaN8Wl0tXuSJ/+jhsGXC3GpWdtKaf00VN
RGM8aQVW0R4hry8DZnSwFC+ivYHPx91S2xsl4ftOVIIi2R8wZlLvczEj9x8rvTQjPE3OR9IcGm4O
gENYvXY70lMaE45W58UvO7QUf71s3gp+iGdUq5KfxoyGPa0+B7GpSEW1H7BIoOVP/mT9F3cPDEdJ
Us9RCn/KkrpNoUAuL/LdPT4mZnPeU4k/1Ja9J0hiuSPEDBalU76nW1B7uLcn01o50hLzo2qdEVBM
oPIk3kAlpgZqfMwEezPc4M2Tn0FLADVIBn5lSGdlUHaWaL+HcPMJGRolPFVPp1Wt2VugCAl816Jd
klbssAvXulqyqtOAMhapH8JvU7v1LI1RwjFgKwDWLmP7NslodtkNtWMw3mXUdnT7o1XFcUb7jSyX
eSaUXr9342ZBlRmRUNmkYIYoq5V3aBRxxuT+eCdG6HxWPwsaSLJtFnq0wlAuXBjnhdcgu8mkU2QL
xNzRQTY9/Lop9SHZTP7ul4euLPw9pVKWNwBh2jlUepYy0R1sdv1K5ijQO6fGsbregYcGUFvxCllA
ehDDbexOcZVxZ+XvXRvKfdfQzUpqzbK0zMy6NUny4WJ8WshXJWtUxhbhlH0O8X2QFTVn8ceL2Dl0
sniSkEh02qSr3/+Npe29e3Oz1AJezU4uxnnwJJfWNANNVVED3tt48jXGBPQvi6NQSq8g9EYNJ/A3
cS32N1CgCvtQB9oMPbOmuaj7MyBsRyl6oy5WshQuzbWcmBdfawP9aWVqleLK7KNsMcfRu6FMcNA6
abS5ME44TgNGdmOFfPcvg98IB4Y/gUK6fWBVghoylInY1ybGE9uNJSMUhxF1Srrsizgz2PhaqKRO
sYT+HFI+qChu/p2gwcz2qnLxNSN/r4/0IWBZcnQiZvWGPTs9HOVMe/i1PwF5mKZEsIfWzM1Z86sR
NwLizLcHPzzTO9w4TX9D7NzT/2y7yHi5YUHxVOAiTgrfObwKQhfZbjppZJ9ePt42N9y2MRjSKP/R
yodr/0VjCJ4bfH+syWXIcFXpGWEna5BGNnnXunkx9b8qwDYaRxCokHApdv/7nseWjX1kPEyzaRfa
PuOTa3eVnT3vnsfivqzaIq2/Ovccwec9WXbMPDAtE0eVRc8aGbKKvryxaWr4XiPDVYerF4GBXFN2
X8IdyZuOU7CJXAjKEJXUgZQBqUaZBtlCkWcUocHT/yV2PNj4xjY86an59GPSzldbxm/DsqRKufBK
iLcBEk8hr8qBDg6CVEbwElXpXp/M48cg8oKgSdZShFJWFdvc4lEXcqhr+dLIwjeoCr/bTG7Qzmo7
d902RlY6k8oVpQvDTyvOYeyS9VLsFoUpHczMqgtiLtTmZU8qJb9uj4xfEmk5tayT0pjX5orZ2llU
oa4nlXwtW1PYbW6xEeAyEr63yVYtnbralCWnosCArS41n7cirFmcWacPsGqwPrvJayse+AqniByt
nrMyABaq8hQZQ39BC2vOrZQ3Ew6NLH6zQiMhUPShy3YfZKTJPOw4WRc0c+1tMhMtuJZ+yUSoIKug
9KxiLy66BlLysFzc/nWyE4zZ8+ERGI/Y5Bl0CHaVjZKw4l+jhhqJ+nq88Ie6FuRCczzWhKXf9L1k
ksQO5XKTHcfWKJ2CoNSP2+YX3hkv659pLLrAgwtrWnAD3UrrJy49pe7778W6ayIqK/UEdpWJNJYO
O7kIH/CpNysnhSQy/Kv5WlG75f3td2gQxExH0qCe+4+qeP8M5kE7uzrRLW4fOmTqaVfiZD5Yd8BO
stePYxZ0+u1IkQ0CnsVd3J3Uww0H0WRQt3yP1JrWlb9B5kEFqUXRLBSeMAVtjkfVf9Jojium2ysh
o/WN9HtqbQu6MvZ762DnLPcP1ZTZZW+Z4W//Ns236ptQduupCNbAxDQFSdFFfKNvi1QxpbYYnret
IThkGbrjCMq0rFB8NnPFg0UFPdVOynPn1SFotyYOW9523KoMCfEzNwuiOxCtN/cvToePT3SV+BNM
DPHvIKRuYgCwjluJhdXe6bC7UHB0QJktJtqGR7DiYQJ8jqeoXJXyWHbfejHpD2My5RVKzAmwM3Ju
8KUJmYFSjMxAALTZbRkU/Sqf82IP7ZkQAKbbiSYtS6WyhYC28AZhsGYsAO/6TROhungqEO+jnKqJ
jTSNABDUocoRbqe91JjaSVtJ/Z8JjTlxTjw1kvxPNNZtdlc9guW0uIE8OcB9r5QF7fgoX6md90/l
o5Mfm7MMofLZBNGaY/7oqX57+ZWLmc+YUMI2R5Q/cAWKqCShf6QIBsEhdLTy2Qz/PTso+JmnUFoI
z3ja0tlKxgJSc1dViSSZZHMrDnqAt+qUj/qGJUPiRcJGGacACuWW0UeAB5BQH003Yc5Y79WugCXY
iV779H5DcN0nGZb6fTtA70nv66VgDkiwjfSizr4+ogDQh+UFA1rQsMzF2Yo60m4RnSxhrUJ6YkQP
2h323eSJKjpjVhRIMTKLrIk4oaOOYPC4O42WRiOhq1CRqUXFRqOC1c72mQrJ5/0QaJTDQnNr7Zz/
LtITXe2gGjePTV1pr6MZVnguUmOsIK5sEL0Qr0sFEUxkLBPiXkLm7vHWoIM9BvyYBwBC46wkCGuQ
cVoHA90UV4lw2Qi7KU9aVtFQ1eCtbYQPkXNNMi2dypH3Fj62lC8YAmMyb7anwn4hhfIHU7gwkLec
0bl0inE6PBt1ZRvvyM8DVLrFYha9pSkMK7krwFLjwM6dsJ3Nc+ZmZD5qJbaqq6iAYx40jMW9NSkb
p7V+OKd4N1xSSIlntmjfJVD/J6Bjdsa7FRu70U/NEs5D3BGJs2rv62T5MwHG3WPva/mSUuk3cCZv
/odyjQjmqF/MbqTynmZXu3hy0IrJddYLCQnOutMA7b2M4bWKtMaYbr2cZedHcaR7WWbtwqktolkB
E+uF4nuFn6jMkbzluDx1l1O2HqLe3zxm0dUe7CbKxHlye+44BBkQbsf6aPJSOi+5PBeBxzUo43dv
lDwShcA0NXB0g9Xc98W8TYYesink/oeaxbm7ZTjz6Vi0SUaP5aFO8dtYpTg86zOg0MqIOBYEvClg
yIULXpo/8mL7tla3eiUFVNbhSBsT2W4kyiPtCHUgImhe4OGw+vAZVYPzPdU6WIeEhIl0DWXMEmpg
vQgFRDv84qDSCVfDGknXTOpxPB2VUt39GnxjsA2l1nsLIMTyqpDCjxoK/Z1DkTWKL3L47L23AUhM
h+sWTsP0fPcs0lZw2VZZObwWMSRCZK/XYUh7BR+8d10Tan4kHfKKKtrd3ch9FVRtjOC6CH/BKSd5
xLxAizHQDWMLwXmwhGIdftwKz1q3l19uF7aKck3FzupH5Vf1iZzMhhAa4tMpOD0HFtDmLBiEeJ9P
3pzp6PQiSrHTbt7GnVkSuMulL+j33DTG10Lkh7Kc8pW+I0/LHiIXasMEy4Esu+fAFmXmpil1TuOk
/a7sF8RxNRHzmQI+UnvMhMaa/xoRujEodjJ2LWMoBJSTlI15CHHmNNRJsaxwqiw2U0Ue/lTX/E2A
jQJj2RpVK/i+KlGy2C/en22qINFY9fDUKxbL6WHE7bc4vRFGorKN76qdqgWLgmtuSekBnxd17ExX
QyvbYeSC2aF810c6OMoOTrMykICuaUp+Uuh208Yh75p+E4rpzHZsPjaKN4fKbFNJT7vgPLFRfUeA
e48dcmzXtM99o7UJzDWo2ZxBb+ShdFl+DL+ZdEnBPkXBCW3zeU709jNV9Y2E0xHM1A08P/JWvvzJ
9avaIBwAaK2DsQPAuNPA0uMh6eonQ5svYs2Fs956Sltn0FI4ybJXLyS3U9qpudc8zj4te4DQTclo
nu9sbs5lb25JO62NE5Es4jy6Unyq3vT0sEL+adxQiwNaIresUA7na9jeNWhF8cPOVbUthY2uxO4+
Fq+/6+WUs3+BeKRTtpH/g7fG+pysNPSviDOD/R2YY0N5Y+B5LpW9MFMH4B5f9rX0VE4Eg1lNBgPG
XMPd5hLGhmav970ui3O+63bpw2xyDkrtCfigD8MeoPJN0JxxpEQ2iZP+nJ2YuXQWiK6EWmiMBvox
WGXf2n3FpcGxU7q/DQhOi+ca5YM0y88y8tLh51EDM2scDd0K8k+TcM9KiELMfo2dGNml/X0840UO
nAk3DQLgtZPEodwK9l7gnHZce3ybZHrcs5/1WjeSkruFI8uM2mj0Zn1nDv1zwfNcnDvwo56YOGgK
HkjkkO7/Xdm5Pnq272Lw2Q0JKjdt7ni1ajidKPLWhCCEf0bMmPSj9b1q3Qbe5/vTp2EZrVQaLhJe
ri7W9+5etddWoiiZJikrfp1Y39/hBY7irOPFRTEgxgLSsV1+UwOVWrhUFkd4fXm49twAEfxHTpQB
H1/fInPpIw1YXa8B1amZiRsi+GM1JwyYVRh7OIQsBj+Ib3ejTWfGhLRqw/frLq/y6IvhBAWgifaB
LBkPw6lcIoYdv7zhdFtRDnH7mMr0ILonbO75MdqIVC+FfrXzdFXNXLar5u967P2lFTNnRK3Ud5E4
8xkH9/5V78hjykj94k2yIOq0wWtGG0BNTd8Mw404F6Le31r2+N2QwP5HzaOonanTsw/EKF+acnSx
GcDCF6q/BNL0oLuNcAjNZ7P7VGKFs/j/RZ71ZhjeLUqdjzq60WpoiRWC2WhwQkNNfWvgH7OlpEiG
OZLKFA4rqrMNQ6XnH8167RYsCAkt7PZR7CcOEIMv4EHQ5GnssBGGc4aCepkfduqToV+eJxGlx/n0
dorI4K/+XJxqdDTnJDYxYtyCD0ezLZIWdPFJDNpwTRHw5kzwZTg4sbg6yAPRwgTjyYB3bTSXkr+O
qH3QFnEpDaCk8y9DaBRyrEdqdcCmn8edKwQNISan42XB3Q4KseM9XySRWJkQEO97APR+4vilz38O
zhwsRiUg8L8MWfSxxiihDLUX5qNo1wFMcht9AumrVNZHvFAEWhs+3OYxffPTqEEVIbYW+xRifqu3
0nM1cKwb3jy9GGyxBZ82QOgNEzxAe/YCZo5tr84i8eOQPDV7Iy5eOWqXq/Y63PLrTNhhe2hs2IqQ
UOan8mvJfz3LPvdWje9VGcu/fONQFjbu42uPphMbvbUnj4f9AkQpuFRi8qS0F7QozIjig8+xshCe
VLzTTCny9rurIMGc586BGwlIuco4lwvQV9jMMFKJmEiDb9syGVOw2b9rzA/sddDiMXi6RTVRLdkX
dtBUTo6EUlNX3TTwPsTfMXYROqkeEr66Cr7wDtDo7SzNTHcwWrSqIdEnZspmSjlc7We/p9YacPL3
z57609jTvtFQ56EV1mT9loaCcUAi4qqMwB9RbV99IL+iMV75fQ6lQod+SaVqUp29zkV7yLrQUhxB
wxb8jixP2pVt6QNJnbUhsB2SQtWA5QUpDsvLJv8e8vc7WniCG9lOOua+YlOXuP/Wvj3n7L3FywgG
v5ZpmZQlHtibKw2UHOunOoggPUmTWVD1OnUxQoStOdQbrTw2yTBecQdVxro0vECsMxJPG9lGqJ9n
xZRqYSR56rQ6+xRUTj7fVUsPMI7u5KowGh2il7uwJdHyyLNMkdBG9OFfevtW6XuOFc17NpBCO7Oz
0a5gmrvOqz0R9gItihZPgySA0SYbsObJnasRFCIw6ZoTyJtdAzxlZIqsy+BvWaLRBWE3HBhCLrwO
4qwnSBB2ly478r6oIdrlQutdf/ZfBWFGepOx9EW61Lm02oOCaaB9xkj+mWvIdgAwpM4zhm5RfnoB
uIrdWP9eISFYOgGI3tFcGq4BuD8w3AOod/2xOE6zOgndqR0BrFv/SIV8+JQEX9Hq0VP3/qOJ/4pa
VHGbFqsER6ackC0789UDOFdxyHhku4XwTolBlWTdm6ttLTwjH4Of03GatH9ehsa9NAx2pweD/Hhi
pWR7NDr1Jc+ncXFG24Klme6GDu6MNDjj3gr7O183FogZv2aSLfbyH61a9dAI5gmRUPkCcGgqesmR
n5QZBWVV0s8obiQAsmu89M1iC1JZoNskByFkFpND9BVa7mUCQw6o7smGOnF2r0Ezvpv14XQzp4Op
TMKmDdnEXFwnhLZxYjS9RwPjMt7r5qRCpqZkNx7v8I1kba4lYjD0chjXOAPSWVlywScSLBqIIy1q
UzCjoWBzPyjVUWxILTkeCKOiBjgX8f6HFsHAP3tDB2msWtls9X127H8WSjh4kvvIMRufMJL3zvqN
TlDy/jNk4XLlA0X065hORKjBsy/gJCHlJY5MYefP0gktqCMm425atECtAEm4KVM7/o9kxCtdw1N5
ea43Mb4guLK8/ZDc8O/d5OFGxzS7hTiOeI3HjpDTzpt/MnV1R4g8mdWqjwtH1b5e4tnAbloZsBR7
Obzkm2EoVdIVoTdacCdd0BXLmf0FsAHOJ6ZahChcG8EXrZYw51YP6zk1GpeqN9KCBAokHjWca9M6
vDVvknFbjWVfSDDvyfrTQSIuaSrfVJPIhOxaQITwI64/Aej4K+oYwCN1hwXQsBvDfk8gO+ShSSe0
+bVIdbTS1AOjSh1SE04mUB2X90e1Uei6a6ijzWA6WoOCAduIM5mXNuv0pBYmDMjgGo032mlJzShZ
b66F+BrBUw/cn4SpFgb1A7GFcsSe1qe3wzwql5x2BjJothP/woO2ICbr7oStgYazk5URadivPCEF
om4I18Mi78wQijGBa1JGsHudImd5XPHTv90zbdIJbTnaagyLUDvLFFwinMEU98Smmp1u91F13ZYx
zTrVwbS9SeY3ITMN8eUM736eiuBua+Q+RPLULStVgwe7GJONYsZQI0RbBFJMU+UtKW/X9v3ly4Eu
8m3ufs1plA5U938Iu5/QRBrLyHnESB16+luDUYa2MYYp5sOSd8DLIXoEpRwKyO+pcmpJsOejaorh
42gJpsovMFoJ7ZnjjfpBKST6CsmS+Rv+ttJcLN9ErcVWmvd326vMlj97ipWaoLTfHZkUBWEcFiNI
4DUFnd1j+Xnth1yCRQaLc558qmyB/J9dDZ0mDtVt9OiT2sD8s1CSoLSmrNS9grL1I3KKvWV5yTM7
w4pAXkylCqXdy+17M4nUaXjhOMx4eZtiWXuAb2Cv++7jTnu3CK0ZPTA4Phhzhqx0w/SG5ptwBxAm
TeAQ8XSfIic0kPH/30y7ZR9HZMckYOElpUDHi9/oI1NFemmSV8O3s961sHZftV4dQiNjL/Y1RYKX
bXvOoUOm3FTZudDVuTQm6xo2Sf+6T6bJ4j0uAfJ4M60YwDIf5DLaAdEV/YC9Y6nRzLpI1k6xx/Hz
51u4CqoZB8DFyn53mmYiXFoxj36/bZbJ24FWHVBhwqBHC8F57803+qnV67vWoZx4DsQShb8/iDi4
QLJZtBSeobnPXMoWTRXeSqhFCRnB5IW0Tzn7+aVmhjTV14TznZ/yEFS+ODmjdNKpEPUXU1SQKHDY
/0gMs9H4jZeSGfvLFC5o5a0fHz1lDNm9ynZE+ZCShn82oN2bhZPjqIhOQC3G27vZIzIXo3HFw64c
rlSAiQ2DWox+OzrYSCuvXPyrpSK7rUeWyIj+OiX9w/IT4f16MUB9YVhrZLC7wTkkKJmyBLeJ+apH
q+B/tH2jfw+shtJd4q15JrtWE4GOT+c8oZXxxKgHqwmvY2QkXnhHbt3Rn0EN3I+PtiZU7A70yxDY
GlbYZG/NPCEzGDub/OR9Lf30c7obzT9iynF3wDMaA0ZXiRrnEgUfNsEOkGRN07Paj17NLfZ0mNxQ
h9T8s2H7n3kWhiFS8YN/IeSMFmFOg3BVhawMRf7o4qImmzJivq4lJHhqkrFhhvc//FOWk6m/TjTu
wPcXcWblwXiigPn56DhN6DIa/Ry1uOpcqoSOhg/TNodP9XSSk9c4jTssxTPK7G3qRlxNpmBIMbck
SMfoLj+peMAc+fbp+3r297l9ej3PV8bOKC9/LQm2yJOGWsYaMw09wbuCcMvLsbHbv33+76RSiJmD
c4HO5R7AHjEpj36z+NyDzJPDS78VjRVb5lxoBep0uwJJggb30iAdb8arhpY1m6zFdKQU6nRLHo+T
nKitg3Wq64uisVtNGKF8v0KuiI6z8o9nBcSc0FHvZ9ZaND95VIULYIywxBgrwUDD2ithWlOisB4Y
mH3u2gmp7ZJWRgkGcX1X1uNRVD6FKKKYSB3VgZwu5mreMoaulgYCvm5T2lkqPDjd5yU4qdI2Pm9O
o6lro5WQ48QoJOLUBVE8W+YBdBHxtEQ11zqF/29B158YgurhMf47m1XgyuCAWpdcFeIV2q9cLaEC
87IBYGpn7LF9EzugiT1wsXcFGgTWq/utlPIkYfCb5ZGKOb6EAi5Y4Lxi+VX5kIzixNL8DlcSRzsn
FjqkvJGSL2tcYT9P7CDdJfWcGZlZRl08vQ8N7VgvQKRsnznbAUsr70Fa57dqU5dE9GvdzIO7Lpjs
pcTbzc/8wvLbzHuvLVFrfol1bMg+vdLA1OmqE8O0G9fOxQVh99s/6AtxtSwzm6pnwWBS8Iad+I9s
MC4qFiDtRAd6tXPV0ZeG4QtTx9DxjSB9V75RhwmGfDScvLXsnz/EuJryKupYWr6TLhsnDmdoUduh
+VCPCei64DLvQ+EZ5z9qGk/hRG0vZPUW/03LigqxJp+A87gZQt8dwDZazVfhmqiI79YICdTFqCib
8hzGb8GX3jA1u/1wq0r//0YEoNrcHQkeEiVeIYq/WLoNrSn3AYDHvsTxagrjMVUpU6TlD4+kfDpx
I4jktz25k2vgcPa0TVetAXSIjmbl7tMjoRldo1zgpjvsIJY8VcVOIkzO/LoA4H0p4De8Jw6MTmzk
nBA42GUYLi+t3xxKrIfBD6WpK+mQ4nChtBMPjHQsHpfYeEBnJ2HY0eUsrDp1Pbn3nA471Z7lCWRG
2kyAfJswus1q1O6xgZXo2cd7zybGbDW38DbWgBPA3v8D40bgZ3B1hl+nnigwM1WYYuDoMK23rwOb
1TePyfVu4ve401ASSZjnRZfmnsuMABWEyrmd7Wzzkt0ltOE3tucAugBKhWdOrvPPQi1AtsuzT9zy
zPD4wob5A5L6mo9pQVQ7hyObrh7cS2XkFSFvs6QVSKjn1a+LaF6LJrCtTqruyTDps8zF6hUyR/DB
ORFiIUFQLbhQMUm/0NbgYkaljzFnbJ+VSbTTeduS3x1Fn4b+1iFnEdii/OKepSSfKixrK5LYv21R
IHIwUkJDmAnNCH8+swjaVzgWwxoTEy4gjqFQpQ7IoR1UbuL5hv2Zp5A3DWQyZTcxcyUZmDRmW6Kz
Dj4l1GOMQrAzZHKGYfv5RwPXFjHTJLlUSrvwrSoRHC5PdNO7r4a9mtM6MqIxMCLVHf1Hwai6OaY0
jooKoBmiR2vzTT2cIO+hNLXI/KtFvlc9CZ1CfkfvabTgXmXxQhEgYshJ3CZp1fbG448C85Mr1xQs
UR+nbNH5qMM8b403JCO40Vq4Q/gRNO6HIvPnUGQW8jRaYApK8IW3Ff3i9Y20SNFwGDK+BqiTdpS4
pxosGXk+ZrzxLf7AS+mQQu1WUG0PIWQy5lfsQhZOmQCUS5yQH8hafl17fQ4RWkHVtyRnXptU8oZf
fyhTzbNVbu33Wx7NcOoE8Y7kaMTu9GCS0a0JgdlHq9LNJrfqphmFLvMcVnUJZ3pYoYtLxrB/rat+
Hk+H0NuYQ92Mem4GWgx2IyUs1/Q6KakwQ0ZQpENhFHvDHEC5bebVfn+s/AeeCKTTJiOWRdvcwTLy
BwAwqj19XY7zT+9GjAMX3vshQD45J9Dd17e9n6BGKE/xOPMZ0haoZ6j3filPDHECI9RvPS42f634
gBQXdvUdz15KaQV0J/X/OwvOCg2kPEWmFf1UywTLvDcKfsQdyNAAbl+D83o0nChhkaKlaNX7aD+P
zuGw5dqKQCiqFBN8TbQWlfEbm0qt0i2Pu0VFoS1Oj7joKgjkVhcxYxpO1ii4siRgfTNriFUnFVaw
qXSTzs0Ox969ATtncNZ+aD3dWTbxkBr+WfwS/SjzHqoLh41kOgTmGXkwpO0TouEOH4sX/5hPULTI
tJVXAfrShvFUOiFq3wJAg3lbqEumdJfFbyoN0AD9J5yzUmq8aEjBRJJqtx4tXNkOZBc3aBcJWs+N
mU1PIjyD0Tt1WgBGwvAAicTvJWae+LQ8ObPxMeoLCk/Xtl7IOwwEi3cktXpjX+JdFoTHQ3GaA74K
V2ukDrmUWMIDeR+O/DLeNF7POnZPu6XfpWsHcH7rdQUuOtwfIBrSBlzcj/dvrPucQoG3vgfnYiRQ
Mh0qhLQayEiQmGP+eXkpVlE1QgNX55RYMZl7EuY97BQIsN13lel2F78cQ3DkvLxaD0OUq+nuPk1Y
0+yyCg8wKyGJYE7bwBXVoYh6rQ8OYGgAHWtLO4GcTt/yVwrYaHO6JUDDBrB3y+rosXskOn0nGDnK
zESU0eqWxSP5Z//t5gU7wA0Rqcbv+Jnq5oF1zvsXQhCnCGo+vVv808iSN4dTe/AHOXb4Yejsclks
pwUxXbKVPHBkUvT3XBRhOxxSt+xPgOYrXoqwVmiGvYLY6Us26Q+n/bno5PsnPv+k3qVn4JmJQFO8
43T8KTC67b3XA7Z+58wFN5kRHzT72qJJ/4FH0ZXhfmy55hwAh3Ktdbz0L9TkFIQco1XImWzAsnhL
ABFKbK3gKmBOxN7Gg0xMqUzqLQ8+MdJu3MUSZv5Knl4fGmEn+V0DXR1qx+zpVxv1h0SAIl9oSIRQ
dFoPRiDpYA6MvvR1xVYGnRol0IhXe/asY+VyJ7s0icojIOLxi85mRlTsJjDb8iER93G1N2O2N9Vr
9nxBn4TuPjEdiUaGBWzwb6Rj/0ZbACp40w3AFglMnce4I8ndXaFBMS5oCXht2A80JQTEtVql+lqv
5yKZzKKA5s+aiQDc20M21dTGUKlo9kt7JMG4glps4DHnbspTmnCYDQyT4RspiVJtlFUigS3HMdDD
nRv6jYLJciVL9SNsHVpHpAiLXUmMpnDGqOi4xLaNVCmEcsKd6HZ4l3KirxMH6xtRTp7biIi9UNHh
Rez030nb5ti7gb49Gfq8my6p1X48b0AW5bOJ+RjtIaI7dkzFgCX07vGh3ow+7UxbAgib+smCH0ZO
/nR6p2nM5kDeTqHlKXm0fGhDVWpbYmM0oPoSpxz3lsxXUj/45oPNyFQ7IpoAqg10ZEf6zgBTA8hT
Z6svqn6XWdAnP+UpXf5Z0P1IvvCGQeAvcmpwwnyhGFpmiAZLJC0xSlU8T1jrfJGagsQ+7KmSb+GM
qj+VUMghIYBxjaBaw08+FKc4wC5Iq24ANJ7BJr640sLdSDy61VEWpwKlwKkFEo1ycnLTmeD4LbwF
GQwZk6uIEuUg5c6fPrMpcssjROQF4lhxi0ay6qlrYGdgyPFITJhnzUVl7lmxxhon0ZqqrJCTsHVG
vfd6xGo0LNiuCGXOoH6fU/flx5sNvq6ME6guASEfS4bvQS/9J+GiVzJAbZZ4sDnXrC1gXhiFwFFz
Um7NJXDX2SQJcj5ik6YuEmZL/nljiqDhKEojB4wYa0R5hay5+93q3UvJOjaOILWOC+LUhOJmcOvH
Wqrt8Ct2z0GkSIDy7PIwehj3QAFMKaYxOHIsD9f2SbcQLbI/X8e20txoXZNXfnttePdN67rb5h6q
6yhQXtXYqHJ5MfGIHFG+B0P7t80FeJZHKEdHRgoqfpqoV7h5QFXAeu4L59sEgoKDK/osTzYWMwRg
jhldUTfETGnooK6RmIju+ZMUO9UivrqIu0MagcMplIjhjRhpUAig2HR43h4UUDHmvFFpwZAd1uEj
7i2OK1a7QekQYygjAUDMn2QdbI4xMaj2K21CpvUn8JCzTVdAGyxqCDweU6z+cn8hP8ZiRBp1Xhyd
Td1NKGa/q3/n1GKQdHNkQoUqHnPE3Vck/bO2KrNE/UgFSgd1Ba/ltisUJUF1AxsbI8QhR5L/dAOb
LqdWzAwT7GODbxaF/ooiLMweT83d7cJGnJQFUMOpbj1rVTwxAMKAEL9cZS5/5va/EutXoV/cRu0e
kqLNisv6MSNPL/N4Q/q+40dKYY5TLCV6ZvS4nrcGZUCC04hI0v8YUeQtgrq6BFdS+ow+oCxBeujL
KoEc9xv/EO3I+jy/z48q+dmFPejigB5j+2VzYywJDUiwumRFLZIULK4o/ydiNtc4HmM549aU8993
RlAKwD6iN4096obY6SzC6XhU0GtDDq7oY0w1EgrIjl+Jf9nIr6QQMxUWw1THx2TSGBcXxbqKG/6I
HkWQ2ZeYlWDQ3tgdY/S2E/CKo+RCG+tm5vJFecHHpkccrRHnrLyRRGUic+yQu6rgKgxeZBGXuc0Q
p90kCjwPN0cvQNCw2nKuoXO0ONy7gBYzsNniAUjPWElS5wdk+Ko7EbKP2+U5h1y33TEQtKj11qZk
eTFMfFgOLWNdoEEIvnu5pZK0EBf+p9Xsx4fU4Pb5c59ZbUWUxgn1Zt2QR4DtaexSrNApc6A7tkW6
h3XikwCaW5BMx4zAOhKes7zff0zCc4AG//N//o+tH9t50CYO+l1CqsZpwpST4V6LVvYTUiB+T79C
jWMYFZ6iD/rTsVgEast33Bm72kc7uofyePncEDmI7Jde5YU2i4rXh5Mh2Eg1tKrK9uuoHIXYKEZi
PGHFHM7d+Xoo95U3XuSbulu+k7iKh40N8ofs1/9JkQFerqIBYiwE4DGaYXKrpsbrIWlpkwOeFOtP
ZnwjYEPeG//PhV/C9MZ2wC5I+0bbzPDwFOfb/oGR/NdxCOxYBtOaERZKrzXWeB11pr6mOW+A/5ZU
KkETqeZp1rVWaTowng0ORX7qspl40jFDCklfuGZTLFqlt0yZa/0faZGGzsiiNfHeiKvDb4MXGhug
fYgWSvc2YdsoEulIgiEf4R1tpeXjsid43F+9nbwFNl6/iploorC8ljqY6RV5NJaSmLjXduWT1LZx
d/4JrLjSTMctAosduZiv+KKlUawfFEwUYmw0uqO8EFM9e6e56dFhEpngX07YVji/xcVQCbKI2Vy0
37RbW3Qsg+WysKaNNLNfpInTknFFVt+WtDTVS1xqkzc4MI0DVEqC/MUHx+cYQlnyF04fd/xyyxQY
TP+yySf+tzxs7eBXYgp9GRuk/GLzu0IvOWyODuuk5XuQRwQGI3oJ1fFdCTGhiLQaX4lmPc4LQrAE
91sJUJavrEUh4OjHKS0tkV4z+hRO+OT4m7VjQVTNgaKHuYvrgm9MXDbjJaXWL/iEdhKCKAReNnnb
SIMA4vMKzuT25sw+5g7RtT2WJpwSg/h+abmCkpRlPvbTMIWey/Iw3Mg8AFODDX87wk12PaDg1guJ
CkH7yDhCAf8RrpndBARlcyi1MHqHA/ESC46zmUzPvATNH73ZMUZHxKtS1JLdnsjKFi1plXa4Afj/
dFVV7lZVxp+6kqx8YTbhh99xzs8Ixpo7OexUmOjvEfqCkjip5L4dE0W8lZ6XoP4GyUYKWYoBWMOj
+T93aR5gOZKFoN5XqRrdUBxGOdk5BEYJ9iM96IImwBeRAT86Af4CsBq9Y/XZc/g1UfV/6LJHwaff
1CJ9Kcl/fFiHNZbF8x+qMo59EUTGUvtlBGO8vuPz84Nsz4KgtnI3rMfbvBHNgBadpgttIfLxAmkW
ISWOh3WLMzrt7lafQPYRfwQMACKW8GpnWcsEM0CvwkXHcqn9Nqa5jNxP7dO9UYjvKZQedBq20/BS
BwRUs5sH40/orjr8Svt8ADx7e0ckd8sUKZxPymiHR2pSwOu/81F47VltB8jadXkRa8ZhU3V4DOWc
IzOHlesMpHgpuy4FG+eaU70SAFK7ilbqjPMDW/TWngz+0FEnlBXNI4KDNNMF9ZdHn7eyEpMMowLi
btoAPU0uLQC0gwFuGP/aS2hM9yZjOFRlBZGThY/VNKDlmS8Ze1gRP7TEIrG1y2bJdT/934rWnQlV
y0ivOMat5D4cM9oa5Ug0TmpwAASzZ/UIC+GaKlOUqB0OrQyoaysgdGvj33YZ8/ynnn8lYUm7Np+z
HhoE+lCOBo+Z8+cUdaL2uA5YHpzLklBTfW3ijCyvN4c67fPFmd2qb+mR+vtVIIQ5XwnPkDqt7TOV
2nh+iS97sZQ4q+Ni7hAiMrcv3Z8SE5z8uSV+7xSKD08OJf8zfuci/gRIxYGsxMCYB3rQP6Zv6Fn7
kRiCkNSGSiytsI+k+jwMWCgR/RvzRjvmr7IkDIWGYSFr5wvoLVvwwO/XHgpN12Y8UvGphV8FWLlS
rUE3ILbc6VNEYct5ZekGWwcDfO2OSda/JbcFScYAPdCcoO2lH1TDyjrwhN31tiaMsyUylFy/0mpZ
Htj3KPb9IfAd+bYNU9DzRyqHzV8UE64KekR9RDOTrj8pi2iEdxDQe7SswxsVfMje/n5+CYGjQzUY
9/lC9oRl+jw24Dn6HjQ3V/BaIxbKaMEm74JIezpIq/btYWARsr5kFuClR2he+GAZkt5qOW64Jiks
HdW+d/4/w8jmPv2HMCtebX7DC0pUr5vCxFaxmirZAmtOwb3fp6m6uAaL7pCRfkP2HW4BFrF2skdA
SncS3rDMRzK/IZYmyH0cs4tF7I/4HJSkdWEDt9JNuazCEmI5Bxr6eZrUJRjoaaPp/j59boVDbtZB
0K0/zTtA9MAuRhcQk3URCCtKDuHMZ8X2j5MkNJNdPp5+R/HjWCu6WnYjpU2fADnBhPQ+xc4WwtLe
7CC7OMHxYEhEC9V6eNvVgJ9HVIP6fmHnVDNSz15FCAAdXrRmx4u2a1UWblVte/OlOi40M40azB5P
Qz4AoZlHpRjMTS72yWj9fwnB7YUafH+89s8jm8eGJO3/3f2dlw0YDZjve9l2Q4W4HRI0Fh8HaWoG
KwL6yKlTXJcF+eesXHZfWb5SYrvTJaQnAfco8gu93piIDsrVYXaE0+jnqmOF0Eh1NHTjMQ0jtCzc
+NO2IVb2JYVYUI6iCpZ9MIL3xm0HlSHGJ3epJvclvliqc+vyd2Ylz3RTHFZkCrCFksC+Ffmwwm9X
hJE3DQgKNLwuozNfGN33HPbWMkzbOE7UKMoLDUUi8gpdIYHr6CTVENSSDy/TOw1wxMW1NBbmc5rm
NpWa52ciSi8P4zQfSgIT0IB1HvhHe7WGNILu+PpaciD/oK+46HbCQEbAn5/VyApNpNWM3VZFZVma
l2NMH86kZBqBP2Rj3/7W+HxSU28I1jkbt9mCWzxU8UL74LqvyPTpo3HX1Vg3J7nxM1vAZ+kRkJ9e
7mNzO43k3FztBg57HmnDK5ghbLaHTfMVo3FSc7t4BkyrXafL2X63QyQUZpQj1EyXC0f52hqiWtFY
8gvp/loO/StU8+QX4UwnFAtfwIC5qIoCJqnKk3Dwam5tLHrsJW7gZOCLsw7lWBA1lPcHG2pfqlpk
WB/uEMcLzU3bdwbktoMUpG+/bfFi0gdSl2QbmOH52W/IkBiapFUwm40UrYi7BkVchJxmMJRemOHs
6S8Sup/dkvgnq+MQJIXY1XX+U/ULlPkNxlw/SJRk7vBIjgb+4H1xHRd4Zx9Mrl/89pOlP18Z/zB2
bccPO0jwRTeHZKJA/IEXb8vWK7BOkUvY66LPjjnAQtqGdtHDN5G4ai8eHsGPyZPCbiwX2MMHCgQi
JqmkYcmaPRuPnIiARqDSrrOnwmdo9UtlkPnoz4WlgUJKY8uGRNEiUZatGQd+mv+AUt1htO9gRuIZ
N5me6VR2jaUaT/Q1lucUzwRCE/+9q2y5frmt0STmSHvB8Dv6XO/ZpUr8BCGLvIUs8aeCQbUghqbP
IVVw1cukaaYfOzblA8f7p59rVemwp1c8g2SPQO/xu9TQjhYD55PW1Z/1Odlj/Aa8hJHBhf3LBGU3
NRfwDZxcdHpp3dl5Lp8zSte8eeZUVuWe/ouc/wDNKpIlQIDN4ok3oY3rUAoTeW0Cn9/USEkW+MEv
UL90znZY/4OIxswvLnCR5ERXLt+NFsOuZQTM8cT3ncWRRrKwqLOhepJgIicoZojOBhadFCDkQVim
RMpvGnqVByH/ar/qSzDoNAKajW4yHJSo2Epz6SQgEdSO2MQ7JeNhlyX9q7wgdtntRhCoX9SuV16p
ZUcd+Q47wAxRooQltfr5hNTVg2CvnbHbooO8+z2ogTVL71kBQ8HhbTMYWvlTOWif05jgT9FAxXqu
TC/Oo3f0dR8JhMjuwLiMMjGLdGQKLGI+7/i8O3exubbKCo+FzoFIk66ZmZ40Mza3aiaw1bdlfCRX
n+5MTkmzClrII494u3I8aLLoa+1hbt1lkUeh6fKmducckBtwsZYVo/mstZOzILbvTAbWFVK0FJwa
O//+RjAvsLSZ13A9tQUGpifb3gs8ywO1qondYn9iaXc/yxunbjn+TZXqogW96x99SDn4/mMBKBPz
WdU9XFabPchGZzk12CtcypJPu5fNVCR4XaTp6ELOBlnEfl5JVlwsoQ15Ri+Zll6NTS+kzDJUMaph
VFJVwZHDZ9M41WEWo8ZyhQl+F3sbmxEo7+kISGfsYeK7lQ4yfmboSUD33LBGLS92UX9gUoi3VOFh
HLozEKTfSGy+rQfUHgAbAV7mPFeBlVe3MDXD/+3y0l0J8z3pIqB4HDJ4zgdTRYfAQIATOt+rk/Fz
QEUUGMYsrBKQczYy9pSafoCCUu1NL0nOWGelvyQwG64TLB61OpTWVKkhKirvCXbHHJBpFKxlNk7u
/5Xy9j781aHost7bkZj7SPRAL+aukNs8n5lYl0RrDvyp5wMQg8YJ1yaClHKuYVE/3vZkbxNWUGKh
/FD/4NNg9Jv+WCTjMgPVGl/6uLZncoeyJ6CV1ISPcqmDNFHUcf8V1FpyyjEDzEHOVk55h8qyltzi
V3qmCFItA5L/7fMxqWBB5c0ZG9s03Z322FyUilGErXH7l27qGNz/mg0mlk7lOZ4822k7GFxG5gXg
NfyOIBxJOf+VLl7/i9VPkyYTbsOSFtnrwyxj6/588urqi01j1sF0cxSPFiwVnmT1zoK/DFGg14I7
RICBdlHYRC+6r0WnTXvbpb2dALjSgFR2HxIkR1Z2UqkIkzP2m5h7c6RELYVK6womRNe9pzAjqN98
5NubxYO6D/0Ie3ZywUnOTzGiM7TBr5u+ZqpPB0R4VWDo37AH11OGPC+O/HlqSbzIW4apdLzKApO5
V1tPxPhDKhEDZPWVsuoZ+SI7aEiWvwBksnRUXbmWBm8iXfjyRUdumQyqYuaWxVK3cLpmhi6fN3qM
e1miyMTEuu9LN35dPY4lvejFGY5taRS6HkYFyksfY2MkCo+A4lD/HNnWiGy6kkuvgJqD6BSgGoBI
EF2QOf3xQ0qhPj4f5kkqwjtu5nHmS+h26FcQ/roQf7Yz4AwAlTVAuS8v0cI8LfzfYk2pzzJexyyP
UpKYm2HeyoO7dJy7CavJw7Il691gnO8eiZgqDk7umy2s33u72YJq8Bk+kJHeF85Aq4cPgVCE9zDR
b7MejQmGxrUFWUhPsJNLuFsP587+LJTgyVhjTz1AGNYdmWB2Q7kxSzUpGsLesZsqgWeW4OTOalZ8
rttVA4MKULnDkCFWXzTbRYxra4YXv4Iit12aW0zzL8gKjYyb60eJXjOCejCoXUGbRt1khZBhVwE7
8Io6CQoyTbhfXR+SAasNTrEG5VtBESq0EZup7DZuhXvoKoPwQAFbsOwUe96wYG2tOPdjrYmMeftA
CVYSso1WMPOAn8S6yKh0TP5LAQ3SJoT57um1eSnSf/6FSsgIZYWQ+LFg9Aka36xyR3KtTb8SkWPd
yc+I2Yzv4z+qOzCtKxDvktvmFy1NNNjXAPPOp0ElsB14ljEO4yy+Xct2t/61AZHED1UGYRTexwt6
IWgKfjnnB1y5sTgPzG7hfLAevyDB+//GqON/hVxgXbbBh3/Jz+bQkS5GFfIX3rDcbJ388JAxiUmG
kLO/u6VOn0lxn7okPBGgmIQ0l3TApOI3WLC2iJEJXkUigYFg1gEkvjMdebOwdIDd2Dn5U1IwP7j2
s6d/4UXe5vG9a4mdG61Dlwmdrz+HOvi5Kh+7Hyc0ZpqrcET6Is6O4WGQxmJdAU4nVH4NFvy3mXMR
ff0qbt/L24G9INEBPn80FIsePhfMwdmJQNpmaxGWa7Y/OvNoL3BbbNd4/UaauxYssjopNKI/7aER
7oxHYTLnd2DJaUZv3kbF3sanamYaFq3E66GsHDrTUolfg3C5h86TSzRGBAibUWVgacmRGgmukHPy
rlB//XFdjyEFYCwdHXpY03lLbR6APKfXaddBjs7rT6Gx9JwLH9In+wi4GJQ8ktjjDEbqRtX9Wh01
kd1C6I2zqKi5G0q5eIIkmiqkejMmFYoSAISY1H+QKEOJgxQTm4Mi4mcZopDw7E2QCmVeJ2iUcGVS
bMsEVLAU1MAFPbCUzZBbOV3rOKhM06rrYvl/8POKkCutH0Wx2agClfwxjsXQmxx67QguHsfpM1zg
bW+6+e8Khfjx4FDI5cFi2VgLxxX8KIVSoFpZSOra0V46f3p5DM4L+eU2z0QDy6zGnt5XmopJNfvY
jXrtSzD/N63kuBDg+lldGsh8x2tfyt7CfSygch3m8reJ9ssmeOC+cpYtLb9MYYGOpqSYKvasaWq+
S4NXoUg6ac4EsGCOIzt0pZc+flSDIM2e/DnEo6bjOZih/l646+5f07iLAQU/GGemhQ557uRfd7No
+AHrMoAj3XveQkX8afryWLeyJ4zZsJQVjU+TMGhpfikVoBhQaT7ea4KpfOjWI1/edsSH8XyUZXfh
fmm8c0+LcNrTvMGzKJDA8j02vATItjrrE+DEC4ZRe/dWgUhF0EDMSSUSDG7JIH2xbfDzidh4mAm4
PdgWOfNkSgO2Msw1VnGaIBgVpGrx3HMAggyLVcWO/mvgxRv9E8GbYbeTIAhgz01lwxCRl5Jj9pcx
axXoRh0xsZggw+2pDQEjas7p12GNXC9BKSSy2lE3h/m/dT5q3lrA7k0Uzp7avlcuov2xtyenPd0z
UVsAVrbE8hT150Z1T1qhzCqUxbaP8P/P2jADKJQkVo1HfktYj7tw1m49idahlxlWx+26h0q3iy0P
5XTooOUsHBoe+lFqtRkhdpjTnKV6y89iMmraBhqy7ZoUrTPyWpCzEi2X7009nRcnXlozzPCZFlht
Z3E7zPinU3DA8C+VUhigkr4d9FCNZVHY8rg/3z+4ijzXjVo+20UfzJOVuFmM/4B/cS3LI30yCQCP
hb3qU9HuDD4e9tA5zqKDDBTgep65LDs7n0KKCEZ5F5v5TX9xWTBty2V+WjubbkoCLI/JBbL0z+fv
gzSpLCAcm4UYoE9YNHJTQHVXeGSBWYxbTJDiL9g6F4r6+RcvX31aH0n5h0odLh+79JtmDhUwrhpY
tEGMHU665gO5ek0Mk1OyV5+foxSSxpVaz1PUhqwn+JGRCAxJfrzRimLrVCdlqI3GkX05okZ8/xcS
PjA8NfjNEG9DUjyqr/A8SvvBp+7EL2N2sNERFFwAidJeHBQLB5ii8ytLSSgyZD4b1xo8v7Bt7NXN
iNz8Ap+PEQ8t/FQEq8ytMzpu+RVdIUmCBq1AY+RxLqX8XF9QouJZR5DWGWS1DM0lHTCZls6F6gh3
SqtahZUSYhn0p1Y+5c9BrOCV5w1hKIxoRLs7MOMkVcme+PXkadG5OKYClFUExmh8Low80cr+LEHb
LwF60nN1xTekq/h0XZd/2tkyohiTAkWvdIwoAHBVd6CeR9aHNDOnJfO5eGop/ji3NDXUKs9NUOop
cNQQLdzhCO8F+1eiBob7UPD7/9eVFVEYzmAu/oM5Ck2xP7s2q26FDI438Yqi5wqzZKGxhb/d05jL
y4Fuo5WtKHon7BU02Js+COd76HWwlJwvGt37FJaS40sOc2TEtbBy5/6Zhq6TduaAzRDEqKwo9eC0
+H1DtDPyZ20wn2eFzL3l0MrkB+XOoMrsrongwPH3W/CVTCk5pE2gu6jTg9c+Anm96v0ovjJ9nv0m
a0kidUUry4UKMsYJkNGVNvZVtIb+seDgTsk3/8CgDtn5IqTan//moMuRSCH/ZnjW1a2pIn+s6Uvb
Uy3MtZ+OA1fN56w4SzkP5OXXPUBOwNiGzKCH6Hwz8Zr2dKLxkRV1mK5vjSgeLoApDTHyIgvgp2sD
iXmVA9ji099PLXkWCkseRty2rhnrJyrFwYhY3KPrioBmgGD41unWOezDln9tC9kA0qt8sW5pWEtM
4RZwwfDvcVjGrtvezOZBqZFQBLDwpvnfN8FYt25C6H00mBnpQbQo2oXXCQHCzZLc/JPF0eEeDU6R
VQJETchorpHqMhhCu+EkB6dMdpzIjZ+KvXElQE+WS1MuYM6+4T+9fuwJvXF9zADuZjQniGA/O+Yo
gmVnBuJ3VSLzmGNd9K+HHsNZ9q9f/UqkoogZzefyy5TpmJn1GbFsVLC2Bq/jUUQjx5B0ULPSLX6s
CdfcrrlZuV8jLWDrmLoPthyhZT9yuPV+/ntQpRktqy4YqWmrFooFrUO2GK14W8u5UolyVFCH8iGU
bwTlqvoeK9T7ZnzY15oj7f82RwXMz+kuvVO/oBHabCSIzFZVTdzCg6e8SSrDBQ4SHaejgJG5WyZF
SCWpEICGqm2r9YIv7fjZTwcWQdsN7NxRvhU7a2dTAn+VwMRPnWk07DQ0KikvKVFygJAJg4vJEdMM
u2kMPeF/Gj26cWtCdUjPSymnS/dAqwy3K+fDxQfd3RZysUgAYcsSo2JQ8mEwwuZ+utFAQp2FqdFf
roSuGdpvsma3yRhXBg7tHvstWq2970IEwLPXYcJZIUnZsUyeFc+IEvBdQZk1FWeLbxVYVM040zEb
Qoj1WDfuH2zP99YulTE9XEOV2eChzh7gT59F3HfplomRlaD2z5rNM16yLPqhxxRp4b4D70gZmM4V
qnP0N8M+aIfC4xuSbTJOQXxxdE5vKL1NWFYfvPJdwIr3dcSxOsQaBrWkr6iOC6pHacE6r7m74Enn
Pl+Kt3STCd52TDO0WiFeyK43r+8wDRDpkyDl+m21E+LcvlSwc6091/SpvIGNZRPbPm+y0WzT56cR
knCG1dnQeKtQ4aHfcS7Dk85sFiVh6mFw5SQtEBIoAw1bbmqJ2zjMYxoFu7slfxCOOWiUq36E1qbS
YCg8ki9tfJNovkAi3fNWYKFQClrNgWzvd3KT2khAQoaVtoueRC0UgZzYMZr4GyreJ/xVg9ClVf1A
F3RwrGwuJoHy7Jhk3eg34CHT+/jlPJPIHaYz7e31MvAj0G2vMMC+/VZlH/Ib7zNPExgEunyjpLAL
HSaRuFLXpxR3fnoPQodsQ3r0rM2qjbHxk//B4de5hRR7wOaixYqquQ0rvbUFHAMPDXqZ8B5l+J49
qIVYOHSUe6EYXPMaob3V8CSTmtVHZr8zvFt6N35mA2A9wWe25zektlVT1+Qrkr80vMEXCBx6ow6o
FmbfYzB+6lTKJVP20TtimtaxkVo0Zm2tb1tRC+KOTJ+BM7nQnWk+ECzX+j0wYVn8M+9NTSTvILYr
HSCsqvJPR3hXiRfeHj8zew1YKkc5hNROOCqS9oSwRHNaxjgWMWrHt5lhIdUudGqot/YzOYlXIdf1
HJoYaiRXZIokx+LjvYSq1QkbxHvBwyRHYkoAuggxdrAOD4ltDMcyV4jS/6W3Cj7AyTv2zunMoe6c
4eMN3ZpznZWcVWzau/hoSAoPP4W4BYyh+Hj0dj0H42KDzzGEjLLOJdkugJU/LIvohPvdQHgQjPCQ
xG5fxr4vJaaFS27uGQnMXGXWkgW5BR16agpSA7aQ9lbxLbjoqGht6vccaHHUxM94NU5BIW041CAM
8sKxw/I0sK/2dsHS9a3iRKU+tzMY++JfjFt7q+j4UoS53VyzZZcd8T47eKx0/jqiFN75/bCdA2M2
OottPDDVwcx5MgW9grvLe+oBDngPbZNkXnzWw7IPeLS0gAKd7yfB36NAE+za0+jgNuDyygNyXa4X
by8qycvgo+yhd2D9l/5EsJFKzh7WJzBTjgybhB2TPJ8uMbn7Ow/B8Xyl94xyKZDxouQZjIh75K6r
4Dwhd/m7h6Ve0YONxoL0cz9Dx5MWqsA9nNkoqm/ZEszIwFG24DTC4cRLlmZ5d3TZ9D4VDtGGG9Lq
dRDCPc4DehXE7SBKx5iar3PVlvHwNuxGLaU2eqJjMzyRck/KB/05EDWKr0yHvTdgT8iQnc+cE+HS
4XY5bRGsFwIkUkrLfQxX5jIbyM1kRIr772XNsSIYWW2q0QAA64fzsto/UVlJ70Q4nZqAqpIC0Qb5
9BklIqyibaVp6QLJRMY+lg0AOvRubux9WLoVDBXqc5MOQZs9i/UPcpvRUJsxwmiqtWP9hbgU5r4x
81wiS4AQsR4r9AvsPU254Xqy1qfgMurYVRfr8+NrkLru+iSCS77+gZYwmDDmKiIgx3rM5zTv5ZdL
OGSazSV6JefUO1iJ7vN1jv2fmbqWRypjmN9uq089vLU0v4R66h97x8Sw6/nLjz7X1V2gLi8dhwaJ
XMcy3P1uzJwHHN4uPFqYhitaFLKqwQZHfhFYLpYEjLM2Yn4TSdBHVOunJZcFkCzrT2PAwEVA/94t
Bxg+NvUTnDmLF3lkv2XFPtpyfJ2HUBxOg87ti3HewNOKX3m9cvp+gzGwcp7Ya7/g2TXMc0Oa7Vl9
Z1QIXPfIujVj1LOahIePWa0mxQsLQOPJKoOPDXLnIU7k0yU1piFA3BOfagLFMuMZpkqmKdUK8dpi
5W4h0ZtvoDBs0NHEbcGB4LzVQ7mxZ/148fKv5wtwZOiN77jNvnIfH1IMcAk3Y7QiWP4qxIcCJCnZ
PMgfT5Cnwwc/KHXQG6kTO1A1yADLIuxvdGXzJP+iZWt3xIEHB5mrW9F2I48ClkL/5UqHQKoeVQCT
CH5sPPdm4xZAaEqy/7qoI+4kmjKPReBcSKmtKglLAoIhZ1pLmr+9k6d1gV+D96hwya9l4XDZnwjA
eGpiQDKYFhgn62UoNd5T20JLWvSy5RebmorL/h0jm0QR59VtKkPgFDaust7t0ed3vFngJ1u+oyhq
AcEr7k7J0yozkHU2+6yxMhKTjRBcl9fy075cD1nWgUTIcaddTVXgJishUZXpO/geayHmgmRjPkWi
LUcgdmKDf81FT1/sTAKybE51EcKyyo5kgyXLpABiZR0BNIj5WYGqv4uVmGrG1uJrrqSJsHbIPzpB
zFZksOW1YtV0TtoV2eGOkYxjGdnKkyIYkObUyGLy7iF9dhkbrEx/S37q3BqptqU5eP2BqJ2cS1Ic
kRCPBtS+KHb6BU3IxJJ9op2C7nuVa0wfO4fVzqBs37hlX2BwY10YT3E+DGO5aEj6fjpGWBSUq5dm
DKeGddFk3f2Lt3AtBXGWE89lD/9U3/mj5IYgYQh4Bb/sAHDFeDew3PKhCzukZzSW7aaEJNz8ak4B
kPC1EG0UK/el/ETtuKpFR47UiYXsG81cnT2xMbMhJoqfDmgoljd2ezhbeTeJJgZXP9LrsbdZGRs+
2gE0c6VHb+Nrqu/W/3YXPZ6b1fJv7TPIkw1SZlwDPTtHkc2vK99k3znLyihfpE65TdwbDK2BT+8E
F3tcT2GkX89cmjbt9lob4GfpfZZ2Oeo0NFb2yr9HMC3GJzXfB76Dl8RAjwv0PxT13xLNSGKEQMdO
SdjhNDUuStaR+nnRdH21G2XCFpPhMASw7DILlJEMKxfI6aQBLI2f1iJKXlIVuHbpNbRRaI7R3iqj
mDt/o7veFidqfg9BxkbjmlvrKvJmyEEfhY9gUyOIMLY7FZz+OuBsIMp6GZwcECwlYeWsxKXn/PsR
2JSJlXiIDv04Cgi/U9AaOPunM0DkeXHL8Ev1AKSjnMQz4yaRHivUW7MnbQXKFnvsGMXSIOTc5itc
Z8oH5TOAb2QQZ3nolBjw/AvqSo4vgzDIfDccLxlQBT1mpNWMaL6DpHCQ8hTUVD/2Qz7xakXBpBqj
ml7aNIQCAYhV5gKelhk9UNCY1DQLmROXPyR6xPjXCVMXkece9YkuGZ1UHdzxspx/KHE/udn6Jxfb
gRw3ZQqe19wirizlpJVJzFyr80h2dQm9hMGUiPpWK/xFqEbYYfdowoBwRSzZnb6Z0E4IsNT52bKz
RYsalUI2UUwnjdFsVOFNvUGbJ/8eGfh6v5v2UF+qoNCMVcRUoH0E7k+mBoiswfhqd5Q6+VjoUqWV
pUM6biPzrsTaabfAbbzpdf3RsSS/WAuexYqjY8KSJGuT8SlTrgwn6bh0zuOiDAX+pQ2KdEF5g+ou
QQHmXVPZwTzlxnyTP2U/NF15gqiuI0ZGv6eAbrnldFf/j1oxfv1ZzuF8W5AD6XTW61JT43MjpWQ0
EveGI4KJI+2f+VoV0xgbX1h7ImrG3SQHmDv9W+bD+c5GsP8fU5tosxTWyPcU+YUXynt1Q13Lyb4E
W8IgrFbJqxpSIh3/PIp0qsrlMP1GCJhemtiYjmF+pJH2KTshpGAdc0NJ/MMMj7gOTcDEVhVqTdrX
3KvmOpaPUocZwNkd3nU+e1MVab8Z2ARNYeb6xU01NYz2cSAYqbD/Vxuo3XmIbuG+VuqxBVf5R2lU
zRzKH8C/IgBTteFWII/4SbzKtM5XKrskz8w1b1FafixqOYM18QQC9T+ZWFVk+YaS8tl5vCrxnD0K
YXJPqvoye0CWHZv74zx+h+2TUCL6/iF6EAaRYwROlfpAdlvnXxa88lhTuY7UUrwd/vgHeJZv3A+3
tXoTv3GQRvLqWFNV4kefGFDc4L5z+hvEkv/HIQiD0jkFUFknlY4NLi+3AHArzCe+oBzOJGXO1sj+
GbKTxDFpAfjcV7H+QxsoMJ77NTmREvYfs9ZB7ND7+wQeZgL/E6H/6wYgLdY1sahE9T2NW7NiMwo7
hGG19fZ32B+NLQw/9uhXGrQJeT7phS8I/d4QnslH857r1n2MtIMbGIWPHhYhMX4Hs75JbM4rnw8Y
RLhm1vobkG1ZYH+T5EB8Q3lgORmG8xuNXRnpDyfsbNTa1aDExRVQmTkHQ0gvkRkb7Q8d4jIL58kK
AAf7/UlcfJwK8YhZ3ntjW3iI3XuJydZBcuF8+7YHvIURu1irrW2ruXYg7bmYdJGm9+roEHyyQ+i7
Ul+ywB7FMTu/dm4fOYbyBoWd9x3gnTNn+FBFX1VbfM/XqlQfspHvXJO7MMn9viObzDuENBIwAraR
sz8+vtee83fo9ujO3BWzCwZDEoePu0rCfR9fvfceHKYkMe496LbbpX8keQrNI+4EKqHQljPWPm84
7s2BxqPE4Oudnb39Vuxpn53J5vrmTbz79T/Wq7q1OE/c/bsd+jMQScMHfXdYWHcZJofVLI7D7OhJ
JteSoUmcXPvtf2gG04Y9+CMQxJAKYYPGwjWbeagsi/pPsZtzsOblB9hRBkLlgPSbv5o+eDFUYg0y
z8DHMi/KYyKsdatspI7ivj2CGWr6tVpT0iThGGZ4MiB3Et52lM9zNjrYgskZeDzTHGlZt/boFg+O
18oN45aiRRovLyMER2O+9IQYaXQPrn7uyZtDTTn5LEFV2vwLNKHmMp3kWB0vmdnjs9bPk4vxop3h
OgrkFEzLttdBcv5B8Yi23RAZPAbMA5jePQtjC1yGu5sOQxnr0X5EYQhFr64br+DVrdXdnbuGZNl2
Q0iYku/9sO8INe4pmkbG6tKh/w5ZPAmfFfTQOuHozv3gecBokXyLICaLdKjEBoZ2e09QuRyTD6YV
2VunvLAWzFk4NgQk/kdNdvn4Rw1vI2ojT+44qav/JlwrsrP8SXI4wqYy+2RfR95qwh4iOGLZ39Ql
e5HXzrif9IA/t4GkNFnLLELRc6b9LaBJD8mcNc0VuIvCcVPXi6JO20n7WutMJX+/GpCaTA3e70dK
kPdC1oEwxM9W+tGEBOrPrUPHv4zWMk+5xd4631f2rspTD6GXKJYV4GIJVFbisikNUWHi6IcTFWr4
WJOuiS+pjrG3KxuWHRu3r1iCsES7oVxGKwNOnbFnYPR4o88aQMxxpwjgkx9tlGjossgxuq67RQk1
BPtUwG513Zex0BoUk7oNiOGH30jgQxwk0QLv38A6PCaZBjOkoCpOC8Zke0HnIKSWhSk3t18n6LHl
sxPLVABM9sZOtM2YY94OmAX7ZoM6KTF2Yoir7IfEZKL1m7mJGZbnqNDN6z3LJ3ANKClEHpHAtI8q
/wPupuxH7iW2+ROjEfASWlsXnC/TD3w5+ZgCKsmK3/ZVuFbpar9CNwFHyNAnmhuFZTj4gOQDoLwT
SPm5WYSouhcFSxe3XeaNNEu/ggTjRlD1oAjNHuoLVWbuyuS2Xkh2TPPtB9Gnd29vo27NDZn2xFBO
L2lvlmXuTF2IHOTGAZMN8sXx/xU5Jam+n4b2RTjK5f2E7t2Nh3KzNhTDqGBNDQF2IN3ZR85hhhnh
dPE4SsLUmobYQOtE7fSUsJ+OHEkXqc33cvlJlh888+gv2IKykMFLRDd48UacnRpJDw0IggTLeaa/
dGYmhhHEeuYXMNlSbQFrEHYZRmHxh7dHvNPWObOTLJakIIz/CZe9FMUKsTtEHFNmy3EZiCPNN937
RiShp/b6dYRRwmt68PPYM7AVGZpefDpPuUwcZ7A89/YojMmb+PYO78tfluReTFOSjHbZTQFOi1nU
amZwguISF0/qu1yx9xD8zyJ78JQpHiOcLhP8WBSIG83Ws5CQKrV8vtzUBSJmkvoxw7Fv7pajIKYY
H3kfKwu3QVQL/6dVmhzS+f2FS7G3echy0PITtIm0vqXrLGMaf3QXeU88dXeh8VpAx43ZS2EjdDfZ
6fXJbwIYnbZXF97AH2mtgKlP+DwHvwSpcOroIG8OVzRkInj4Bn+tUThkBtEbpaseN26OMzRRn/PK
QJth4YFwQMA1jAhdVTO4TMYQycUg9YVuYAO2Kd4VoHw8xZEQWl/dQ6V/8QzaJ/udIETbHwoGkb6L
iJSGtOp29WXFTDe2rDkw9HY1Jg96rQRu96ZWDcYoMCqRxomQ2Ww59BOm8cShQiVbbQtMM/BEcBu+
NNl6tY5ShRGFWEx6xcHxqOehI4E/QL2mUhl3jEYWBn7dKdrYe1Z4IAYeQuSlqgW8BDU7RXxY7U9O
imlVXbad3DGri16V7jw+wihLngvOFt9fPYk94ce7swOMtu1K6ItjhtWkgGRJ8W1u2o1yJkQph0IS
5wXviPM2zEBSa5ecYzseifJIkiiACUjpvT1PuZZOQgwGXdW9cNmA8tsELqxovYyuVozuChD3DnMg
uS2c9v3lIDcFEqGXbmucZt17N0/mXN/r1slDi3v1BTwNS90ehiwAStxj1YS9l/qc6idfNHSQrmvR
IwRXFsrUEeGmB8yJ27aL2uLDMYZ6/Hrwzz9Wils9cprNRsXYEu4jyVof8XUEWg3we8AqXiJtPLJ+
ESS93js18yqjzJHgMSt+58forX/oP0iZLYShvB8pFz18K6azo7TkZqZmuSUNC8qgAzpVdxrYvYf+
fMs/YwnvUnvu5lkyO5gz8N0T4mM+JcEylWsIqb9OMQdi0M4OwAixFaCedpJMl1mc13spEp/skElC
vocDa9LVlVvsgIVxlx0Oo1umXbH06b9A/u2uUPUcSQLC4j9IblFJbPtvrG2k14yBswucSQ9gN6az
c4MBH1XkDXXzoX6W+slYs+9geF/l2t7/wqZoTjGw2G+MoBSHW0wBxhi773E/mLdtAsjZbQQIJpxK
VJ/0GmQEvV4Uc1+eFsCQ7sES4VMcgGxQfu2UpUzZy1Myzq6RmwoJ8l9h19LseOFEs6s+sNDQ526K
5junfWeU0Xk7Qo+xfpDGHs1ZrGgXfrNhz/WGualyGzfgq6hY02/Vyxo30vOxWyn18QIWaTA15f2/
zaFt7VZsmwDWrd8hGr/mrAW6LTHmZw3CT0cGKlTUFeiJrqlQVubJYd+XoXLNhFlMsVWLm05XWrhT
wr7afeOSfMvhmw73qGeuxveDzlnWbIoIf/rIKnZ9lDZ07BO68hVqASZVC+py9eJ2g3jNT3hEahYz
Xxyfy9vnuf3A3NTirzAMkB0Wk20806pK/wHiat2QB10t/kc9EGXxWcFGZGvUVOyGCvTQ/PHciXdX
mRNVW8DSYH2AxKjm5OWynavJTPHBk+6cIubDeqQQUnl4jFR+JTn7BGmmOXs0Sg8uiyHBJw1vqerU
duIh46GxXXHGoobHCcUG14t8RKK3tfLLfpzrmyECfHKu7Ff+Xe1/LM8Zp7FKBUsBbsXtnceAGgFr
I9oBJXYAzDy1MB2AB2wKkF9VkaXVtWx9lXfrmrboaF+gX9qEvjHqW2RUXSnNHF5rzGvDgMCvhX/p
OgzrD7xtugBR4/xaOxqQvulTQOb8f4Wj4phKXt1dWh9UxpylTss/AvJ0KsDtweAh0OhM4DGosNIL
othhdisSaBFwjXoWu9cnwgpruSt2zLYqVxlrpoTU7LCvjs9Ap49Sj/RHDvJU4MqxnibwPreFEm99
UGEMZzhUUt/OWf9g1dO0r73/pW98/JsroncrLgvft2rh1yCT2wGgQz95FNZR317+YORXaBgPO1qk
9pIzT1v1ph/fjqjtLNrahbJ4fKvYmzojl01FMSa+usFGvktM8b4El9W3TP5o+h0IviNTQdJPb5Fz
XsnPjEgiuGc11CxT3yG+B3ilbUPY8atRGOV8Sv5er5ima/XH08tXhTJeOrmi3+6C8Fb1KvtYsJK5
nqPLk9KT3HU+ElCjsA2NNcsJI0pX6LtFwxBqPOeirQvg4jG3JjdVq26ncfKIf34d2eRqKBkkzVuM
9Ac3O/VaIcsk9vunIY7nFAkqwk9G4cTRRGRx1MPU8dS1d3iLjlSWkH8hId34B0stnzMMZ4HW2bvk
YvxSfm1m4af97dTdNawAUJ89GUsWRRGPJ4owPcgZNhvsDPkfn3cKTketG5pDR2l3qw9+LTX7RON4
gAPreX7dVLIFtXfGoB9MmUSEr3HloxvRKFWEcKNmJkTMGP7nrrwuBKfOp/s7Uz1GA1SILqLxZy3D
RRg1N1JH6kEfcjGKQHkcakvy9XcWFj2jmO2LmnkCcQzVFel/1apJ65JkT5bP4vuFUPYDCT1LUS5U
1/5k+sg5SZVaZGJns9IK0IuxIFzUVdHulQun6gVuUBsWfnLJQ74AuQrHU1VJC4kgVc0CIkgNZgi+
QzerxVtL3BPh/Zt0UNP9iAQ17/8JMMlsNWEbIfla13mTla6AtpjLgo56O+4SE2s3232md2Vf0nDR
IPUZo4EnnMocD58sKWu/5urOQETsfeS0L0hQMDe55+YBRy5q+farCalL5jYmLzsknjQA
`protect end_protected

