

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MndbkmQgTx8/SiPqHkiZOQc2Og7HsnPGv6R762YhZQlkd4u7VGdD8IGkiw0uWRUu6oQdsfM1OaG9
WPWL29c2eQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uYgUbAMBWB393Bxd1Uwwk/JZMU+8OgH5Ff0hIkY7hTLYcp2m2I3qH7c3ic4QoxZ6Al+voEtVdAk5
Bix21hRZ2Y0am1rrEihQmx4ePyGPrmsSNCEQjGFVhcuS2jdqxYRbcztvxPnMnmA7z2sGgxlBvDca
2LUCcUabhGetrgqLRPw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oqgsGo1FvkqYDJXZwYKAlm2GwQouVHyr3oWltCkQfy4eDiq8e6dZtMYTvS2OptsCXxwhnt6dpFkV
aQPwWgI4M/EeWoFl0sJqSpzuKxw3clkzso1m+60ALM2kbDdmCRiPzqUp/agesGa5v97tktn3T6EU
BgYvmTcBujJumX/2YXO0JCzvDgj15zfmbIwFlBOPlf+5lHj1TDCyJHsleQSR9Aw+OaqgMxpV4mhY
KIV04+MC8ksfeSYXqZM6GbEdoTuQXQAZJzv3f93bNIadB93Qjw1ApTq3glmk6F504OeL4H4uFhb4
yrLA/+YVagpERJJyxq8aF8jV2cf8ecUQVWApJA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ot1qpsZGNYyIou1IaCBBPbZ84syWy7TKG1f/JPbtBkfaCKsScSnESpPe9sIEyscYmg2MtRaPN7AW
pPElR4ydaedMQf+P1JcgNOAfE7pZRVY8nidFZsYHLk1yqIYc7kZjeBd60Wo5rAwgqRN5Z5tVa1pI
Gjf6BjkRcJxSd3Tu227hWTzk73NbqcSK0eUT2OmuNYVI9IdHb/PF5TW46MpIdHW1dZegcarbIwLR
bwe2vnrYpJNkH1MPBuSnZN/mmW0kK15ZEUBpz6MZhQu6b5tP6+p4qUumkx43xvPki86TqWxHvjKy
yulQ+bFIKH7nyGHyWzM2izLOJ93wG0vdK4K7/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PbJi+boZI6/u9MDnTENt2Rcb6pD7iRjIlP6ME83AndD2K/54TLrMalMeI7LTsr97UwTKUFhzjLF5
XKAzaDRI1Z/F0TOStSdDbTq2p7N+l9ugTgoLpWX5Yq3/aGpk6L00r2Fm5gSOceZIoCI6E6rvaEZq
2fE4A2nqlGPY7nD6Tgo=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U41YN1XD2lvq5ZBC1dknnD/8+1FHs+DzbJIA/qcqrsNBOVhBgQ6QTIJSI1PPcUQpjrGr3zoN/eN6
Otg8vQ/qNLepw2AqzWc7J3PGDNuxYxVfXvNgBR5Y7czpYRo+g0OQqGUkdOAQbsfL3tC1KFD2mwtB
IwQwjBoP8jx29oDmAEUQ9T7Iv6Doit8ulo310hnw1KbbW18kAqDiczZLAdBvdWm9gmXduuf/XGv3
ekAT/xoctRBzyMw6/KLSAjnx7HBmWiwx3WDkoPfl2jfgWMmneVre3c+6nnHhmu+fZbx1P8zovjz+
gTiE+625Rd6WtxpBJM5iJaRSzwPBrlPDT72Lyw==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nvjVjtChOYYPiT3W2qQsbIogwQPRl90aNdsik9o6NVpzDFwS6AEfklc1U9kUuyE5ZqdYMi2XL264
4VfeTmZOGLAnNXvF+1qv2dH7JpycefgUtOdavuUUL9ES5QLHVP+imBnabbIyNbOtVt6lIBXhicmr
kwmT+J+dRdC2FTZ7hZhDfQRX/66b033JcoXE+EZj5yf7r6DC1f/IWvDOHfISdsXcUdlU3PbalCDy
94/1SFMc9/N/dnqYuxDczKydEBuchZeIouIdQu2vtSsoO9qNv8bH9eR3vXW8VzdH+Yf3W2d/FyMr
rwEaWhDQ+Ftm+RGc8A4ZXAj8zW/r/RMuWf8/cw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
brCdM6vu8hnAr06KwbGI6icCY+Q4rv/VITZPcy7/Z6aDlmsxgz96AuAPZVs7C2cafXg5UegZek1Y
EFhkIirLmjoPsTYAkmrMf2l/v/HwIusgZAU1KpriPLypXgjyuEXntQTnYIx9hNjVe9252xXf36vH
/XDflv9Z1YumzU4GMmYcHJiz5UHFxwk/87AWqlH6Hfn7fhCGrHoz984ffImxmPHL+cbGdzbcyh+v
kmF/lckbOBTnBfu/92OknPpBQFhAw8ZFwNyM2v9TJyZTwHgdfLLgG1H3nipJGCSh52D5OjoGsBQz
bXFA1ydpE9R+BTksgUhjJig5Oiv3yWHuu0PIyg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BS6u5oDcP7egGpSYOQ+FbufBNbtK7LQ0P9+kszA+El74e/Sv6S0VyssuMGoaSJ8MnvgdnMFwhjxU
mZKo0GLtlzpNaE0RBile+d2hI8zREBXIwJcwXHDJKOQadE1wYhW+zsKRkjDgzGjLDicBbCi/grvC
r2LKMhUtHrtscGeT/udYOYiKOanwk+8PtmKh8shfZY9uvWocb8mfvEN4lwpxkl0c3c9X73MofBU4
9uPLacxSDOEsH201WRf+r5psiNmY0WmDZRFtUVIJwa12M73Ug2NEF3Lctmn09U/EtiPZHXEhFxQ4
ilXx2ACgw52aYJnXoGowv67zfz1dMVKcT9W63g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74240)
`protect data_block
b5s4xqXnXyiivyzy3zCBbzDVEx4+qhszvWTcRVQEv4mzrCj9LUGmEzRS3xPRV9KNP0vdDuzeFotj
dDwBNtnUHDDjdPwfe2ZgmjAeStte6oeC7xW/y5YnTwk5CjbPwQZm69tc0m7jSykaFu4FKxVEF+6r
h7sgrGO68yefv8WQ6ceWAQbcfGKkgGQUQW+4oUoKqj4zh9pJN/ieZDkG4sRQQqe/4HmWsBcj23lY
GhcHF/Wj7vunvaN9z9/1XALFgpSAlTNUlJwqmc5uuMgsI/ioO/Sr+E9EwZrXqMoxiBBGYFEae9pr
lFIMhduf2xT5tJW7g8QQTmlMm2wnjKLAfrpe+1ht5kTsACvUw+zgp5SdPRQuTorig9uEoA/ug5cP
+cFN1A4MgVl7JDNLhrjELncYdhFZzNOlfI2mlE+ZFvja05L/qMmsX05tAQqlJpC8gfbSk3ZvPv1A
PBPt/nGYCYTeHVc9dH4FJsjiOnEznjTyHJ9RUvgYpp1+coETCBgePuM6I3stdZ5MiuQA+7cSuDKn
BQ3TaOALvUjLhSg0Z83qYJnl5nnUkgaRGdTkIAGug9GLpz4kPwmGX6NwJ+aPZoORX8m3bXQaJF8L
oAIJWSdA+yC+9yqp4s7VvU5dRWJDcdfiyfhls9AQKrb2U0Bb2yq/6o3L9hZQ2Jvzjtj/nPA0ju22
i/V/3WJ4sgJ2x80hzI+3TSPOyPrORZUOwYr0PtDhY3FMgt67H4kBexrYN4kNxiIiX/pYn43IYAqi
y0MRe6iXeHr5OXo1ZiL9FAfZ0G7dBHvDb2f1YYwQIfBKZypG34tZwT/7YsXUTVnVS1xmwAItyD4N
pPNvHFR65UyzVxOJSsoCa+BsLEw5P7qE2iul4FAzEaf8lWFORbR2jySXDoDJeXsBWpQUwnzNvuAp
uMrf6RfM2/5ezCUG7UCH8Ky53q/SI70Fb1bnO98IyqGUmwV3FhxRNFXdpSA3q4EtWWgXwT29DQf4
QHVsP9LipA6luJsv57ZXbOlqjfbnPAJaKsEBm81IuZEXjr88bdywOgReAi3g8EXdSKl0fHBYN+Md
E0pZvvRhnVvfO7LoOz/CyWWV5QnaOWUjfAuEYtgfam24Zks98a/mixdZgS++Osl7vN9WizGjBHcK
YiNl57YB7Xd10/6Yna+BUycgwa3WwUpguXhHqUgfwOE2yFP7Nrz97a51wEFmTBtQNcPLy02iLUNp
zfTHlmCA7ICHbxcurb8mwyPQZmYWJmHqyHyh0BOuWzuhjTM8R+Gpnx9p2qen2qGvtYwiKi3f/mOx
aHtWu8TPzydkhbOzJba/66YOoeM8E+k2prffCmZxdlSJv+k2d30AjfR6ozvfWpgB5VzhivuejyWK
67tOF4tDLPwrCs5gwh72X9r94oIaZxlvh0qoS4QWEaiATnosULqgtx9GXHmlzLAa5wJ+5q8q9rw9
XnBLyvIJJcFr46KQ9G1dwN6zmVP9sJuq45cOEfHxymWCsMUP7UxA7nCcV9YBqZPFk4jkXhogQHpZ
RklADXuMUitV0UTWee3xS0lY37fK2NQWkMSSPnptRp9tey69M3A8/f9iZul/K4cOMbFa/HpAnaxP
RkpZtp548ZXEaa1N6suLgXckvIZ/TP+RyKSRZmuchLmu30zWJR5slpASf4nl6oOGvwUU1iGyHRSL
Qxntnv+Ejp/uV0LNzFYkBhxTnAV7uvZKpu5Vf3ryHUEqpJMK1Dq1K43yjeVNz247FTdURmW4oqBw
3LcOmymHngDlnb709z7M8tyouhHvUeQCzNTvdddOMQaRjduGhK5MMe2Zn/jmHUfaCy1pnN+0ULDM
Z5Z1QxZZacQDmvUqtGRv73Rl+rjnaMn9s1gorLatH1vCIOSG9KfnGbSmOta9lSOU2DoHQSm19mWS
ru55jeqtSDhicr88q8Yqcr8d0tbx0/2XUqI3IA3Vg9Lpc1hqad/SBwXlaR37hUxILmCXGZ2n5XhC
m3byR/89RUkzOhjLdprX7wrZYYKjQ23tQp4csuTvBhZ3nxi3X0at4upgq/E9q96bHnJ+uin4wLl/
bxcJEM/ql1k3F3RxoKiam4dBLmNkijybBFMrCCN43uXjfofjV3UH3LGi4QNz7Y8lMKbyYY6Hpx3B
Cq67sb227B/wKUtnEVNSqDngOmU9RVpFp6IORzPqsBYGLbVbT2dm3khnzd/mfkI1MuNfeswjc7xy
rjsJ64Ym1b9R6ASAvZ5Iy5KoqngzYSvKlJv2KPWxJZMLnfLuUmZccS4PlaXOxkg1XVjcTAWCzRPL
DqM61wlByzonlAen5LKajBs0+EMBGr457/Rm0gU1ix8+zGgg6P4v1h3s0jSjnRTxpGqv1DWh7N9n
cbq5qxxIPLpW4Eoq/ukZO9GGT7vCCCX9lMxeboVagSSrBdGV+r1OTNrxauC3F1/RJWZ4Qs8LhOWs
cDBhEuau7yrhAgfR8AEx5evJwNLjMCFDl+M9nR/FRmatFo+rROktIzi1TSKgQYvkW70MdXLmfLcc
zh5SCByNlrZ2EaI2OS4tPx8sAPtsfnx0ZUwyMhb8Puk5kc2ZjU7npME8VG3hVOAsa3sViySILc3U
lhbNUxyBt+XtBR7xdHD0rIVzK+TfqMbj+Rw0XQUQO3Bo3m9qVCbWijJtWY93NsDWpOrnVacgNOa9
QYi/FHvWazu3JLu6rA8fBhQENnujkojoOTs59RnnVfGelJZVucFQ2uvVL73GkqaZRP0QkfZ0zfpl
nFsvq4YbTsknRoUXPhp56BIFRy3OJnWGkBqX7TdiBJwYpOoIEcSABv2rl6HATd7IWZXEAa1TFOoJ
ZqZjsRNm89Q3wRFYC5gnRKnWdBkaGIpX7np5s6bxc94zjfD0oRxRGBNWULh/n6Efs7dPeSSH7J0I
WF8lOYXazwTTwP1DQDduwrOagrFsb2VnOrmpMouBW2dXsZZZepSsfYypINOQN7ltycncyFFmZMbc
U3iMzQWM9xbq7KVrYJaBPDKrd9W1XP77yRE2Iy0jZuLjN8YD/YOkvAC7Xbjx+bKEWQaLxljlFuMR
KwhuqhPSrt2jpU0E+gDw6HmU817HcWi5FYj7hUplRa4tS2YVJWHqJBXkzDK/Gzi+vdLsMLBQ5pWD
XzHvd1ed1jf/w+e7mb5aSVzMpC9yIkjpqg3QhtlepnDc/KSAe+xOopLYsB/frvQtl5VsQ+LskUdo
McgIMKXy0oCgJ4wl0rMs9y5JmaOImDpAL/NIzp0fRckebJSa26I595dvhdbtwmpUoilwCxTtlRJc
FLTwlUgZQnkXtS2iBFCD0WQr3Gzjza6CkEW+EVGgx+Glzq/UgpZ45ZaPp4lkY6eygMWClJOYqhGC
mpbD4dD7ySZqkyNQiGyfiycp4DoqWV/7t0OlLCHHETuwLOGV/Hrlt3iL+y+f5UmH5yePLmG2y8wC
9W7akbGvJK4ZaKMun2+JR5RAX/JqMc2ukh4eHT7Hc6MNUtmuI+PliqJ1q0V8gfeKIEVRqGsPvnFv
eh9XaNU2gpwxJPmZnQGlRj0Ocq4hGh1No+uPOJgXQTftYUMMB5aI133/tiQrd6zeIZVR6MSKMa/P
4vWDNWSCQbQrkOwXgBXlfOgS7hOtDJ66kHy9hI+yS+Cm1QJsMp+lN1/FbJ2hxirGZbiRfTfxGCoY
oo0kCSpxQhz3UCNS+A/L8aSeBq3+kf8F5D2mR2Df/N3R76/r403hvX1jQnU08GfQnsyC+Rjp8mWh
IA0DihM+ViX8LHSL+TWW/udfqIi0a8/a1wdZepbFkolzNZjHTP635AczA6G8QRJ1iseDPTmvXSyd
IinI50nlcRgsI5AbAn9gpJb00HvZc5OTT2xF5sHnjPsbmyjw7V5z/w1K48nnk2aCaOleJaUwn/GQ
XOREfOcNc6Fa8AzZaeJwtMB7KOANVlRpcd+4OHfujd8u2a428AT4KRLC1vhe7K5tsSYqoOvYn5iw
1HiMOMtzem5+wT/ZIpiCKFe9OXkC/a1ZC6lr+IJ0ipPu/RaTTS3OGM9Bdc0XeUNuabISjCcDWwjz
A5rP7H2XjfDQsdkoESxXQx4BgUO+YD5xL5bZpf+PDM/+xWEBZf+4XW5Yvzn4ei9av/V0ceIke4k0
k+T/IGICo6ITl7SjXZfpL7IjeHRPxNmuUzzzayTrJxmrn356eVoq6TnG2Y4TPBuDoosEUxczm+RB
Sq1FGH9vsrv8ZjG8mpaZeac3iKnahz1drV/IhxGFKvLY6fWvMySF+X6JEnCmS/885sdCJEgvhkj/
LMvsIbMvRG7h1HE9aT1GFqM84QEvbmvxHvafiFsomfvhuyeD6m3vEpVZnBChnuVG6BuW0qhG0OkJ
MGk2ShaSDww3oqAZPIDuPZHSwV45by/JIe8Zj5pmXaBL0OOoaYLh8KYlaEESZEFD1lkanPYDeeoc
cP/PcvUtox5k/+U9PRwmrkGPv40+wcTSaWnzpEJLz0/oSPuZf3t7estnITz/JUPEUsecytxxpzG2
EEIVl8ktkQ/B4UuvjmjzYHcBAVfv17duttfAJTzSWbcwxn7BTUSZcI0B8P/voYJ+H4QyqdpNmKyI
hF155vzR2Rw7KQ/svNSDGFmji2r4jW+RlLkvitmqXoHRjRvVpastchA2jsc49lABX7/x9D/5PZJB
LU7nShVi506VZTuBaUJO3g2pt8flR/esWUZ8ealizY61npbz+q2/XQvwzo0fs6mH7awftxgOO8d9
NtWuV9Mba38+50PTzmMQy5HAmmPoGkLgNGdCKjJVc9V34yCmDTEhOZ0XvcDPqG+ksl9fBms70o51
gcypMAV3NWcsofUcHlUn6dutor5TbQrAj+TgJ9SB4V+otdecv6ijoCAfxs/auAEqxFI6g6MakGG8
0I1WPX+aE4WD4uFZhRYybgnFB4pSND5BxJuAkMnqJhvghpqWOdliLl95BfhTTkruKo9A8Gl6AhJr
qyo2uwYWjlAFBqs/pmJ4o8fo9UcqOy+9xKKelvVfuZVoX/STNXbBi7ai1P32SfUVW+vkBnhtcUuw
qAyoRwfE1BBpSeDEMtIKMEMv8/UXL2fTuen2KinLgWggGFiikwmeblsP8/Qi4l7MN8+Y7L2nwI+T
FbdP2Hy7V/oqRdc3POp+uCLPaNXeEDBeJcnca/rbiHRgsKCVk0aQwvhwXi76ikK5gFMX+HUt/OTW
NXzMs1IvQrRMbbcg4+5makwoTWtpIt45pSx8ax5BuodKHwpFEosXJaGLESUyi/Z+GB1c8NypwSro
bRZdZFIaqPjKZC3f0WqCs+bwr5pNjhLufrO0suYkbaUrExN2/Bq6Qbb11xZawk51Jgoc3wh4rPFa
rEoU0SU3LE4G17cURqJpsLpQZ4LsnMKPiTksDsUklwvSDdUeVUWfvT8luxf/tw/PoUif4F3vuQeO
UWQTjU2eF33JXdmO31jYdfh9YWCGq9dgYKBPMStocr4tToMy878BobqIliUqiloZfgswnJcfw22m
msmWz+O9ErXq3sbaW5aPj0CNg1F8BsbYQw72F/RryNoUdIDdng1rhQPj2LC6eHl20I3rAiaSTgJb
nLTiMt+6tvql+fyDgUlalK4OrMJynlcZfrG82Kozb6ad3myrtTsXJgk/Y+X6/3lxiLfjZTkbldjl
3rmhFStAzuXPbbL/k4M88gl1zwvOmb6NXHzYvHxvso0LnYgkzOwhNZFW2aqD7KgoEKh2uRnUQgql
90vml6wHZQhhkzYQS+OwDFhI1MPm2ihPn197NuhccnMp/f3uE46ThvDcx8PE/QCGa2pojj1iNtyE
ZYxp2g69AyAQbasa+kPfRQvUhhZcv7yz9ZlHup58ie/JnO/5sg1dG7riHh6FwhDeesDDhP1rHhbE
YvhFESLU22MWS8HK0CJ7cnn4AGQMNGSrbg6s+vzYf5mkHgnd2c9He/iKsgfwUCSRDRR7o6UNwCzF
zIpb5juIdD5VRy7EzPkadP2jR2zT0VR2mFZyLxuf1HUScJy1FqZTutnVYm07bW/oVI1OxnVrzHWH
7dBYSJtb3EUESQbQfPAEs3vND8084goqsH+GYiCqHAtqv4oHcefJHDKLpmWMCJIw8PI+LUfAYQjK
/a4PrBkJLZKyCKiS9oDJInrKsmSY5Bi+T0cqWvIKSeSXiQzacBRzi7ZVaBXFZQeeTY2dqgbFL02h
oEq6iSjfu8iKsvK6+nv6YjCVV82OSsQ8aMPEvph8Eh3HAr3neh1V9VbunJKIlWyTtPVen/z9lk0P
xfUnZ0hgUWZWeMFKwnXxr9+1tm2soIISN4W33h1YRZCYe7d0+jyVBqCBx1ZE+D7/FWWQdT3DF9eO
M/YnEVcnSLqeSwL+1TUIunVi+MBn8JbEZ8+28T67GH6qUl4az0FAljLXt+JKJGQtOU+UHO+0qvg7
bH6kQydImPdONdUt76vtUto9dGfDl5iQODvByDM88QSygLTdHQgie5G6LuYPqdwJCwwvDIbFwUFp
zoRDbJ4/4T7St8E4meV5H77NFaIRffhvsMtXbTavY53oloSiRIqkjdcNXrxdDr8FM8HwKOnzwvw5
rMbXurPS3ffzAm67doheQFOb7TIwiPlhsXkGejL3/pZD5Oyb35a0q2STMR/UybHhnP1wlt9ZbP+5
Xl5M2lVEIccYybk1mh0Zhe4vFJD9J5xfD+fzqnybkI8XIeXIzkHp+6rc9976ml3OJQvoj3r/7jMv
dYpmLwHPs0PysNnQLN6O7Pumgc6BynRXQSfP98conVUpUqaVTJBEpXNTaBOrBKlwL274GPXhv8Xk
ld5GL798byR/XBgxI8L7hn0ywA0JopucF/3ovdOs6C8wEMmaUXTvhPBLnpTrPdjVq2RZV84fbqdy
JLxAzrHhrw3AF5bqY2PYDlGu8d3qz/dTFRFipB3i1k2qym8+YJHq/imlSL/wAaHrnNm2S5X83NwQ
uEcAMF7fc6keL2VAp3fUZWQjpjQ+LAESIu7ZU4gjOXyQ133EbUfnY2CwpX0Nn1c58YBAR/JzuIwl
S7BiRUJ2aTNJY8gVz82aQ1UFNxgf/uMfnWWO/YKwasVqjezXkkO66MbjjbFwcz4DI/vh2VWaFjPN
kcKP/XPsr7xJz1p8uHJPjjp7Fwdp2jQUP/WHvfYByVtuFrCrY6DnEscyEHKtbna+Ss6tk9b8j9bU
AxNg+42f41UCBboQaXg2xuI9mGvqMVOjz+XwfeCRKQt8SYfauRUHmMjE+w4LvXWaosivbwxQNaJ+
ho4fYrkF+EtM+XVxQeXNER9HOnGXKEM8aeACShYt5+ajOqBxPuif4V0yELYt/goNE3tOE2tWrdLC
Y9W85cgXjHRs/wXpwww+cG7fUviu/F/7o6ly4c7PiPVq/i/OmMlE7j+Z/7W7bv7XGKJt0ddePdOV
YNtLz++aJES/eGy8h2Owt+Ft9WY0X42xZM2MNu422hrDFEHcCn6OAXvlRWm2POhDsCy0lPA3ttb2
PxAdPJ0rApSm9lT9Dq1kmO2DRspoUf3KigiCwfiT5VeIlYWbEJ8gyvJ6MEO75kaFg2B/HxV8SeK3
EgHl04BOPi8D6bMzCDkCEDDba61CqBvmm3x7IUo2bmRJpuCgYSGgzy6vPeTWSUSfbOroO2saoCL0
kKjk3RLBaQh4hpO7NFBAis46Hw/Nv/kMNY/cf4OpIb21E/Mb60a57WwvFde2mYrIjNEmUXkEqWEB
dCZvP0pfNfnAyQCen+2cJStItql+RjY0cYdWzKz0mPq7jK+2pF6jOMKj4T9YWjA5xYhusFJLKL9J
ztAMu0uBfP9Y8kCU8SY1xQN132QCSR2RoLBe3Dihqo9A3Z0l0nVy/piWPufgrenQDo3CIt37dI2w
cdU73lkRqbV+eLteBBhWRdvkMk3t02Qwt71d9FCmin2AxN404PrV8RBncsME6/TBk0G7eTwp+Jkf
QSKuR51MTaXRcuCb35q2z629/msMY+il8aMZItFFIoEn1VLolYUs5r1eM4b+4za6eNY5U2VSEzK1
/cRchq0mXjcDa0GV6jNsphatRIHv+zKQYoB8EJZlYuXjPdLK8o01x+sFRRC4WltTMQg4O0FAY0Mc
yDNs0KNzLV+mlMHJP9607sKO+AVNQb11Xyl5s7YSgfT5dI74MQAtrttUUuaxwd661CzYbbphIqkA
NBu6vbNeT0X+DjotuNi2QaEIzp+OJNYfno2Pdt49OyLLXQVM4g66fw2IKCjBx26kbTsRt5rUCX2A
Fhmt6pFC5LVzo/MhNWaDFwn4qrV7IXdLBlhPvdqSieEr905ZnZ/KdBmtDa+KdTNgvDna+Pb8cWP0
XS/8RW8SK8EknJ5MZeBQQxpB9CXzz+2adUwOdOFyiFwA7VFLzqMbfjLqt22fGt5uw51kwcsVAz01
47eJ0vijHzy+cSI0B8RQKyeG9H3aLJtAeWHIB/2g3blaJuUYE88i20PBM9B5b1OZ7kUQCGYuA3nC
pkDHd06yfM/etWEa7HLA6LnHyKlHnk34+p1BhtvzT7g6T9IXRXgqhP+HQvzCOELJeLkfGMWoYkjc
f/0UXyayliGbkv+sidqkFhypmUoUyCQKH8SQp9yGncOMFiai+Ondjs8aIPD0Il4iuwVShZOv9uFD
GGiiJwi8cBZ1czBtp15BJg5HvUaGLvn4/lFuttBGkByLLNn6+AneS5k6J5yblndJY7C3IuNRvRyI
pY4tC8jF8Lv+kzqgdTq9azJzdoz5OEvbJ3FYSt1KQHpDHPf4Ya2xUxFyeDEZOYCzP8QBioZFkkF4
AzgB4m5i+IGZTQfbdL7r/aLY7P1f/61QFFMYQWfRo+h0ghn4MrvYgGsrM/0OVrpjY2S8ry8R6TMH
BoplNTXyocsZmoZZINsH8o/T0Rk46wUuiIG6Nwc4ScXd1ZWOnjawjOF1/X/VF3HxnxGFmWE77SGk
53FFVns7OhhHiIUQBQXcNO/daxzBuNsaDcGjxlmKoR3cJg96LPj1de3oQPnj6r130K+GQAWnqwI8
07VZEC02fXveUyUNG5SLhL2nieYQJUvos2l6UcYUqhoU/dRrqGfHu7Zt/4QyWp2kBe86Kl+zLgbU
iK0vXwxp2C6vvoC/6ZHKS2MwQn9z6UTmK5K1BEIxmpbYd203fqGvwKPZVc41ZSncUyrAVAe3pmaQ
WWeklyfbb9QngzWAY2AuAwAh2BuHdyadag3cctp7U4XsIsH4CusbdIH4RNeWAKpHjX4VzPnRtoWK
ifNhT1UrNVB4/cLivzsO5oFWht5pnIQps2advHz78R9zxDpn4+MEa7PwGDT3aYPAta2YAeflLv2p
dVP0ZOxnydg0p0C/zYNp6B+H3flyZlDzQMehWLQ/mIZztVHujHYq1jK4zVx3kCbADkWrstiUdBYr
trPDZhyjSAvbqHFECBThUE1Bq92JEGDp8d1GYLyLm2TQ0dcAuRcwca+REGIRlvKWbCY4EyxureoT
LLStAvrZRatSOO7QmnCEgv9UEotU55THTDMOGwRdwXs30eQLZ0jPOqQiKfNz6uLS40qcwUo0jRce
abbLNK5UG5LCu1e+Bq4CWAg0spGu4YciJruSSRfWEis7NX018cqZOoNXiZWtYSDZD0FbHhWkwxHA
BABpBBUHNQGMqSd1nTUiC6T8elRljJhgnV0bxHUkf+VsZ6otgWpshpMIcGHXC/qlFFI+8qS9dLrE
UiV7nkI876K2GKHs+/fm6GPTKi5baM7S7HXgDD3zNfW2sbtTdJi58ZmRTlmbIAh59hYwdsX1T7ef
deQmYPuaOUvE3KrlbcAHT4993gMwc3mdY3ghYNf+G6mlWkFeqhOQclput/UjEPwVJVmKBNTaqCga
vq44nBbZ6aBo00eYGmP9h28kWXngi+zzgtmBpJ0ZoNrSXN3ZFZZxcKOXKGIhYloqoQKFNQdX4yT6
Hf9+MJ+3f9il0+mk4IVX7T70ceVm7qyZj0f/6LmxuKyuCRX5rubzSdK5rWF5TIsBqTj3Me7CBwIj
Cnn0alAwp/yAssScqP21EpVv0difcPgVGpADht0BJ1etkHW45Va81P8E+VnYCXzVM/msrH9NtLgF
u+Ki7cpXUJslShzk12t3KTEBPPisIXIB3+3tFiia4MBQTqXs4X6ah0aUqdsWVkg48Jj1t9OTUz57
1gGoTDX+FyZS1/JEzh2NXkq4ogwPyWbqSIzo4j7TYftJyvdMEByW0FnMv4Wlu+cPiM8g97zu33uS
r7uDRV1366VkWl9g9CBWw022+UBKUIZrh/YQyXpdypBeU/tbiYwWmE1gPwuM3pG5QQ1IZkyA0kXh
poWqIKVlJSrS/0lVH2FcR2rKANgyU1c3tHj5tAdvJwQgZUlE4qB4X+45WYT6b/ew0qgZ+11/oARr
cQutaTmmNWaz+MjZY3NMDOxK4L5lHfAbEzZnK3ElMROqT6wa6yYv7qzyy5FfBEU0KL1SUxM/Iuiv
ReZDgAjepH6owDYcSD0P1yvCcuurOAKG1IHs2UvovqjfHQUNP2lX/XUu4Tee92z05X44SpVcbcpW
g0PpBCXl7OtTTxg34JGvm14YvyANVTXW6TY2SoWfLJY071v0gEbjXZ9S/auoVnmQoZGSnI5F5R2G
j83Jht+LfXd/qowzbBMlrwlFYdhZyjBS3efrTrwBOdVgxFy2Q19d/fFYXKZr+DqzYRjFPEvg17l7
km0//Di+lNrQVvsKKv497161vQQrTk2Uh7WbyotBzoBFHbUqw5SkxnhSxWYXD1Fv8SpZYB+nh6Ce
Lc0nDOMKzVu5Jg+0EZkMT9vZYGQq83M8F2cHsnNalq/VAznp1dNs+otEpXyLV09DtSMiNNWbkXk3
voBJ/ja2OQbkRNuTxDOEVl6DTEHHdled9IvQrslGsDTDj6kf/vh1GXu6eYMlw0lD3JKIkB1H1EmP
9+UojkxuXvI0t56kYIXGcAIl4NwYnuxu2YJ8Dvou+VZ0Xe+nDFRfjyuZWmXjNqM2/V1sZaTQiK/Y
L2l1eC31wAJhJMwIlXEJBTYBNAOYK6dJ0aIRpTy5pqucSoonn7DWnXrwB6zzRKRmOMQUi1yfRu4I
e7BoqNmNYI22hYF+6iazuTKgmKTX05rjuE9BmktWrcsj6T37pBqa1vfMlF5bN9BarsubTactLXDj
uc/SVKr7OHpRqj2M/MZ2xDP+lqcURNN51+lmldRhuRteikb+HvQg8L3/El1A7Z/tsPNVc3olsO9W
RzvAykC6WQb+jUzId0ILwPTsw3Mq8G6tegXghgyLySGPMt+kb1SeT9ZT3+wbw4CemklHd8xajNQn
gei6baAhA6W8XiufswxkPLBjf3GQBQ+ig/SDZS42rw0b6Jv3HJiHb4k6SudZ7MIX1JfeE0FIYk64
xOvcBB7RLcMbqMqEhqqOAXJj4e4pKmSRTjRrXnHDCNz83ghfCeoRBsJqK8BDi9uFx+y+XcJReXZW
2Dx0z9peoScs46dUsEj/Dwd+ZW1tAdDEy9mNMZrheWWgaq2YE/6TsH3/ebIiIrB+znughPYi/Yt1
yA2g9P16sjWBw/3AFgP55Lcr5m2uLd4rHeZ+0EmCDWdcLO2SRUyp7FCzi3Gdi14WtAJec1FWkgI1
zCpDj16wBUIBiIrp5top4WSPqG6/ufZu4VdUzocomtVyL+2B1H+GTFZUiO52k/qsPjfkDpp3GRWA
DH14uMmzqCDhreBEzUt+UEf+m9WgOOxlCficefbVx/vm34IW0ZrsOWDV6pt7KcABkP6BCRdpFNyp
es1JGL/0VjMJhO+mC8q6+uj+wR2nr0Yz+o8PZsEfm92KjNcf5IvgJQiQmVBflXqUumZyx/IAWGsS
4XELCfLSVOhvvUNkFUI1nKZ24nLFjyYgvTez/jEKSR8BXyO3aXmpeQ47UOv8E1Q7hkamJXN86J9K
0+88x4TkoqNHX0CoX2XoF8/vcc36HUC1JjO0y/yCUr6PmSn9xn4Om1/LByy9Xtpa1t2mXDbg3R9c
yZ4DBNfaWT9iu36yLYokcStDdbZrEKadhZxHSBVUkRcA4HTzt2N3Jtm1UvcAgBGFw2rfQCRqOJ0f
tau7KIHPC6+QBUdU8dcj3On5O9P3UvXGBnz9Uu5JgN2kEkI+O1f87W+BrpCwH7a5Mu7l4TRPyQ/7
Xxiuf4Gbqsdt+Mnd237rwFtyCiA3Khwd6Xv5UtMGGeQaq9QPhuxJx7ayPWT1tVwYzgMbAXdsOHJd
hGinHCLejBDkqw4DHEt8PCLwum6cuJW4z3wNQ7gI/JwYUX986FuaE81mNWdeD5xe0Jsc/N2KoVKW
0YJFaBnpZ9jZzmM5PyZp5lP1CX4R08chstz3XoXYe4m3YiUeb08ZbC33KdSZi/oxNFHphO8CMqAi
L9UgSE0Vb+NNVxJfXgu622u0R02ECCIfWMdVwM0cM47ccifAbcRNlgFI2q81q5SmyZjueMc3T6wl
Ds4e0SoG90vn5wAdkuRMjGMo1PfZQfaH69pIwLWfzHe2d4fk6wedheeFo79vJdTOpL2O1CWsxTKh
yiZ7IIIw1OuQe4dH6CcA5UmIr/xFZP/BX0WRitaurayOqG7prP+Z9DoHwJaHD/tdhLflfQzpOZLb
Y2dkb9+C62BMI+yo9oj+Rws3VPvdHY6OQVDsY2t7QHDwT1Hh+I1Pn25/xlj1ZYyyFfWscewt0QmE
1fGBqIsU+In3Fh1kCc6VNtcFWRdv/Ihzea0CykNA5LaDqQo6+pyNDMN6BZ/HcD7salC+B5JtsFjR
fylkLKIHGL5YpKMOYx9IyVigO9WzYgAkZumw/J4xJrdZPUBdI2shihBMk5oulncs0duwrygjIkIx
daLs6lhrG6xcNc0egOkP1s0YPE4WAIZ8sj3OWJj1G3INDZdswvh+s0rJcHIfYSqa28eyaAI9LySH
GA46rU8xm0OkXrkDG2VtiByopIjUIxMYVN0d9AYtD2bg01R4QT5CJP0bSVgaIuG9BwHiqLQNqzVR
rmoQmqj2NDB9JQ+z+TsEE1AonNx6bs81H1S+IIIfFChkXwoE8W2vPER8TlIP68H3k466SSaYrJ2f
v2wgUGL6wpCLP1P68ifHmTpjOvncorC8jFwJngTrt8UTnn6kpVN6ZsrITV41AUAfiCgjsyHrqKbK
s3KsD96vw7R8g9q/Y+0FZFxWMqvd9EnB1bGjgiphnXV0W+ystxm1/DdFqLiXiWF9+j1N2HnbNwqD
82qSa3lKJvPWVraB0+ujSPwhRzORnLDOIvmxgfogmDnSCmsIroZNp9gHe6SX1sd2u32suYQLPgyv
F7ovQOHN7aAvFser1lX7XhiNYoSkcjWZuhe55LSI4UhRq+PQ/Hv8sxZ6zQ9ydp/FYFHMSkEC2rOz
D/Wu1lUkcP71TD6Hwg/IUCdgpz587WFDY9am7RWunCJC4J9Ya1ESYsE1jgvNMspDLjo3MhYz+Fm5
aF3axhRMP22trkn8mR5J8rpVuU/fdnF0jO1RQ1dqp4dN5gr7Hn2Yk4Ebk8WMXv08aH5yJUmg40q7
QX8S5oRMpbbOF+iBOdt3DV2nwS+kpMTXUV6N+cfJZgwG9bWmYAiCwfQ2cB07gEcdaSnHFS0Svut8
KSRV5W6vgjVlSqxMTzQ5UKqOKOAPM4REowaIyV0xZr1rRKh+eO8qeENBUxykwlakTAoMsjtCVJhO
wm9yzPIq2H52Hz0OArxNxVbjw0Zw/n74PVWleQFxyOWucuXKUh/dW9tXaFGc4lRaVrgoX+d8Gzmu
5mCNDxz0yD7CCH/DdGvM5zZZVIbsXzCYwT06Dh0JwsFa/WvkRriOJLCvIxkTXdUIgkrCcX4KvB2O
lngui3Ay8nFGk1jDPNdMCUhk5NATKbdgmJZhQzX+qxil85peFBL3K+PyGdltr6XzveJYRxjjdgM3
QtkGcrzDRiDOxJxbMiyozblFsoFGA0y83J7jzKBjxhdWGYllFTENmRw2exSCXYQs/yGxnzg8IVwh
OhmSm/B9IzkC7B3NtetTnpP/uh50cJR733VrCJn4EPvmqXkPw4tFKT9S41+z3BSXzkbGbydCIfRM
ChDLMRwoy3HC0exBe1BROGOeAe8WeyeBLJ02rWETh6BnBcGyrVBhhUp2xknheWdCWEkfpq6a8gN+
RH2faecrqZyPP+eeuLTdMRMhkVFRavX540Qzg4Q7YETBNRln3naeY5Z39mbR44Hd63xnwK/VM3sg
6JgPz5DGda/+7c+f0cuDxXlE89SqvniYghpaGodHqXMxdOt1nB9n1z40IGQb9Ls8L1be+ZpqHMsv
ujewpgVKrmKqc8WQBboXiB5EgACfTRkg1zJBJp88r7uDOQ58aqH5lyR67T1f5Ks1dghFGuCr/iwv
msxLMDTNKlXqbVhWgDEjjZTcq+i/DkBUpW/iCW+KVypFlrmvvPb9wqu+phMOQ8wnv4fNYqwKRslE
IHf/hanMmhsyOrn0yC/F+etbAPWjEphCeQZ9JQ1hPr/cyhoyOMDV0T/sVsZQnJZnTg1XOA7zYsxe
AJplYkI+5RNiEpSe8LFLMfS6c4sDcpPkL78B3ZgH7juKRD1i8yP1/+LgEIDHtmXWsCBAh8b8ioxh
gYf8wcqVa7rg9oE6I0hE3I2dCe9i4YZNl4OSf+LMISjY0eI2pAigzTloIrblEywqhgv7QYlhUx78
JPpwhTgxJoTTVCgdoc/w1Y2xVC27UQpZBfAs71UPJbwm0HdEoycaKyE6tZbcqZpj5uazKkwnHHKu
yfKK5ScaBSX3Q5jp7QY/pT5Ut0C9/YirNsuFzonRa3WqJxOji8n98zUoCI8Huv98OA6cbHTynQeA
mF+MBH9AWsJDU4o+z84y05WFCEgIZjY6S3bkqniV5RNg35aG9a6ZfnGxLpm39+sP1cOsjONb59eZ
ASReRhVXh3nDzmSmSnyhxGYT7QS42Gv5pvmSyxEsxmgyEE+YyT9793lvYjXHEwJPTWk83gAd4f5G
3E9FM2uN42JV/Qc565jhdqGl1i9UrwJbRwuGXkV7GU7tzoLKt2BvRUEQcYn/WnX9maAXlx8c9F2M
yE/KZqR7kBYPvAq9APZMEwQwQUMkGdCN4RaQ1sQIcaN8ahEuJLiDYNPad2SlsstDJ9odcMILaFDz
78QEKIG+0fT0DXp+ICANg2WEllOCVqUt2hef5R3vSfCaB4mxu5FPaPOkzF1rSOu3ZYZMRxHGymQf
fDBsFIS8AX41+iV5jhpPRrYWFDE8133RUHCwAjSe3fIdvv7Zo+exbNwwGA4DgDiAx90EqW4vwVjJ
HY+OnxVtFcampGthj9BEmViRYc59LT59MCSlN9jt+8pb5MDqABQmTxJSvphFAYVBaboay6JGe3ls
wWMskVlNBcyx/ydADxwbBthrEnhHqIZgqzn+D5eDgg58MLzsnopsBf9gAMVnyRFkK6RmQ+j11rDJ
4CCkBPzKC6hiNvgjdWR7UOjAO9BOsAJV52QloExRQ0aN6ftffM8dwZK0lxFeI/ypg7cXm2KktyJ3
v06M7sLwJ398tcwi3iEeQQtjNRRgNPb8/AAbhW/a0zrbLUkPlGmSJd6rSIPxUIMI8K+p9YheQdJ6
0Btb4mmV3zJIt2ignd8aWNYyGnzDEYi+xLPoZOA/NnzuyYCSE+Lj2k6at02LymSvZdfRtfN8rHMt
f9llOLT5WpapPnVE01MYkQDeBVQQGCe2OynIpwcmNVX30eBLh/3FoF2lQlrmetX5oBxj7Cr1+EAz
FKEWg79rUB1RSZVwb+0+/dfncA3W+fDkP4l3mjRldTK9x46iQCWExMrmiT29awekhApc3q5cayPb
zSY7WExXeAcMCqaxyHECG4DtjEZDfjMyS11uvZ6Pv53PtgYb5GAk12zTuaTV77gxhkLQzZ8Xmy/l
YfBPEW71h2qJjes4LCqjyLKHGwsJ5OSXOYsewoTX1M9rih5RZTQ1ltdkljFZwC1yG+wWzYw5RZkM
SON6nD5LIh41Izq5fgr0OcNWcLAaYdpljKiHI3rkWX3C7sQ1EqDIVVXpshpk5rK5Ya50K6Y2hpaF
pKvdD4wRzap8XkhZow9ljTvmGhVPueRdNN41DL9zq5pbpel9qETm1ZB6WJxU1b+H93KrZl1gF+13
mtxz4hGU/0wZtWeUPP43cwPCZmqtfQJmH8BQIbQTMh6pPASPtvGkZxIhHzmrxKNLZeVkzVmq0s/j
4KTtoBa2XIWNxNtS5Q0V0CuMd8l7BuePkG/sbfmcKsV9ayI77LYC+P1b8Y3lrQ3DsxeFuMGQXVLQ
d20ftDpH6ZRzediSdqEezTSOSJZ0YXPHXn9Glz5kgSQiL3VgpJcX8R41b1EyPle/bA01Q/bkjPGK
arJVfFlutHS+XtsdC+MqVwKmfGn5xMmgXVVeg8a9EgnpujotA51PV0z9ZGsdEuYUG55VbNnvb0hq
QqcPnu6US5wBj9KeZBTuL5/WTK8VxjGGWddwBkrruJYpywS8WspGD6aFUVw+aC+JLtDaqArddgm2
99Flgwilmpy2iblEPrHEoe5SVpUaFizrR6c5iaOtwJet5Q0rev9upG80R/7Vj9K6BLcJMSCdKa48
N2YSXSU30IR/cH29KGoUZrqixB0AWramn1aXd6omgsVZAL4vh/oIlMUErzPXBP6zzotWaMU2fl1u
RcGgwSK1w25u3F9tHuaoYTuLUFps9K39ym0VZ4s8X6/qD063xmr9gqxuFJ1GJ4CIq3Oy9MhSm8o2
kwXch29s/17uZWMZnhvCbfAKM8Cr3TR3oBQYMCs8kos5rTyW9Ovsqw6ImJLqrVO0pB6qYKEvHXeo
L7X5Q1h6lM09YvmGIijpw/aHmTFCVyaBRaUpzNE/Ex3i+NN0sBzOqay5Cn1LsQIl4A6BwWKqhE3w
TO/1O3FHqjJ6yY5SZJge5USsCs5IeZxcDT8gDn8axPp/s99jaC0V32ZszpE7rZGMmRbdC8535TxX
137c+oxv9sajchA+EZt1Sa5/NkXu2jUndSrLPAmhlyaEcKA++eapsBW3jTS+t4fmAtTHHhlvIV/Y
9jFv59OaUPBFS5j5Z4lUCSS+RFVOjJxi2nNWlBA89fKnOi9hTCCEbZlM89Ywid7bS+bezTn2mT++
hJZy1ndsrPfj1Ed/Fy2RjflflPSZKoYndtb8wos0nXTjr9rKwqxentLBOUr2IDKrybvIXxA1zWTO
FI64FrnIVeUrHNHPrED0QRsWXVLyDXdrORQUwCrV/usQED+9NYlHOsbtpT/yLs6RgwQym4sF7HCt
H3PL8+t8K1wpAGMxhseONRGCyLjTT6OAgx9UDd5+hLMs42FT626IqMXbUzAk/omG3Ns7OqCsOrEN
tjTMnUlS2dCHgRdso3MQ9Lc40XTuUrQJspo6ssCeU+K0f5FwmxeCI7ngU8RYgc1rvpTskia1ZuNJ
0QGpB/MbJ9gzTgUAXdxr7Td/+rfJjlv/B4/ttm/TYJRbURlhPQIQRcuDq4PfyO0v6Ugv+1GIXmgG
Om8BRa8mn9sZ72GhqxUn4HE/jl4FyQxTVLLGHJVeVkEPgUwkygHK/5QUSGsfFMYTqQn2NK81N28R
3jbt0d85A6o2F8fE/TJ/uA9+fE4ivZtegs0Xqdh2v+HFM2Bir+sqTxJWYUTgq6B2+5pay0L3JocY
fu1Ktxi5n4pVIbY5ceeV9AaNLYjKc/cMNZMf9TJDepBrZVVWPBqZfGlLE0/7IHaorGfyp5gc0l+V
iYRyyHgP5MWO/aFAWZa49s0Nu5Uip3MvER54PnS1dzVNNcG8J3bIhP1WoGDFpc/UuxU4ZjT1lO2C
X66XmZ0EyRMGJEEOM2QTVZ5O9X4rZu6P5sZG/OIKWyhApUsNHfTnEahQD/TDMAMdW1680CeGt1ez
X7WEestrT2VNlH+V5LW5CPePqywmajA1C0Uc8iGqnyOcImCEnsMLCB3QoAzInRiGpvonZJa3J88m
Nd0swQOb40SnOkNy/Ehjh5L7aSO03m7KR8aNDkbKmXiIhNCns8eWslCqx5AAhexzlSKt6vLGx76D
Sdygs+zELAdShfRiAB/Gb8mnZCsq/ribVemzCcclxXUHdQ0uZs3K82zFMvjHz6fBIP30BOyPwlvt
Bjim1pajVJ7moAylnfvIPSYh6lioggMSTgvwI94OU+0A0ZJl1yGB1atOgFCe4CFk0wZYNoSH24bk
O7A+5Mjm1Qc+5PuHcYBt3RLg4fRMzQK4apFRxiEhgDkmDBVSmAKLjES00FfVJfZ6Ax/WJmOXLNZg
G+9mLMQYy+aFH4qbwoW2cqHdLonLccL5dm9oKYAaweCIyI8g093shx4kdh6WH1TRKAlHAt5n9zY1
YLXTZ9J0p0tJvEW3tLOo5loVxZY4L9GEWjAHiSUjBS/chbv/sG6SnEG9pq2JSZ1PeAKHw1139mIq
jXGIaJVS5kwu1MyBaYWM9ljXeactFPIsEq/iWxWb5k8skLQo4vDLS+s2mxPg8O9eLzWQwllSiB6X
GaSnNDOHxKLdALyvJ8T5kr8QUKJdayCz+sAlT//U3FZRCyXBGQvmP9FWDrradRzSf4Lpgty/82Ic
OHROcIIUZ+Q1DX2jVDNtzSB8QQIJmZUU6deK8DpJ6xAwzAzfaUeFq0CXs7Axo3LmChb2fT5Zlo8G
9HVG7dS4BW+Ay1NgTgI4SmYM01DA5OJ+XuW/MeBXSgedIU1CU9HT57k+Wfh0QeZehZwHu4tQidVs
vk4CaWdRLNpKZg/7va8z9urX4OIGi7s9LBXEzB0GAc/tcUHG6uSmQphSi4iRq66ae6kS9nh76BBb
6I66lDmUIMUwviOQ6Tq65n78S+BpMrbZfyY5gJXefg5zvtr7AUiWy5uaKD02D6JYtbg9QyN81W/S
JDmEq0KRqIR83cKnjdquoFP/7XgIoBti6wwVUTkMnAXy1W+zaz9XpZKKTqjA8tTptxPY4GqwiA+R
lfdIm71IsoliR/OkUE1KDVZPM6BT7zlS+KoiEzFk0tChTzPgfElKKyZUsWrIsHa98Nfz2Op2m97G
BUPHax2P4f8xIk3t3kMzm+3lqdzzsEQwBhEOz/gVRaUjOFPx3vVt6dyQtt6K/RCg5JDZFzjoNoKe
CPJgFWeA8SnDrYt3y6POTxFtyfBWYFrjtX+9gjxN1u6mmJ4m1WyUBehd03tJV0vMC0DCZ8poLxpE
r7vsvT26nhw+22TNzeAnDUyba8o0245Nql+jQK1M7frhupBebpq5b3qyD6dawSafzRRFarJ0YU/s
zsMRn+q5a2feNIDs3H9mJNdXM3Zqh/IBRiBv+hccsBWaoFXUmaHZyXRrdqyg+WuYatF+UEnAd5Ja
8R/3VSYreS5TZmsW0GjrIdF291myihU8NTkxh0e8wZwxapgy2jPnnAJ1+djkIjO+DVS5ONdBZXXg
ZFe0TJhUEes6JWxi/vq2T4SVp3BWZFPpd2H/2tiVdmFgeB5iaKq/vo8zNTqT8X5CS97Rlv3qZxcJ
ZhtJ1/qfehks2pRIwmoHkbFq64qmUp1H9sDOcYKsj+xsARfJNlvuUvwE3W0i2wUTT/dNbPN+QVJO
5csQMmOeBsMAC8LATcP2wS6KKbgQSkqO5WrBdm0NhV5GAqTLJ49nQG8fWUONkpYCjI6G+ZGGjwGL
yTRrHashlFfUsey0crQ/nJxsEejjUCG8e/yimdynYoeQ3TZkLwb7Z4dWfnLY7gRaRMSor48ubixF
s+YgEBdwns/enP2pCUMNjRcS1NQ5hfBqTcWV6ONpA+YQ257CWr5VrqRiFNAWy8vp1fyD54hItIjz
GAzsiAp+fCQwCmT7gZ8GA1w/vmmHHjnHEdos3R7HQs35JtVYz9OdTp98wfymGYu7FvVTOCHgfTI1
32KnM4yzro7+o2AvGNBA/hXguXzB3beGHMLhSLIUZV67Zp9ipgWw9YfE2LL2bin9qQ1xxQ/Kf0bf
QO8GUi/vIpABQxAdrNQR05xZgurB1pGvLa6WYEnKKvCgiJHqlR/7iBjvJfcv0D9Qwhws8Hxbwjui
hTNLZiK96UZeqGzKCcybGJbPMXc07C1n+mG2gNX+J1dPRI48KXWzeUPn10qDjtT6FjdSeQU5JLal
orgmsGOx5XXIbiDQXd07U37d3furE503bvAma7haV2j5pjlFDHRF3OsPTgKaHDs300o0vP7y9+JZ
UqbRu+yR6M5uDZAALaxm9spPd5k/k9Yy3U68gLHFRqwViztuNgUx++eagDhneL26hsFM4W7QVkSH
jp2j9R1pfLkUtFxU+0ZSTKR4+U/2g1z1pyXPNbJ97kKW+a+SlIDuoikBujzuYMki00IHXaSlLP7+
UMyPIVhjuQYt38bQpukdhXcabqTtiNRybPNRBlvkda+JMMTRGRMGJvvQE+FwRxNNJiyAAQzsS2Oc
TJ1fUHqQxT4fLiMq+sh4gn4G5U2iStzHan629sbgIMkyjLj+zcyGZKuA/Q/M/QkUgnTCghB7ZIzw
3iCJ/HxQgjJlJhdOdBEFaGqipkmUToDf6agRrcwcTtn7VzD7wfXPDQ/2O1QB08qXHfQTRbZxq4ID
SmJr2DPfYIlPHlRE89bcu+8DCBq28COiK7S7sQxgBsCZYwSwUhkUBPVyuK4IfBMGOuiZIIquKeRh
1WS0e5OjytY+bguG4dACYJYa4Sq2Zos0Pbt3wGyB1m16gGzADtBMV2uT3+K4a9LNwS3Hs5+tmtzD
QoPiH4cW5K4jPcc5sQYHu6rYUUjTfjAjv+R9Miwca7Cstr9bQ1RrBAgFFRNYZBUl17BSNF3Tee8J
babyVd20wPav3TCvswBVYfER5fd55Ia6evCnLg2/hB+2CodmmHf7ibAEQyFKZP0sF2V8CkSKSC/l
/SBhOjnsMfAPAmWk6FlWkcJk8Z8JDNb+feGsrP76RBRH8bvbxpKZrjVTBhBEc3S8TNAyiQ7TJ+fq
LySspmw9zJAyfrzgUorq0uhleFjs7SHj3231WtrlNobEsB7+P7h1miqymz+BI77wDpcThN1oHoTi
OGbKafEBF8Af/8d7lc8e3MT6icmv2pBLjuML0oVlh/kywagbEZKqR9blg215lz9GMYGkei85OscW
SjUikTawVdajXTh3sFemAadKHL1ph5pFW9VyVrrZZShOnjFrugNfke1jJ9UvwL3dEbW8gtqt+hu9
xQ1BJJoHTbvT02xr1qdh85SKObzf4Dk/oSRomQjNZ0L0fnPY/2UZxWYr7lnmMsZdEQ9k5VShDRlT
Xswr7xV/p7PC9h4/gEZGelDUO2tbZaH/+j0JBfAzyXvKAN3eDr9nB/LmTRDdHqQ9t1JEeoxy5o3f
vOs2PRpNohR7H7UokyvBiMZlPCdGwXaq3O0DHf2JpwSv5J4XMzMvbw0bbkXB8D/l7fnF3N080F2V
tNWqEQxIWnLXZc12gVU8YuieD3E0z3ZBAPMDmA4O+vvUZgYzo9tn0LwueomORSOxboc5UuTsg9mA
jgVQRs/pyLdwhBeevM4O7ea5EaoTw+J2PaqdcfscNEIN8HmT6Yx2gjtDGzJKdI7MhGbNi4xpgYyO
lgv1/GxSiTKDicdv6Jpm4AilyJacA3IpmboLnS17fgC+l3nvqTM/Nq4jwE93yitc785a45etj88f
yQKj+nuIkGNu6nTtoEc3YR59j1GC7GqCba5sBIMvxZ07IdAZWipzDvttW9NvrfxuOI2Otvbu1WvI
sST5OgzQlQYqPnzeRSuY4Yzyi9Lz0i1KGYfQ7BEhAE5b8wWPv6tpM3muSSJ7lTExEHl7aIrwVxUA
OJGi+il0+G8aoXRe+mM85DyND+dMf+KGtzaqwv2l2VMJY/xTJMpeyZVrps3QGyCBDakvTueyn/xC
qJvdRH/A0/4Xe4626BnJVGdh5WTexB/iFux+dIoXzCVMbQttjKbXgC4ofjh63ytesp5SEpmgA7tn
keSGa6l/TiiHGfiKzcMnZH8JeYl9d+qSr4PvsreNO970jREOuwOKe4ueE5EIzWE91c7RWDX0SSvA
S06wOOuu+Jloqdgx22l43zVwcrRDf3pb4Bi8Y6E60//ReTVEA9pxy8M36NXMO1r7FIktcirGHAz/
sVGwmqXiJu9nRsP1SU4wtb11aukO47XwGw5alKv+xbJ0aFizZiBCgERZNZR2ucgwKqaLpYHbOoWZ
YeD5JPxqvUMUBmU+hu3mNh2gtGdGqBFVps5azzsVCS8RzGO/BIFM5uA5JCjaTlaar0iXIPhniMOy
bm3c71NqBHA0gxbPw2b99mREcoAoD/JTpQ1l3twPCMUmKCX9saztPgmjX6ImlCOqVVBKdveD0uuV
aPnXpG0ZGjmfVfEVfC4C+V9R24ehil4aGBhbUhZs0Rot8jNLaGoVUSoYXcGzhTVLF/nWe+agRiEb
xrsfWDH5UyD35yKrLM7+GWp7ZZLThYM6hUJwbLqIjaARscycpKQyHRDm5TXqAEDR52aMbdvrD2ac
x6D7Y3Pf8rmOz5pskZLAWgMtdl21XhWmrKyHwoOrhzIvTk/DClShOrp6E/4fWEt6L7iFvjaBme9b
/n39EDqOScxTxDwtlLzUJ1kPvnvNssNS2MZMEoo+9ZLr6iIKrIHcZoc6Vinsu9JdbwvznI1vzuEL
/1ADzcrDiL9iZZw+nGUFUXBbGytMgJpxkmcOEp24Knc6zELbKOE4tsJz0+6Iym5mqDmNc9bg1DOU
qCwLFwKfCWHRVavW7c1Bp8YFpQ19ZyAfEoy+80Bp6V+GEYmVVGPh1GLA4yATkB6DJpC+prPTtd4F
mNarQnHLgCob6ZK5GCSCQc9Xdbgr0wA1sLd6bS7cbn39ly4Ckl2qSMw63XbkJUcDDaoRjIF78+2V
8bjQkQjnt9abm2y6iuZdc1TfSzwvagNPLYkAZ7f0gNvUhXzbrJb2uQAc1fVQ0xIxpAy6xOrGvuNA
Kr1Iv4GDznGK5AxIi879Sj1LhQBZlyfPQ2wfXHyjFD5X+3f2Ji9U+S+ycVhNcHxaPjQl2eko5mK3
A4nnmtLgEKP5RdZ5DunzRlQFQ7Ql7L+bohYqmRaoq325mtphISHF2Y+Y+aYmxu+FEQYPMZHS8U5i
LX2Cl52rJzZRmvBCbf15lDP3Ltx/4lusFAZUR57dyMnYbDpPywUeJXUysy/mES7RiTe/pj/O1E5g
TW7ZxUf5mFQpj4nEWyF9BK7ZrCfODcXy2+P55kPjo5sF0U/SBSoibowCCo5ROHQW+rMzxZ7kQCpV
FCXNXF9SbEpi2p99fO7UMuVr4OTFk0tjOHZUDVHfB3RdV3stwLFFGa7ZV9pq1T+0Js2Ni6COK/tm
phOwYv0o67DDPlg53xOOyWzsQ6S0LIvVP8IjGKacinPcHsweqR+FfL90DEsoGVpHpegKwN+1bmQU
3zSYoIWky65FPirqmuhJhTLCqZMlNC8G6cYo0hVYVH3mH0C75UCLXX/GpiRFbZSHOBXUZ9wd+eES
XYHnCgHeOidl8a3bMhqQzX00MeHqBYRI1z0jo6sRcwo9/WdZdlBywf6hA3pmQTLkK1xDyrJXqCat
Y0gEOZPv65pKcvel7iGhv3In8XSMYu/zw2pokzwsjCbgP4vvZJ71YKBZibIWbcAOLOBwDrjDO/9R
FEaTNN0iUYizGz+LG8OnES3y3DnDRdYys9Zt6LElhnFvSNSAk3BEqRstm1/UkRME6gUbY3jeh1hF
/jeZtgJ/C6QwHXhX1rbXNUuQjDARFuwJOJdy/a1orU/R7akufuBqzhvyUJN35GO5ROtc6yeAKZxi
EOFvHA/j9lrTfwPIkEog0pc5yvOhTFWcTxgJWgfLfOqsIZSFrL5iw+tUrxvv6Q/YnVs5UMa0T3PL
wPJp+tGmxNVLTGIGBYgO1OjW39b4PCCE3RcHyaVeU1q5k02UDracUnNFtcJg9YkKwnTawZFE23lm
Pf1jheZJaB0Iu8U34k4rtRJ/PCml3z3hIfKt1IW3tuLhibWQBTZ+ApsIE/Q2xkaSIwjLCeiqPWrn
W6DNe7p3ky6w7KJIQzHd/QyncbLm4AIv+C159TBVsZOWtryAhi0afL1+FBioTf5Et46dMAncwouJ
FTHxtwNZIdwT6SBVNpZTL7AYx2XQqjvRB+WemTVniWiwzdLRAxZ/3Qvs1N2K15jRSHgx2LH2pEL4
h9QCNSwdwVrCnmBk2RrY4m9qTpYvjeNF9d1/CeuztfVB/IIEvZNoaFcr2pv+p9BH/PmqhZptru52
bJv0rWnfK1TcHS7rEbopzhTwvxBO42PDKbASaKXF4znxpw9ZwoqajszL/sKuF71s6yCz5gmB1/2/
0rBNhcVBC2k4wQqoOL4kYH+RPqcR7VhcZ7FezBeSCkVeGUvnIQ1Am3r5S1ZhNHf9FdjcCv7Ah2rQ
dzki1sLH7DrEc0tCWOpSbFq4EyYM0zHss4eLVQvctL8jDQmXH2OJtnOQkJSZILUbUQ8FkMRTMl7+
zH1fzueu7/vTte1gel4icmP4+Y1RnN8k+vxvjeWjIjD7F1hITBVzJDKDCHfrKpYVOwPmtBK9RWa1
lmdMrmLY7Nrzc2cTi+vFjfeKM7ssi/qQ4Y7b3qGQcxKXE3CvA8JYB9hmKY8cawShZclcIxOaj7qC
+4VYfDWpadRiPUIrChL1n01Q7b/3jMni8EO9ZlXWwe20W/iG/Q7jaw09/476fTFGCHsCGhn7H92B
lmO8peZfuxJr8OwEaG05ZN5SiUgP+F4nneEY+efmx68GwIr8ZQAjdqX8F5yYNJZKuPIin4tjUp21
AbdU0kM5lvoRoBE638gbSbERPvM75XmJROgzTCVK9yVefh2KdPYSgaghg+mirHHCkAHMB88/g7K0
gYWfaLipBKh7WtqInpxeAR/MMEvH+DmCZZcPn0VsAB7I+nzy0taaccG7kaEgiTqN/qfG8aPkGh4W
huIZOQM4JWBHVolUh8wiySGYIYNwhv4HtQazyvjNZJXUhsKmkygmh7pEnRI8h8Ukeou5KHANZYmH
l9jOMQUDc4nzC82U5CXSVE7z4MdoT27MJdVJ1XZvvyFuz1+SA6S8CLzwSuWM1WuobioVDxYonVm0
RL5cGQQ02SzMJuz9aonV7wEFg4BaUgeSbenoj5STvp58jQ5Pl7LuvDHI34kxaJgy2jHXqFQAROxa
VO+yNUfTdtNXgw/fSwOsNet14hsEptFhlwLulb8xeQ/LP/5LfBgn6DbPuIsxCT708xvXeop4qgDO
8ARh2C/1XuXI17yj6klCXHm9S6zuM5RKS9qfrY0Lt0xKwKJNnOc+zKkf/YE62QhCKyPVVA6a1gq9
KC3S7PrEcmRzqMdyKn8gamd08pE9BD6jNDBfULeQCpScKXHd3wyaaOh4/rrOmPt6MM71ovkLRlN+
bQSKF47hUYkmHZvisjVG7Yj0XSBHK64Ni9sr0wDBjP6lQQ8gHP3icKbpw+NN5yVAMv3rOY/kwvvu
hGUY1s7Ivx1kzQhdIx8KwQkUevSwq1RYCM3T3u5R0ou96a7fX2unCUuod1muPTE2pBIn3/hmgCIE
CYDMZh3oPJNX7DvCGCoqCWJHzcvR4eSD+Fx+xPumCRTn7cZZeiENQYy1kwqaF3YMekTeqMfLrMXM
E0hP5ZJNWUYh1MntdpIRcRGn2xA/CsCiz6Me3K1Txl9/btarOzQXixoh7ZTnQ6pdJ/6hmJCQEOGM
BJYpw+mUqtNJOaE9g4KOzihfyRfzRZBonHyt7VfuSbfE598fChJCrEYq7N6+5Ff7XbSXoYZW1bVt
xUIDrsdO+YvZIvbV9iaOzKqoM5D3VGIb/H18MzQ+bsQuevarVYvpwqCVTEF/6aVaJzH/PRrZ4cbG
hdsTsL+ZaFMF3O7w4i+Rceh9odU2xj5fdsIjGcKCjXadRTtXobR1wQhi7RCzADjsxpDrk8nEsxIo
KCeA0UWxV6YK+Jwt06c8HSIBQskLv+MBw3YS4C0P3HFlx2W0HlJLvbT/cC/ai/R3e3MN1+/mRrB1
s14TiBFk8x2YALkrjPLJ+2t9Qizegwd73BrbuakvOgqMKFA3hFapAuoFeJA2DwDsqZgoNGy2uUhz
CAAbPWiy5YcyGFzC4050SxfGjskNdwocE6XVQkki0lgM7kCTk8inz1S6/pGaREx4uxKc/KSnGSXC
V+SajSeP20PSD9YjImGS8yfP0OBcbRpkWzb08AzydhAzPvFdTS2To1wWY1XanJpiy4VC3g80Mx8/
W0vI1UdTtVwTytmS6QlWmkPKMBAAKUxQTriGb9cG1uKYwAQnJ0X6lDZiyvR30aNOrovWy1zFhhiJ
Z1y/RAfsnbHE9r7p8xV0XzfcsJxGH1lWUCUeRv5NJ74Kn2yqPGOQ1B25qULVDOIqti3zvOFj5cWd
eKtmExPZhUTw+RbLCHJgzLqoGGtodZukaQWjEnR7P+p6IfhAGEOx94KehQ8Rlla44GzTvgOzCR9L
A86Y+FmI+yOC6axrbfkpSSffVqwxYUMjUqd1SsBWfNRA78DNCyGWqxgzcVdDAeeMh4swPetew9Ai
0RxQHT/s0AofuMZWbirdrWP7xkB9a0C1+SKy6XWUEvU52yOyq4GLo1s/PAGx9CVA1/todDFJNSDY
/Na2K1SxWxq5PRQP36qkgP0Woy8eSBitAj17C3svRCUlvqnsJoTC/vFae234mPLWoc05B6Ygbcqk
S18M/jDoAdUJXfmTZEKy2DRHtupiA63xR4vzXNaLlNUVpVBL+T2WVAdt0HawsmcSKsaGCuSpNsSh
fa/hdC8hhbde/hz9j1KSKD9o9d6VLiqo2LeeDF1jrOFmokJq5/9+P8KlyxJXOkaphhK5XbmK9i6I
aGX2lzDsYPjtnNguDWKTDSjIZthenHnaENCE1jgkk1Ojw/f8nELu6AdXXME38hXjRJkMJmytxfVc
0bf/8VPSgje4OjMFSGdRYmgw1tt6URZGqQBidCXE3PaEpvAZ4sI2/7VFwlqrsXXG4Sik0blYyPnU
Xkb0jsAZHQYzBepEF3pyfowu9g6ByFQg1Hwjn9tMcToBJNd+DxCDd34arOf+iOnCVqyzjuxbB/E3
TMTy87Plf3ZP1l+Oy/G9s31KQPf+XYsfB3lYHWIUfSmQqTqHS6yCVoYqC1I7HqCLHKhHPhVxxOF3
xxhsC6VXVH7I4Yl967MmTRQqMvzS/WChFJqtqVlNnVkYclvxWvRX9ZMy9y/YXaYp3/uyFvudcV2G
1RwfZYMwx5AsHzw1s7AIQQbQGfJ8BRNb8TBd1MqfAKqgxdEgU8HVODUvlge67SwjHNJQurKjHnET
9EgauYfD8hXmPfOGg4w9C0t0/bP00/WxeIBjah6et2wJU14kT6bJWKNIPbpnyZBzxgAkE+yT1CDP
byCp7ULrHNnKCybs/I8fKTKnJwNHs0Lh0XY99hIrcpMjr46/GLB2j+R682vnJqL5Ikc4FU3ClT14
x0rgRdITaQI3KyEA0vzf4ihpNBr4Ma7zNEqgMQnoKaepGMhvuWF7WmkVYilUG3nQDJ+5cHesvkNh
k3v83wjCHr+Yw2GpWGblumbNK6Q8s7ynLCnRo1NskXMvNsVLsepLHUplRoRLmZ4q0p7LUrLKozxv
wbwcaNYreZ6qw3pGwYJ81CgjCMWgMJ+q+6b0nmpQxYdO94ACBT8eoQI6SViEmHZ0qdQwzHxYStSQ
v3kPNW4GrIfi4nBYaT4MQgWuY0BNTbQ1z/iZCcYqzRUyXQBml7bJ62oMEmGTNfGWM8Y229jmGjGG
TyQQoQz9L6xjnCiKdbY7/KkE8P73/pJwrTOIH2rR+yEqJY5Q74SBUkvfOskjWChhZjPl/hlC/E4T
0xXD38MWGKjoAiYVk4pRaz752aE69LamUpEZjqWojVJo0pVOOoTs8et4tKgPbzdgpk4Bh0OarE9T
BCDxRTay8jDKaMsBQd9zutCa0GrPbAOlgvj8QMX4/vx2aI4y0VKSK7H5vEL4Trv/tTxiEcwpcACu
X1jsZbuiB6Vl0JUIxOeyFaP/LkOz/Z3uA+EwIJg6QHcZhc1SvS3xS0NEg/LKCp0D/pdryABnhne+
sGtz4hfVJoi8uy0RR2nV/kMCOzlwz+47wWWZJ2MWyDu4c4bo+Yb67XCdDIMPaX1JolV0HEp8pSxH
m6U3NJQxpfE1tJTWXx+j3rBEq4UlR8b+72VGaCG+HUl1yO4kZs2QnT1pNZOX3YXhUiQbd4RNebIf
qSRzKtMXOvrFDynOqt4Irp0Xk4R0z7YbdDoT6+X8IyyO3DsOGW98nyGRhQIjvvIf67a/kJ0dtyQ7
yX5Bpumr1YUw28YBi+sibxAyYTJjOhMjaJ8uoyFkM/iO2e63xchnQ1D0x8UBTp9T5VIGtzGHfQfY
VajFtm+ItYPXlSuqK5VOYIeUbPp0kB6Hnbg3JyWuHJRxIkK7kl5m6c4d5hw7L1vMnsDE4a7WxyEy
GOo9Gd8e029si4H1pMoE3k2XxVxhu6M8TpPa1Fo56z3aeWcbfsY/gYmOVn5srarTvIlQTdw7vYAt
Q4bGKYhgPmMiiMM8/jwyu6XvegjnEpSLDXK9glEXdDrmy5VVHWiwoKTXtEC+IjfEZPuCePEtsW/q
AiFseTTZK6lopzHntP7iovEUZod5+XZE9Vo3U+gCQucYQHQUfRWQJPQz8PfnkZbJxQKtm6eHiahE
y+3vOIaBwzffFsMJHeLR+jqt/XmRBLWODdUbySNgs65IoDEsOSkAfI3wTRsYFSe0/w2ozAVjgS9J
zHe9jZqCjgN+303rU9IIWLdGB1gfJV/WGKYmsX/Wxu6RJtGXTqkdnAGITM7IRBcuXkbwIVF4W04j
YGlOVfALS79gcG4AQcrhyrleLjO5E5ysRflhWlPppyIYtkVr+2qNRWx8BY6390N4xpyPUarWiXI8
twiTr+KWyQkRjk11n0pW+N5mO22350CsCHP65r871lC1QcpuNzlFNcAj7oMSGLlo5xYnpVr/X5wz
fsTBOOXyR7YmA2+jTgqLSGBmXYALVk+43K9yKl9l++SPX1fL0/GrTgQ1vpfG+V1CDJpgssI4ZREp
oj8daL3oYbdDOwl5/3xk1ygC3WLcywa5eaO9HZvsd3NlplDdup281UDGI7xCygvvYOFKiudFM1f0
fEwuO3WL1lNx8PGXgznSB67XaOstt3Yn0Yx/DDE3+vgpnVNMc0/vsmbvOntHRXYM5VJ4MNggzD6q
envVcoZ4Ib6i2yoADj4Pj0H8E5kupS/EOglje/A5bUPW/3YfdE0TIrjJOjcJbzJrSMJLJKiZCV1q
WvPcFTHWssSkvIjWdA7nBVOYPGYdLQe2x2jRDyks/hU1eEXH/Lp4/lyKhGjKC1R6y9x+9IWdg44I
nGSEDPX8moHScZS1j4a/f/o+i+9UGowsoh7agWT7ToSECpHxdhJPgYN0LB0BRwl9Qcey71VZ0l2P
3p2ORJ4TkfuPE7ar3keLaLlvzPm7Na3yRGeOBFlAQ+gleDHImOajB3+HvfSicNnCVdsdrDO4r+mL
wgfU2SZsp53n/KqPSgwlAu7esiwt0b6JLWW9+kPBxviW7kBjvXZrRunli/OBraHkaDtQVg3GOC+o
tRK3sagPwpIvkfYXqRFIouDXjV8SQre1JhZJpRZObmzbMu/RJlO9xLxg9+mAqGHEz9jHHRTELtEg
Vxm7Vgs2dYf+VW7Y2LW4cszs9moi5FdjOop6k3tT74wuVl+11WFyVbW5qbuGoEYNwH1nx7Zoac41
wve1XcItPUdOd5OpZN7GUlsI3h4mgLfZGbAVTWMZyBrSXCYKe1O9YP+C4hWoFzI/gRsvWbBaAJp9
qBm71x8mfr2kohUkOZ7XtkVr+QSvRlb4Rm+pTivbaA1EpZyt5Pe79nwdjhUXjsw28Vsut0GVEyMl
90v4y5ibnouf2aiYnY9E6hti3tnmK26CRLAL6VD8Ajb3bhp2M7yZvfMr5Qi9GQlwUXKGlCmTut/W
G5Mo2bgNAVZ89d0VgtiZPq/OrmnTtmm5xNblIljuNwECsBM34268jwnQfjp8q3PS0+xPeG8BajbA
SbA5jh66GKN2U4KxnWWBLY0vJEjRYQd0r0FE40w/gv6+kQr+vxv516LGFkT8JWAw7aOpLyIjbNTd
Hf1OAxSi+bWN7X/rSd+acka1bzapHXnLNX1f5q/EEDqwfdkRXMBxZJhOYnQmSHaZhpnOOIj9N7MJ
PuFiKMriF/Y34DMjE0YJqu9qhQ1BETlswZftTbhT+8ZZ3QVQLHAFj+w2EnQGJo/QuI+yJgmMYMsI
ZgT+hrzSHRiaOvsqTULKQGFIK0aQ14CAKQolWecVv3pan/hBtSLx2ci19nagLKpZsVPmndSvZc//
CClpyAfWZoiLe8iaqr1V5p5E4Wb0N/3Gq/fYVOwuMZrhjHgRoFuk9Bsfb6k3txp+JBJU++LOwctJ
R64PzTGWEuT0PTi7yBud2QtZ5LRixfzblumIIx2V6EYI51n70OKXOGt4jgPGgdWhapNo4nII6IDB
6GVnM/hTMDFZZIwjWdP2TqmOPCmF31urz8Fr/JKqshlHCDNKLVlj3FjhBXSBnYXNBtYsKSXzxxnl
sdueB8cslbXNrTe+j3aQDnTZ0Bx3HMt1EHWXNZF2zNamhgUbtIpqFODlOm/u7JxG4g3KQn40OAYh
wRG2Hrs7qbhZ/r0/C9AD7rgwlIEzjy4cj6lVezwVfpZxCXckAJHoQl0mhsYfO78gGJXtiivUztdF
zRgrc8ld1f4pShmKpXy0Tvgke7OuHydE801Pb1ZuilzeZV8ZWO8fnAkaEBbBlie343P7owrmfru/
Jr4IbR9PKXHcU0gEfauSVmf2ZDoJhwSTXaXW00MR6BjjKCGydSjvfvq2+10y134HMzgMLqJZgq7G
bsdavtjEmobMlYfq42Acv4u+D8+Qy2N32oykxmNmfAN+hcRMzYveJ6JNaSdnh+NYXg1fHYjUyf3R
kfwRWWQRa2jKbx25vtHamB+1kN5bnAefwEd5YodfI0vffpWFsb5uF0aZoIqvCBfyFax7NNIzZ9Ba
3S1aJobTU0fzlQlPIMiCUE+tp+/q9y9Mp+Sz9tbhSLWsSYP7mQu6YuF87imbYwE7M0kSgypPkacO
9VcOhv9BMfeqsHa4m64BiTzy+4IUdpu4vITdFlygSZvnHFRV4Yj04nDCylOxo/YQd4wRvTaYUCSh
CIzMU/7kERa/vP1G1ANBBl7dNfvbWQlrP3mYPvy2O5xL7dGbOWq2YuHt4H6K0UKy8RFW+ppA7XxY
qgiVp2eXlKnEi6acE5LXo9PR461rCzoERBk/5w0ZFKq75BYCuYe+kSeeJmUfVNufLira4RYgvBUf
Tz9j4YonZjI5vjy6npH5XbIGYYwAbln2xR919mpJY5kS6SkuYDZ0+m75/gg6/Ba/9/d1FLi2eVvS
nXpqjWmbnseP3kriCBEyYQHfJyQPeXn3CCp7NRR/99pobORpyPGUCcNYuYyjKZtoOxcCh8sl4RDl
hSBqsx2dqB3Te+FOMuhL3uMjuXgWIu47mi4yPiJWguWYiJuSnHAFCuJWoRGLMN8UAb0O1PNWg8q/
H6YdsKd4aDKWgarEmcUFn8WFdlrx3TeciTW+LBNSyQnbh0Y2acYderHorCqLdSRxgQstgiQ5CV/B
GOzqQISh9XPqN2Al+8Ecl11ifn6F1W3fJ6rivJjmIYu7OZZLl/Xjs95BgH+rDJj2acGUVuW23Ngl
6K7wmYKizzmlvT1Pe8TSNv52f8WjEBWZGOcJwbhufORlp38ynclO417vmINceZyGJ4eBvYBm+yuJ
Y1R4Cu+IJVavaRRUFbcZV4fcCs7oi4hokgsj6r8IHIuhtRmltTUpfEhuxJhN4ki5v2IBfEoKHonP
WJBIgemSi1/wWok+NlvZh4xSsa8Oj1beJ4Vd/Xawl4aeIoETkbwd4HEMrp9uat52tnVA4Zl7jkgj
0MXaEHaavMvyU7Z8oKL+4kHQ8Fig47cdj7rOHW+tzPVMm0TKfrIN6mk35NJmJBUBkaY/i74d3jDO
u59y60MTXMN53Uy4rsrujpxN0nhYr2Appks6ojPzyWvpKlWKyzE96EV5cq73hrXnpZTAXZSWEG8s
SrJfb34xtlaXmau2ZQf5i7bxS/9c8YkkyRAqnP7AKDyw1KAOTOmrZrFDr7t7oZFCZ5OJ3KvVlYuw
YucAHs7Ql18LicEbOYtip6JDql1F1u+6l/FYjaj04cSau75SxpgZEnCBEa4vRkZMa4cX6w1/6fHu
WnUM+5BeHPQyJ/a4t3Pln8cMXyu/F3t8jocTslhk2C38cRn3aG5tzlK3j/6JIhOqSO1n1LETzM95
CbOBNk4XYW7EX3pSt+LMwLZd3XXSY2cKtGyAXN3NciMis9Jlq6AriS4EZ0Wcw5fvazYq7AzErd+E
iq+gIeuIVrQcJQT13AXfsUv4wnSpV0o5StANTijd79m/N1n8gZ5pXzjCnNTJr7KE1D6Jvrx8le8F
OMW9SSLyZWdfQObl4AKCPO6333Dx1AQZQr04z6T+JapPYsdXOEMoxTO0Xgs5WusRsdUQe+5W/tNf
1ctQlt8F66NozbUrNnigrO+gFJeKdY96xwqzPQbMcOhe2Gdy30IaHV4MRCuU3B2cbTZYRxU1NIkd
Bj8pfPVvgGcwSTZSSyqA7gCMRg3CovvCExsu9cX8/WS8pWm0cRX0nITX7N3jHbp2RUio6rNJFMt0
xnS+jIwnOAaxBP8Wwn/rX1k1yuImf4iSy2ZSpGHwt+jSA462ce/b8/tbfinI8wj8pUnda712AdF4
1Qvr7MdgufxDFCpjw1tvU6UQk0ei85z4OcbW8fTUjBvMFoKe7XBn3Tv8EkRqfff/iD17XDg4xVZH
x6R8duF2hsLB9jlKdhmKTkWT9wWYUPaCSWhpIwitHbcfNZwu9+2lTw92NTdFtpw7GrY9FHmAwcv0
vvnYq2K/Zx5nrQU+IBuAq7sgUcwC/OZvcNbPJu50E0ukyDA0Y8vz3v+fIBNMyZEMPlpuykCGW2hs
979/WBu9sbkuOs1ofgyLxwrbwGXusx/t+CvdamC4+aUKEmnjtGJYjPa20E1xTVqcM+6GxsgqDmNb
XHmWGjoENODC3m5jl3Q25C1JIcb9VUYooyBmn/IkvkRWJMZAF1K6O/JPckwoYgSa0A+RwnGdWBQ8
p1F/DHX7fAANokqiwP83oGbJ7oa5d3N9VFjE7N90wtlinLrFC2Tsg5S2rD2hLtcKy3VXxMpE13M9
ynH1e65CC895asu3k0b+mhGo6MeszMYHND0b/L3PV+T4BuMbiz4+lvElHtGcoayaSjJYdGpzGhAC
MT8gMS9hlehhaC9y2h9wQxNLPcRHcPwiEu4maui4YftDAgsnFBXcMrIJLy3sf1oUy0D8gP0ktX6e
NF8rL01h2INAg+UFM1fTG8FxmWYBIuvPFLe3+60pPTKVVXFOyQIH/v0YPSpGfwy0qhhzdHikI185
XMAOC0LQ+F1b6V5S54d1WxSYhvquuIWelNGfkcSNpeCX6dRNDJqfiwudNQJG4sNDCDlGGhkm/LbX
xmz0kPaW2HChmHx4JJNM1yqz2L8BeATp2SJXXFmSVZp9g2tMJJr4ce5Ui4gziQQMSLj3Xt2cr4oa
ofEjYcWjGy794JRMOP7CccBFcOi6sVShYuPSLawBTAu3qoU564r2GcO72gPee/HpIsbLqeX0tQs9
p2a/3S0lou9TE9hKmNVOwHFBdar1XNIkJT9plqZuIWtXVEjJYciWBtzKAyp+RoZ43inP0mZl5lwI
oh8MrReFcRmqaL4hGY/yOV4VqZM2W6BNCc3WElIbEsuWVXM0J7C5CfZ/NqikShLLoqbRhE+IV3dr
hlgo2N4GjW4CHkZqPFLzlLEUf7eXnDHKLFZsdsB/QqoDvrHkZpO7RSkssjN3OAqRofLFolalLL9D
fp5ifIzkE5oP4ns4rnOx+bGDYylEZi6cPhCR5eKCVGY9az17zpa0a73soY5tnJFdC0rWo0aP0X4m
FfgnuBVzp0KEcPqdqFMYSj3kHw4lHyYYRkESITk/rlxTD6AASh8jEtSsdLrJFsU5y5YKpGTJ3MRm
KmknnH6m7nZfNoZAr4eQbiTvDWDAoqCUzTV2ni5DXMmaDpnZLOy5ODLQoWnQLq3mjdC9DKu9jN0H
Q+igrCCC6fj3YnCRbPck4d8Gy1OBXBTmSn0VKv24PozV3D91hoP3MQoUY8+pcZuclnwlTU2DUh11
yxI2wjcdE9JNGqQRwvMPyLbPFUHfeeWmVpwt+VoBQst/gdUn7EQrmVwTy21T+TjcgCyU0pQS4SNx
icgYvVAaBGdL+waiEzt+VNt8KUZqsXyBliCzdO9b4m26/5MEsEHZpTnQIxBm8wfsfE4fwABmtVvo
WzwpB/C9ra7pGy47NhJTGn1q7PSWQKFkTxmgZ7wG6uxTVT1o9iNN/wAQItEZHWTYZknJM/NybiGg
pagp6Mc71ioK6NdjhZENYhTYLz3pIDUzWqyxNwue9u7/yUfo1nN0XnkH9zgGK8J+00QkIo4Xvtx6
KOcomjwNmYwaTjZRQnKZTuBTPxqm1O9kXaILNv6z3wZMFd2gKpHqThdKAmY09rO4N2m4o8ExF87S
tiyp6VBLv2CeAiMwqAyb/gemKdbfDEWHsA1SifBiLuLU5ASzt2r94ZQBbt+gcZOebFzN3BL8ctCH
V4ev252j9oHtKO85/rIbaAviHSPBXyeZeSBuOqBAQ4w0ICQl5JHDBwI6YF+q1XrefpT9LUkUD/sv
eE3rhv+ggqSK7hQPrcp9+RkOvgIwmI//erVr7Pcdd6TBvFj9ohldSTIRYD2UNo264Q7kIIV0/H7Q
vUDI0hhqmThmgdFYaFbdZmNYVoNBUcm+9Tr/3Cg/6rH4iNP3f5QrPJkGvOXGGce20m+CmXMy4VjG
jaJHG9dvnC29sS9xBaP8tTPTn4JmfkhvVb/6QOzePq8P8nRBUDj+seRXmzKw5RCCmk1Csqa5GvDA
zvXzCNQ4TbnMnGvkqIZQ2JayIL55C7MiiqF8lOF+G0QGgGQujLeqtVCgHHVMt0bGnGptu6Ei+2xj
bkrOr+o39q0fi35uID3tX285HO/lW51NRyf1gvQGUmF4qKqyyoqxnFxWDD/1gig7NvwVag+27rM9
MwZuMkrWkmgmMFlUTtGbifVF5E7rTJFNhBe5Cxs1FnX9GVSvD+1PfrfpdsNuKfvbaV3wozmKWdzy
Y6+9YeMPoAFypAtU6lFeoEeHh7kUjpVizOFkRf6mmuvM8ekpZasBsyOuQH0v2BANNRoh+biGFeBe
3AtE4bx/T9Jd867Ompf5R6R9noXpP6tSlu8Gsdr6QrKIqjKfAva10tUQ71uJ8gSTxhM+JB1YMjqX
Pis4AmeTgRnUU7S1PJN7Pk6uBUSf3uKtB5xYOWtLaDy5jEIBbtG8aZKAHT57uY5QvjEnPqZG8NpK
r1wYUa1Jx5NUHFoyiLjGBeDndj1pFbfa8RRLmE1uMu0dWsz1p2gGpJCk25+LwogeucrLQLQ0dGwJ
uunTgM0VZ1DQDLzUzdjmmBAgoXSbYxTFyNImiYqLDiAf5KFP/HBPdi/enZI/6RhSLjU1850T9Vis
G+I0BCD9/kcEUce/GUArDsfpA3zvVnBrGeNLhAS6If7rllDH4OxxjUGh/dhJOMPFMf38WMSo8GdS
YRAPwVkFoPPoeLqwXAQvjFEpyBQgF0UrzhqnSs5xzlRD4mPAOYV7acXaqh6V3e1POXxenvw1Puog
KQj234g0E0aVA4Y9v2xD+y3tfnjkfYmZofqQkkakh82X57wVWcxRrEj+6zDGJyHjVzApgL8fiyiK
UQtDZqgAx8hoDHTPeBm3BflobuS+ZxzW2YqKX6C37uWSZNo8a+7cLAR3SN5V6dvZYPl7iCZPgjU1
p23qVwiYQLl/0jPCOKBSivrdl7gBP5eMT+/lq1GTn98cMXluMgZiyFsksp+YVBJIEVLWogZAYbjU
l3VAbvhKQdCRxsay9C7v8LBsL67jlRI1j5J9HXP9eIC/+FBtAuCIlti9z4hZGMoFkTFmRB1bZuYa
Yf7GztFNDZd9eKvYSC7ccvPSzuidHSfvwW6hxkIRs0s6bRzoGkHZA3dylV/EAn5o2GpeYQ+g7u6e
+YBUnq+C/3X2s2zWV/yPyyR5VZJdKZpqLZys5iq1vyY4Xh2xM8KI1yQEfHj2ipJW99rG3nZ32thj
2iWiv0XcJ1j//navTFn/fRDyt6KjiT2g2+bI5+7Ovs4Mh/bG2mQeUQ8VXS7x3Oe3fVrz8dfiwm8a
HzP94XTYKpQEfr5JJlfbPipw+eI2YHOrBOi2oaiOWVZe72D669ns9EE598TXyLf04oSw3F4ozojM
5hJ5zwXKPFuzigAIz3c8OaD15P/Vn1gn6h0cjPUuLokij+4EochfAeAdwjY248Jw2rgwwD+/lvJT
jYUt5+K8yRVIym6Twxbl/RPjOTOjosTLbgISRFsl4UCYwNO08x0jilOIsGJ7wFPID6j8UeGIPTQL
dWfAZMSgph/0QHdbFCkQEA/f9i4l5pj34eQFMEs8hG3tgNDQoacEudRhMxfO0em6re0q1jbsxEnC
ZI5Md47gC9LFC9RK5EeOj54Ha3kjKnllwr0r5gJAhQaT/+eGJEwpLKkC0g8vpLKbfaYzqwS+l0mv
G70ykNS5Qm05C1TPpClP+5idozpXkDLsqnWUsjDFAVD10LsXhAMS8FOGDSM0HGi8XPeRievD4cBQ
UfQddeiQaJ3eihqlfJa/wLIUKswLeuk4w33OnUlpAyVXiW+tzli1ocWCbfXCsHbfLUQUkkmC3k21
DmYhaL3weLCDzIXeuAVH9nUpNZ8SIAwQ2dTeT9S6H8HDNZta4BwxjLp6AiM8tixR2UcpveLZCUnb
iVUi0j1XTX7X5GUBEKVEWgB2JICzFseQjs5ud6bTiuclI5nQSIXHROTsdmeTxeSrdrtSdZnKcMXl
/kONLM2nOKBMrYwHwn998e0+aCoxOuGQPAOz3kBhmk8URUFx2EdSbJ0oMSt0OidDwgqqYMb3STVU
N3QU4vhy8iOSsD8B8SpGnDJZkueAhZlo5OUQBX0S4J4PVQ3qHdlQyjdrohShpL6Tix3xpu9XLjHZ
mqzvb5Nt/tgFPNgudWZNsy1uSsbiJtLk/scjeKs0KndswjWVGpdTANJcRe444Dfil6fKSkNFkrMe
roNJ/YBASevvKxobfMzjn0Dj0b2J3KWuXGahbLYAnfh329u/ZKMPkAcEbfceOcY6HLzA1oYoR9A3
nMlZXIWEDvj9vlpMONJCH/YJtXlHKMeo9CiiycWqtAl/D/i4aJVhw4OTL+E8hb6+PmyYTa/4Y7nO
KTatKXW2iZlag3+QLLOVN59+rZZlQjEk4vX1/kPJ8AWJQoOafQ5CUs1Z6rQpE+sDsGGchQg2RCv6
pM98I2zmZHRiwco2ImEBihmXV7GcsXzvAHc1pipCJfvk24hwtbGfut/isnkkaUKZpPOsrJUvBY+W
H9xqJ0gDk17tiGc56j09h1WU2OiHnwo+Mrv66NV+PcvCGFnGPG96wY4mNfVEQl5DEqs+D9dLlLw2
yHoC4d/ZBZq8U9wTmngVg+pQvsjt66Q1o6wkgNAKidGEw94oiD3HQUIurEZsWJCjUyC9HxFd5ux+
bch3xYD15YPehUTVgVywtHfWRoHpWvX9DEHABx6TpFU90ZnZwd+BK32K+IrJJpctfcoPAcgSI5Xb
ZnCPaN5rVnELVtKHIpx1s6CBE+v44I+nwBrEQV3UxxEsQ9CWXX3IN4nvucq2ZsPKGWaLHYC5H1jM
Z5WQjCzdOkvW4Y+zeHRLbJHMqIyPeilW1eXutyQM82d4uHD4qKa0ylPypA+0nfNCudaN9A9JccS7
fUD5jeHH3XZyv+SaRaTO7QHDlG3XJnw1K5YwUnp2bpclrKAwLgGWffiktRE6aAePumF6zKPIIXfW
5w0wfSfbbntc69tkd1GY2Vttd7F9Ebb9cOqSBto6TdwkSgpBojSzOudj5Ao4P0qQD4JoLu0AaD3K
GM9/63+a89rKktWczUdoCttV3To8HI+qNVhzU+1O8w7+wK3EhvLwTYqcpDRB/dBKaYo57tDhOtTe
VD4mQX5/6t8r24KZeavcRRG+7gWXNYu1vCYKcClONI2hrmqibf1eAmMxQ5yKAdKVTNwdeCNpKHiH
G9vIomj4LMgmqbJX7jQ4fkXZRoKNh6rKWIVAyrvUcFidWnvvd+yhZzm1MixXxKyAE4FL+uuahLvJ
taFYvEBxDS7B8DOALX96Mw+yPpDusPGdaCHvItwG3RUQNRTVP7hYZntccFFYy3j08eG+mQ4Svxom
q0zS72fp37BbbwG2uBuW9QZYn1ReJjbxagjDKN5y541ymHNGdYKturJ2Hefj7CHal8OV7jn64iq8
YenNCfAsUm8vyd7VikkguXjoTh8v0+DF1nnOlkailEaptdvehrtEbLuF2uFDqpZ9p04rFd+m7wNV
CnXjzoqtJG0FwYsrKnaoD+6N6iXH57PoYp3JoHLUvcX3i4luZAYYgR7NP3KFJpBS7Hpi1p6ArbmY
vG84cbgCghJiaQNy1Zb17hFvjCoQ/KIXQ6vKqQy6XRMVtCYyDGErph0Sbvx7HXkY0npJ7ZhjgWDq
6YCd+cp16vbpj0kZyKntzB6v9hmGps1KKYUHOTyaj5AGq9QsH353OxHdk2TTOSNhPOxSpsSD6nP5
Frh5bvIdExrEzi8AZ2j61NyGJ8cYj1YMjFTiO8KarVVIaoX+uNJILmjesbWBU6/Kvfmy2KTTDLIO
QD0gfzSWrJ2Gp20UwPTEmym/nzzG8wSEb/rjpSqYYy/L/tEqr72fBO5/3iR+pmdP7LJdWbIuFQZx
1kqUe4Ksq9g0U2jnKSFpX8WdvkMCXX2cdZqf83mCfQ0HX34exkMRFxyLX/KqH7aLPz7BTWKgaa2d
fLB2XzjOIKJWTITj30LJ55otebWprBjp8QlmcoSv2y8P9UyisL4DwdWZsPMnt4AYX5R6VpcQyHKT
brDQxeDaSK33za2neNb+US2RfWj0jP8ST5eUX0dkYOJpJtjOUGgryAueR4/vFzgGvgnG0UcNpO5C
5Mw9ozUe0lixeS0smKTbQwE/ONEVkeE/NIqNBAOzmrX0Gyx2NK7OukRnmtEHiFZn8DMvMAtYe3GQ
fRnbN74fOfk9Y5PvUXYL+aR70h7H4BDEOig7ecTZ0zYPX3jAetol4d0DL+tgmjsR/9whIy/mI8pk
vkuo/JltUypJtBN9z+1CE8fYA7MJExmc57H8bvLXGsobFNCSzrp98uw0+XLRvY9EDe6jjhIN6t7i
L4AnfZSMhdr0HgMtMoZpKfsU/1CHSeYo/ua3S5MY4vID7ovJkfH29FNxu65M1lOtVYBUVo0xOwKF
1ji6NzdrO14zDzYF/SbxMVBN/lV/JtIzisJNr6kHOJFU823R1S1YPW2o/JmqKBA8kX6ISNMuewyi
gDyCUWbmMkPjPA825moftagAlfUGexe3ld3mXjBSdbHKbU5pFGZnSKxK3WPWb+KhTWg3z25cv6JH
Vxk+yjyzR4H1h6ac7K80txqoPfvbdFEndXWqzfw1WwR6o1CN91hzMDTYKKdlYebHEZhsHzWudzb3
OS19L9oJCWlPN7FIMOG6VGc8HYWk+DxHC2fgFrHCSVNdcpx26BMIgR11A5uE0ywglH/YJ8vRsslC
gBxCjOKSmKg5j4q2jhTjvF6kIMSAP+dQK0j9fK1WrqgGp7JUeWoy+UYhkyzZZuggF77SqlTC6Oj2
smTyQraXvG6nH49nUpxq9Z0I9F/CEAXx5QuMzmtYyzJS4jc7+Qd6X3zhlxzA7NzgUV4OFqyex+mX
sRmBCvEaft1rzuUBftUeMdoobwGawjD2hr+SVZJnieMqudmVHYzfNZXH3zxeUdIiJ/rOFif0tjJm
t/5NmVhnjQ1sz/U2f6tUHi9GckQl5qHrenTLhmrFc0KDVRrNMblX6/+hQt00gRbxcq7tWUQ6myx4
Q+soczg4XleLKNFxGuq+Txs04j3YaGR6WDuxCDuSUYBy7GNi9Y+QpzpxHNZctVoa6D3qsIyUZk5U
YZqZPNZuhhkv3vKpxJ+K1DtB0bRZMyH3q98OVwZ/lt/v5SH9Pi/jatJ+DK/l3Vt//gShf/JJ9JLt
TwH83IQ8d4zU920iW3MOe/AYaiJ780WaWDtM9IAmQoJtwu7bE9ChTYUA3fl0z8eUpk9fxTi5jX+i
UR3RIY6Zof72v4iuuq1ENcUYqtY9WPP9g9yQRkHxNsFQuiZPpsepzpf9/JpVaWGqWSsdhX1sVivS
SDEbC6nTSgmBRDdWPBu/R5C41l2Mj93d3sOHhXvcznwPrY0yzibWoOVMR92GTg1Km/NyHwIADe/B
nSWDLgzwzLRr7mrklIgvObyOp4fW5gCJQS/vs/M3GW7eL7AQWECPmdQ8jKQUOC76rQZTKKKfZOrh
QpZOkVNE4rojWWOeYV2QS5fOdgtGAQr4x2Ipdvw7PueIPtd4kMBhmImwDlIImzXl59tBfKdgrk4A
haqw9XIozkrmVaajsfcZAwUDGRj+HbuySQbGsKYAU+KCmHJsP3Am9ye/yP0HYKHHG9qTMiZClb76
0T7MCG15qP2SkH2hFUN2zv4OqG+KvBM7ywAF5tSlWlp6MVNtcg0fBm9YjhRUrtrVbuKXvdMdHfGt
diA41WGer+gRF8uMJEc0jWwBfCDeW93f251fNjV3ZjEPS+4yokEy3wYEc1R53Y1qcs9w7Bs6g5qC
My1b7fmHJau4vGtEp4UVT0gjE0owy4fcaFY2/4Plo83Cpl6GovJxHmtvjp/VZFLRxsFCDnvjmge9
gjVWzkuTp2n7lvsfQYFQfGy+doKWB8cxTfer9j1fbRqHT82LdGPwh8rkPMrJSro6aaHgASHkMScH
QcWs6Lv11nCDbNohtvENqXIGOhjVAIUiwl+HmqN52CifqXUx73nkxTv6a1Rvv/tFz8zjLcmXKzuG
x0LZFQz9ivpFNGxLzAVgjr24iBxPVLHwajiyUPe2m7KXSNTTxJ8oZu+xzXhyrKBsvBYYF2Q60ep5
DdI23SCH3qXsMH5llYAaaU4q9ppWMC8JSs/OP2U1v72XJWKDnclxouyM/906X3hXygI3TQmxVTEZ
HOBkyf/yyZKQjSUQ9bhSHSNf3DAXzBzy0O3MwUqVoFzEoIp/vRPRjA8oXc1ah91TUbon3G3lQ3Vt
/Kl54Wu3vDpWCHnx9V4ZA5bs1WYQ+cVoVAs8zQCkN6asDofDWNhHGQlNMI7E6wAxWIUQ8cVu8GKZ
GuXJ6vfGhl/l3bjrwzsXOwdH/CYCd1boPOoDbTwIpJ/VbbUgT8lfJMDa48F9TGJR66vfJHhJ7Rz+
EFnt/gCxh/jnhILC7fwmi6LWW3+M3S0wF+L+Jlosw+Odos9x8tlPNksU6ZhIIFfn0hoN8asTYuJI
f1rrRlEXRJa/7SNdQbMcKHRYMw8Jugv5cTVksJTn7reyVaRkAvkIaW/HbH9QYYDVnTa6RnpzOXBC
Ql2fNkAztOk9v44elfmAaeA3JpUUs/iN3r1oO+tIpG2tjWuNxs6zm4FkuiuBugkEjGh3CB6Hdh/5
tfAaL6NBGwEXHX1DlJP+xHqFhfaXFXGHy8yniKLNNmn+LbakZ+F5axSVDqrgTOifCJGvHMkObNcj
NVUni/7ZupZLWyoplPhe+E+Tn31BXFBEiXTouOkwW5ExkvbdcgXPqGLcaXKGihpD37SF+JdJlNw1
n8UaNkjy7CZ/z/+02Mx22vfhzc8RTS8vocTFTBDj5D3V56O883Bh8TouWQidefKEKpvABy2UwncS
q08M47N/DCE6/oS08KXVniQZwvjlzhXtkgkZw0jXqF/1vdgFYa/paVis1xX3ukXEWL0nxW7u3U9u
oRQ7aCVXXZuKDzT4HEe+6+UVRC8ozGU+WegFixBMtw7zBgWJmelg2LJM4FhoO+RsX1XJl+K3wUqQ
9d5NCgPQgLXuwCYZ5wzqjt5Aj/t/BObj/3TMnT1b63N0xpXqcuurYvt4HlrHZT97pu/VKQf8wEGc
2I4MoCDE6sJX1CDPgXjmKaLC0GRoSILoQ4tBe1HXC+I/fZeM0XCx0WAXgU+bdOeHDJha45vVR+dl
1B/thjttLdEzNxbHmAAhvM6wxj5SlvXSLbesqi1l9V8bqhYWiZMV+cU5xdOXvvuSuF3aIu5ex/Ju
0DNYDmTr4pXZu6qx0Hb4kxCQ/MdyIgf59zhEYDpVWSupZjhux4on2DVbDKx35UAEcc9L5gyu7hjR
VuvzxWM+8SeCKTJKpR1AYiVoqNNZDPf7YumG+W0dh6GoI4BQUM5kDdtyNReuM8xAtLaUKAz++POM
CvdmmJY2T2P8pkpJqP6lYv18s1L8BwVVCNVNfkYrCAf5rffgZzu/XKQlNCsJF2rBSRWV1ZT+0EFD
P+ff9/1lLW1pxb/wa0HKBwe1peSOK/8AwXjcvgBCD0c3cJfb67nYMJXkixM0/hPN/eGBDutR3qRT
jWFCAlG55loWME+qRM8eAco3MCnnDJQptwUu6pv/tPqm4LnyWaWM4rD9+IC1LSX2AvWpqjEsSyGr
NaBdjQciwzaXh/9GTQAjaSmVyd+B5o1lqr8tpWH+7FrQCxq/md3u/aMCbp1CAr7ect1MTS5ZZxfe
celJFtq9qdrvrS9Gr2mFoTWsOnt7aG514xUuHCTSnU35+MmBxH2bnX05FHEJAZthxSWg2cKjz+MM
Z+hCCmBr790H70ZNLndpPo4sy4tdO2eEwzouU+ZKiWIT7PQk6vNjAT6YafcdBgps7JU11F6ADra0
t2BkhN11/o+IMXsF8Wj6N1mKpwtYHpVwysEnUvRuBVHOPuusVCLBnUBgKpnVckP3Y58NZlAa3kgE
B+v+CqrJlca0+HUPVaJ4HORg3jxktYdoRAxV5OF+CE90h5Rzxex5lg7a8o9bJGv4scfT+5ME6HSc
eLlSv0N0PRbYxZsrWGJHHq2TC4Oa0cppezOce1rguogtjooWEIMLp8S8urLrnpTmAHH5NxT9P+ox
MLkpiBSNO/PpeQM+tmH7xdLX0Gdwo7V+oCwDapxSEsFArqSwfvdYczasTKKMsOgNCOj94D2NORXW
+X/aYUuKjy8uyWlS5hDV6LFsTpTVmAElG6soqkZm0qdO40hJbnz9mfrQDebPmpkRwozKxl/KNbQE
0VA3XrDZ1qYgFZecK2J14W3/c+UfGkz+NNDPCIzpKWrM3e70ekMrNT7HT8OqUPrlg1zCOXNlIU7/
VsHOwTSB+YeD3UDtFvdRNK0g1m3BKGNybRxzsZ86ePSXdaoAPKCziyDTU4yfp8N1FEGgzLq1eoyg
ra/JAnFdcr2oao8p44OtNAIIvN4C0ZarLnOx3ly0ClLJ5btOgV4rkRwx4B2QgxUvO5Wku3cvwKTM
PRq9zOjnMNs1eWkN6YLnMHYSojSZt3GGE3sDtkR8gun0QQfYlt8CnHe+0S3yNjLAzV1XzEQXHDbA
PEyq9zHblD54d24kol3SRo7wsq2xBxRoSHx2Nq/PymLYAum2KEqa292sYDT21anxuYzTbU7D8ECn
7S6Ksn1oAJHWvdd7CEcvkxQO5BVj7vqCIAdNIPkikiLMSw/rNVHFcTEnmc2yIgd4gtLT9LpnDPlz
XrV7ktHivI6GKL0zlfrRJWWql6H0Pz8YwScw9WxqceADqwr1Dp+9MMpVacIDDvshSZH9ANHU9Hmu
8JG+vyyVNO36LLsoJ/NmiCYBK4Nure16hGAsNaxAODQ5jDPDFc/ZR/9NDDkO6mQFJxdl4t0oOI+O
T15z05aHuFgpa+AvSs/4RysJHQlQxNYL47I5atxf2z0gOVMb8A70GDxIl05RDLIiMEF+SocVWjnP
kZmTAD6Rpgmoum3rESwx0XwVjRb7Y5d74GRORM66kDHJEiw2BzcXVWhX6zq0wwvF1iiK3VjQMDsr
I1yniW4C0GJy+xkotprXJg3U2Zhu0bNItsQoyhz7P+4pCz15jRhn3a3oKTrOYId+sFTf74B7Ym7g
nasCuHA92qRP1rH7OkFgcg3Yc31VtdcqemEKEgLjNhiGejA28N/RctAhsi21pmmt3Ep1zmQ5nvzR
S/hNWoAxeCOLl+SeL6r2P2jYl5KhZcVbAOxchraNNb7JvtuYvUHv8LyFiziWLpnEErxGVc1DlUJT
EFyhRgifFCTxudYjTExGjdH8LGQ/vXzOvNM/KV598onjE/dA8IXxgMhEJpsSGLShI9cts8X7qKTi
RqhCxbwMtq9t02urK/sK+zKavIl82YElqziCtJYkmpXvqLsqO3hyjRJO7PWazPTECnvMnaOg3ykr
8TS1Kq/6iWxBekpexaEjS+OKDPWYp7IAu9JUCqZ4Gm8I/s/kdYx9E6BayjJdFsAuSO+inXPvXKef
sVXSin+7w+Ze9eagYzE2JFuiNPilz28OVB/1H7L1cE8aT0Iy7HVCp7Dg5AS9auZ5P76CsXDwxjXw
cCGjIOXOLw0bZ1QZvHmFvXpcAtGoXqrJ7TC+kEsUh7l1ANBxjSi8XT7Q0FUtq8vIDAXjAeE8AiNO
V5794DLAd7mijJwiMuFN8IaijsukHt/3eClSfwauiL3T0WRtLfPx6gIDGLY6l1SQ2/DVZ1wxuJui
xxIvRzIOX7dMfOutv6ZN72dR7qmMNwAyWLwGyi7ZubB44rQNX514433Gj+v6Rh4Ku1/RqRxN/PaF
U5v1Hsh6xEZdi6pgmQTa3ychPmpthC0YgfiF4KtbUfFp7NYA/J2CTjQ5Kw0LVg2tbnrnMy/iALHQ
d8sm9Zs5n1XZcIvfkr7/NKs0+tnKt4TLN00bWveThSiHn9csaDK5QNO90r0//0XF3f3p9g7f9UXe
W8zZsEgNuE9qoqrVXzWe6Gr6BBi9eaqAzOTPsn/R4wdBA7//bAbCptFiaDgn23xfJ3ETBsQwHxPE
OXCqk6xIFdUDPB4OF2g6U+LZ2f0EQ75/0W6xJJ/PZHpvZ0Uoy7g9EW2ouA5JaSk/z1hOWU3XEPSR
NxNu62fD0mtPfJ67mtdH0Yqx6EnxTw0wHeMmWkqOaPmgdckBNtsjYz41SSmVibXhIVXTI6lG+9Ja
besXiaUVgPJypi7wwRmO/F3VrCyraCi3aOTIV8SMZ84OmsPZ/AMGIijrPDIk4Dci/aN9I6qm+x/q
2jrJln2w1Qp6ueDTABPZJSu39tTuRbilhgG05t7TXmq/trvx6UgtmnpLFvZz7Snsuf6yl1laarbB
K/qyesB4Y3AcCsHGjYP3BiXujEOzcaW+zAUPn8BWoiZzsCgqtC4AqXOgtoKX/rkuOXbui6tA5b/y
luhtNBIzQiOhgolh8u2ba4yXXeRCsTvXu5CrXSbIe7OEdEWJ01BFldYL9xFiJ3lf7j5SBS1s1S2k
pIVO0JazNbrNHIVhenWCFq9+cjsXyuvLfBIR/UCp8RabVKpjB+/BT6zf+RRkOeM8MKX1St8Vnd86
6HLsLv/iGIG6OYcvMo0UHrojuw+5kMLWxc8m4GFmAiq22LthbPTM47kLdXoQ+Sr3335OuvHGQszi
XCsZMUNBVfQHqckRWYmijXkj8O9crjOi9zg2qsOkD+V5mZX4cAxQzl6jtqVSqr+/icvoqqK00MU6
/4UkkjKsEYvvgBTj8J2xj1ODICd2t26dQs9hEXZo+c/hLEXEPDnlHOgWYL4/Joun+z5jp2yGcvkl
9fgrdxgQgFCgg8hDMxhdThS8uJvuj06yIYW9QcT0NtaJ3PoQgcc5brwRb6G4qV++N1ey6hb9Z1NP
4xjYts8EVOTplhT3C3uY0V+AMB+fZISj62lkZ+juFT+rdBYdQazBqsEBoL9gi3s1bNj8ANfQV11k
7fdHpMt1fSytOscodSXXnfYgFmruAlivXAJCDWnnTrnVd85ku4zQsKo/6nIfh2TmeAYmPlzSUhCi
7r98XM+8RNC3QB1i5S/8Up4EM53ajbpAphzEdE6WKHopIL0fxsSDQMw6FIwtiw8g6WlhOA1ivH7F
CD6mrGuQVLeEqvVpNb1qaAg/klMk5OXEyEUP4SxYjrFmJz0PQgl6xllpf3f3WoTz2gefosZWTk79
IzPlx69qaf/NhWFoAf16Q5E6C3xeIQt7skp3RoWaWEBKwhhhi+HW+akQ5WhejkvDqDqzq2/x+JPB
ykj3Rp/nhQVv+fnrO15jY7O+SF6ViS9ywCY0IXWLWxEMvkqF6nwk6IHgACMxdbA7ZkmqNgZ2/4Hz
wlXHwPZt9NkEbYUrSRQPSgQOSRSnsFsCg2GhaqRNAE6xeMhuLbAqJSMJur/yUqA6+PaiccsrYQpr
/An8T7vl1NnF7EJin65DqmWnLXQ5gX0mWO11ZjRreS77647uFosVPbP0Lv3jtpwSUIjfqwhOuTYu
bsbrowNYR6BoWQAum4Mtr1CrPuRUzMA5UphRej/YfwLO+KuAUn1w2afKMDOA3LN3ka+LvtnZ4Pfz
1pvsMG5zHRGarGhZfjQj5esa2InTrXEN/trOKmtGLjDWtw02p04W4FZQAOxwJnI47QLf9cLfm7fQ
edefTEQHTsH6VcCsaR6WAA11M1nF8Ld68i1THSjaVTUTSVKdQDMQKrdjYfW/TcIrbHUsh+skpKQZ
0G1uh2ropaFrY7GJr8QgX3BirmbuO21kcwF4z3Nw/PmvuSwmmztTUhP7Mi0bcDhTFRUuHOgVUJ/B
nNwCKhUp/o7MeQ4Ml+7mUFOIYUI6ceVsz/mkOZ7VZSfd1pQiQKtk5k8l2JSZoeqyaomYyTtPUakA
G8rgtKVGZSVn2ZCF5hCUGzFzVLvdgX/GjVqxgO1PXEKWe34PoiKzkPwwBsIVYv6MHRGeP42Zlnne
OPhptCLVf9id/OBT7GUsppajmOfHrtb7DmRIzxxyhIrwSla3e4nuD+JnhijOczFZyzVDWOfkx3SR
9yN6fEtdvxj/+KH0vqwdN2sNb5oTpEuVkHYoEGTxejTJVJgEfd1wWeMmiWojsct2cLhvJ1ARFPoF
ke5MfoGt6vNJMiP/QGqqib5LOO7celato77zRh4S1+fQsOyO2Yoos7Pa/LwUH0+xHPy8eiosgslt
yttGdLxAJ8fPQZDZDzz4ZvpkutaqwMmogSWAj4KlOHGcy/0s06Rb4v8N0WxQ9IAESw9/1+qzqlgl
W3n99uk1KFNU+HEdiLbVzj5r9VS39zr63aFWCn2/hp1DeJAneuLlsAR+qQKI370hm5BW4G8r6O83
zkq6IaCLkwjbn5A3tI/pujvL+7RKZ5JGvMh8MW3niYZ24JIt5WhFWmDEZ2+kRyZkvxTTXh/cye8+
Nwoh6p6dktMEzfQ+hwTLKmYURZKwCYr21TuKUpmigJ6jhnq8/h6DW+JrDo38d3nUOCPX86jA5ft/
3wcG+F4wRq0cCge+0i7bdkHE+jCbKHXS473Gxu+l6rnnTViDNKWu4oQMdsZQl2ZEw6H8VfaGqWlc
XQ4IENjtvRRnDOExE4Cu0OvHiveSvuTNA/X0tfwQe+M884+7MWIMEHRdvk4+eFOcqEKtoWQeD3G9
q9fVFgqUvcAzv+r5Nv49KuXZnIEm7GjAXvlqh0ycUvH0689Q0o/ZJgQNFI5IGMoloYQkviM52EeX
W7f/i0NWxvhDtx2yzCut8XjZQwSuI1V8c4yOLx+KxaGD9M0/3XcwVFaZHLY1YaY45ZyQFVYcO5tT
fjKsYW1mm8ZMm+Nyxm9iR0Jm6bi5W+xqqeZR/7emk3Cx40a3MbqaVbZ8bBnocMFXNY3Mt9t9CXsX
XZIkb157N5EhxBWgsbxdo+LGsKGPLVHBY4Nhp0D6GuSZDn0ErDqzMltGXh1UL8of8XER63cLZ/e1
qpZ6cBdkNupJK3Arl/LKWPODOQl55M5xnAcsLXhuqQYiq7ZQ7XjiE4Fn1iiY3/j3UOOv14c6/Xx/
zUuR4n9YLQvDiWJIah9Jqju8KfsflTDFPAbiMVzQ0S8s2P0WEgLuB8dHhowqSAYQSoZno4YcIvG8
Keww9dVHpEDHS3s917BaLoC9C0J+dMRTXsy/bF8l2uy/sHG6E071eaYJFX1zN6Wn+ip+OZp8cqTh
Ivi8GG2srwdHwIu34/DWpQh3yx2D8cVvGXBbhkGgx6v3/kbT0EGaZ5ImyM6kBZ0kBtf1NSp437V+
l8XZoqIpZo+xxDpGXg3dQclKZz8EEtbxsaRdS6boji8mfgk1T3NFhxu/o/CraWdBkVdxhiNmknoA
SaOBc6hOptyV0SvcCSxZTGqmvhK72DsQUp9CkxQAll66tEnAf9IsRMbOhWx8Nd7wdCstpxCTuLXo
YLJQVyswMam64fB7vWNYyUOnefHAmNDe/9pVxQLF6WLE8k7tpZ+6xLqwHHNFroNcLnhb5ou8bwCP
6Ew/tNVHx515X53T7R6zPe85OzfhSF1T8DuriUUvmacL65sSeYT3+ALiZR5BrAmib71LcK+kPunH
RdPON03Gn43C9V6v26/lnMna1guXYqNuO+7gv+tZcjki4xLkz+NCIGVYaFMmc2wjNMWBuaBkDkY1
QZys2qWOm4MWYsIGrzXV4xGS+7KsqlEMT+uPCLP/f6HhUZlRijB97Ih7LkuVstGd4D2GoZ5376KM
Rw+3sVe/1/55TYDuM+m4Y0L4wXIohagCY9203uiHRUZnT+4YsnHJu+c/IXsucBuYYN5wppysijGf
zfZlRCBp58UUNwfT4j9JyI+aEDUx3NfqDl0/5sJETY1kex1v9zUaSUMAvWbyU2fl1Hi0qzKWm9XE
Be0AVcX7GIh3K5Bd4FLweCvzr54ItdTsDxcb6DxhK9rBjfi9wIhvD0SL+SsIM8IMsYykiKkHtkKy
ubr+y1UGmgjMU6Drl+BDLAjpjge/EcAbZyA+WuQOsrWrMfjKTCgEnH+q7NKcnYEz+D54xjqSmgT7
il0CveiTpOECdkfTWrYdBzW5OxERSGVOKuBZbkNyzrgZV+wa9b0zRdOLqRLKg6qvgpawNpLyjjqN
pUsshd8rhz6mmkjLnOUJTxRB/E/pkoDeb6xXOgsfSFL3P4bMsUqWBkqpX/oobaHFaLolcRqFp70D
cd3IB5MKxBfi2c5bPib4q3tx+UVETxpGVxPIkZ7q37F4McDWrkjLPD5vVylpzzMDaRi1vwJOgU5Z
sEzXexYfLoB1erwvtTrfjHZW/Nlxl64wdB17wDh1120tEyHVmWMlPql22lIPMd3mQw8OMGbv0Rzw
7rOoSdjpcq5dKv+XdQfyvOlPUH/FxL18ubGPTCECkaZosmyF425uPhYFapNARoY7SMSgOWIwwR7A
UVoM55oBHEK9d1LUyu0H6uswOJ3Etugbm3JXTQr5fyOyhG+7oCzTjIZPaXH85mG2HfV8xtQ0LOUu
Cm85i+Vy+brRnHjlto6gLux21Eawm3Vv1+TbyKYuDosKDnrLr13ANzc9LBnmQfL3IlnbFKOQUzdd
ehRvpX0fGhHeBhRk0oLsBtFt9doXxKKhatTvnA2D6C9rbx4Qi4BwxGeNIjdZwldCfRRZ5RckiRy8
cKlAr9wjX4MMFFpLtolVtkpEiqB+MfWFIkVW4GHdWDNt5c3uZDNAMap5M9EbZ3xNayW5JHWaU5ay
rhPTZGfdbao3AkPr0UsOkoCndwtZTnbX9xKTLkfTIphIQutiOyKJROZNzLmZxQMt1QWKZFj+9Q8U
TloghnJn9oqvYi2XjDe62P3Eh3hwG6JINMt3PvlEAvrBjoe5PrJV+9D5SchF9RGoGOAOuGzbFOGJ
djtUsYUXQKqf0lwL7J04T3uB+0XRtuldtWbgKsSvqovRoUjH7UGF00VyNSQxbu0rpiyup7C/Aj7Y
pTLBV1FpVE3JS0K3XyQWlIVQa+HvYyJrVWqpU0uWGS6OhlfPZ+WWht24kR37QK/2qNF6mIdWFZsU
xO7l4fVPn7SaTXGbdxWmEFAyoJZLmJimeN8SjNcXqy3wyVSq5Q+Th6rTf/UWsHIdGSspgvusxExn
iMmGV9BuoCaqji3hHveHoPZoR6r41xdVcgOEWTN+rDhDU03GAc8rBMOWfcpuQh87k0ahT3M5Tes6
8qqWfS/mEZUK23xvh6QdCSOL5RlY2vnA/LSFZ073gc8htab8Cxk+2Q8EooEoee4BQ90wqFSxOQkg
W7okpZmxaAskvdNO5SA/wWfAr6HnwhcRBuPyV88dMkBxHB4BzREn9ZH+aNzJ4mRrfyt3n/Sfa4hv
YwNFKA2tA48yy1H/bxfu+93Tc9raXr9fAYO90meSxKtDMewUxeb4pa5bZ38f63mzDdjveUtA0Gy1
jj5xLHUag6oaqqQ/+nVxUhSQyV5HDIk61pgdeOajzqkz36kEHdPBdLrugUiWHbuVsedCKhsq++O5
7Ae3RIdSu2plwbWgE7tg9ErKVP7g6NPRrQdcl73k9GbaI4BA0z1nws1wGl1FJaDCNAOxImeyVL8q
4o8nUzdchXqwAmxvRepqEn+0IgGd4IJ9gW7UDOESIIwon+ScArTEtuFrT/fEjQTjMdLekt5du5N/
vL0nirhvLpZuzaw8PTWOWIJ5qrrXqiHi42mNXLL15DZ2dCfM6L7oyPRNwvx8FTnvuj4gcvIvodUK
JhntEad7W+PywsZjl+IVnhmgid/j95MqxqhrbO9I47G8p8vNCLhjxTJv+SmFol+W7B2nLu4PDGIN
vJ775FKWHmFfPyqL8NeYU0bKtfTZkUS0Fs+xe/fdHx9jq//Gn6A7BFRRoV9fxs7Ob+y+2nX89xTO
8zF16ckCsIpDYi2xKWXB7i6cxUyrTLdveHQWxkKjzhAz/gRshPk4v1tGgzhCZo1e/LZUz5R3/8ba
klybQP7dK5uDEVVCpeHnCmlm731Z56iJrh1+pF+C3Im4jb7NHEdalFhvxY1XcY4Og06CzrYBaQi2
quUZfcq9k/x6eENZyJRQIrzrUF74ZL2/dvZQRX24oiHXxerVusD1QeEaAG+h7h/GA5wgPfuRgWum
lHzAWWaA5EdhJ8Qi3r9LRj3v1bj1YDA5fi2Gb0dRJa4yy+mYYhfx332IDSq8PIz2c/hLoVzLjOnz
9dvziStFKf6CFsk7P6hB/zxh4ZoMwsLbbo+8BvB/xt93DO45wONxqkpdbAXbWGQ9ZuWSf/n2o5fH
olktVizc4bLuZcbJpOfgzh2QxLg/BpxfkDaCAnhe7XsowZOM758gDPF0R49X2zp+p8sDptKd3FAP
1a4M0hZsTgJSUOgqmmBXF0cxlTo+V71YlT86KIbRMel3jgYsL37pNIUkYAYk8vPL8fotcOvBzOlJ
SZPSWVQ9BFWQHGpPNy7JsbzQUfTTPwDMC4Uq7GW2K6x/hlAojydfAJOn1c4HifUpYXea6zTI7bRp
ga9UFhwwUlqmYgQVVUy1+/t5oS98/MpTmqwYYbCd1zQsxVbp7zZG6ZOjh2YdStNPUE6PLj2brrh9
iKt3P0IsqfxPDEraXh4aLU4rslTv6GMwZxGzrHn04L4gUKgko3iOR2BzK+S5DXCR+yD2f3o5oP6S
sx0TFTwkKqHTR+o4YOPgnT2+snJDNi9KmqyBWc+Va/6o18T554/VGmps47PxBa9ULdmsKiJ5QapJ
icFlhiyg/N5PAaQYQXHlio19vH3r078QwiVzmA6gn/Hr8flrkjr6xJwuTuPJ6GKugzLR5a9VEYXn
/5aKqDIz0QDAY4OrHMMJbIalaV07pfrReQCNyoZQ/VwYHuIZVIe4sayTVWVIrG3s6Bp87I0jX01l
3WTYuV6PUOf+2+g/XXUujS5cteSU+nsvokVZ/PlZuTssztT4ao7vm9X0gMm03gHRGu2maDCQ4pTo
aAT5UpHWvT4ke3YIsle0ACjvLd04LjA9G1aP0swy5+GklIH4piy3SHv0knrcfkX5+yUplyorkhau
vczge9dmH59PTW8GDq4Y1zZF9WQRnjCbCdYYDJq3FuQFwBt0Au3oQXt7k2/B8APc1cE8cquejWCO
iIoJztPwvdq7+55Gz3/Ijtl5vifPw/DGVpHHT07TbCTTzEprVWyp50qos0rUH0H7N024eg+yK2Em
J6jrIZdsmXND6iMTxe4FFFR9QLAz1iUVm/CYX8ArMK08uBW0PYV2Gso/wqCzn9Ve/zWZT2Z8MPL0
sXKxjA5kXwNICbIir56v7EHB/oIXO6tZOSRnxHVkQoK/B9nr6xju/BMW+oU5XOemDQDRndo/jfh9
6DOaeQJX7Jb+uojdPb7L7AbtoOzM+V9iQLiyX2nsXG7y1tiPDD8gZz+cLlr5prmhtI4bK1culI6m
P4ZLDJe/i4QaNHGTsIE1Id9Iqcd5H6Bpkhk8t9CGSehm1VELm44mYiFY0tE4ZmEhd5IYm/7sKL5R
v/4vGOCdl7DcH65xmo8JgB36HTR0Qk3dxKbpCJt+z0T1anr+02wt84AwVg9hjcA7dXbAXXNhqHkW
OWuhBtzUJ9IMaDgcAc/EfkZNdW5qz6YcnUrjkfgddmqpAfR7/1szKz0qRtECUAWlbwAhOsc7yECw
SxEwWWWtzaNBC0Wl25APSErGW5ZJiueqwACDg1Yg7yerPwsvq8qTDMNBYzxL6MFN2eaZZfdc8FkH
WKGXSbAWdKZNAeLgHl2DCaD4WMyMiJ8NBLOIJ3KT3goKjLyNfKjbD6IOJ7LjoPsclA4AnUHu/XYB
iOUdqKJpHGbOu1jIOAs74F7Tp86eTznF1NzZV9naI34veVOmWfUQZzz8zk7OW1SmEaAVu9Giit1q
IetQaaa75+DwnQhtgkHBf4wzc56231xpMcQBz1zjxwW7EFIochUmVoYczJGArhxJDF58ruK7/7Pq
LwJLw3oAUSpYMK7wKR3BqLJMoluT/2fbWvQtxk19wqT7q7NT0oLT6twZpFtS2kv6pVgsEOpwGt3J
DOmegNxcmCrggNbh+S1T5GnUmmdL9QBWidhfx9v+7qvfYzi0Ps87xQKC7J91ng2Yhvuu/UTreDEi
LH8fMrAH6sDI58vR0+g+03RbJZpgb0LvLoGHEnm4rbmD9aOpGoSfIl2LJWDpKmpQc+T9bdSychsY
0omNwf0i/PxHC/dzsTJAiZT7XaqTW+YF8lk5/hjWNwZQQbY7rF4fqNBAXtAPESojBaEpNJYem18v
Nv0xQfafvFFjUpFUb6pfuSZIHeoKbayHptMCmEzSkekvNNtVbCwn0ziz5OUbLmW8zgZwk/A5IlFK
1B7xfI15IdlReXhg0V4rOBD/FnicNx9Afa2Wb1kqR1UyvEUQ5Rz86oBx1Ns9UdO8SRO4Vsv3E8D7
P3dTKwmZoNhtKhXuyrhsT8qd6DuRK1JqxSGT1wIS+EyJ/6NRpvenu35LERxEVvH1fu2krScNICEW
xzzlHvGo6xO0B4/TvLvnwkop7aER7YP3Z589DgdFTEcxdJFW5kNWD9zGV8dThAG1HjadoYpCqpzI
8B8wnTIURCTo4huO/Zk1ceoxlvmpfTJKbuhwaxm9x4cLc4ezM7S14IIGXKqfPsALBIOkEzRlbe/Z
NjiftSzJA/IWJeE0lcNsFfnpeLIHihpdLDUoFz/3lsc6tVjBsxmMVv67HYdMFIIa/ntI+ATGk64/
uyHAMMvQTrV7sKWYxWDvHwjQ+6PJz2lxBPvK8Bi3JS7CG0qVraqBUBhAzWMMQUivzyUKI+ljg0Mc
EInL1DH4Oo9aIkXRpSm4+xdOkqeR5xBGVcZ/4Uj/t0u106kYwKXoXIE7DR5liHNH1x/bU0FZ/74z
/Q32HZdXa9Zk5C62rYXZoCKvfW6xL9KasOw20sDMSyjvOH1EDdZmzO6SQaKk5EFmHboyqhUJWuB+
ffuB8Q0KRMk1qug8DTsEa4WCDTJHhp864V8qY+HXfzSn86Uchd68DnzvcLTrDD47Q2ISluUVpgF1
L9pb4seBTdlX9rw2bV2iZ8SyhMpjmQD7Ek8/hgBB+4WMrZk/hE58V5p8XHGy1bICD+aGtCCyRpsd
wu34+BEoNxeHBFUFNuHIJzhuvip81h21mUFKoeuhZRy8v0Feq3I2Iw5Snab3NeXbGus0lna85p7f
Iy7gPTnd1TSCiQ043VhtWS9fBenKGJoF3wk6QZeLTn0Hi4nNTPZsaCQslwzN8BR1zfTOkXIucDvW
THcBcLZ0Z4R/cHedsSug4GTNqEeidDQ2xSZc8IWsYQYcHg9Aa9w3SOwqD3q6biQjucbiPf+41lbo
eL6xTMPuqF5xTDmXWD8Uc7XYI5mPrei2okSzq8g5EWwz1T8OwtXTITya6I6fTssVXD4FyHxqHqih
1myZHx2GntjZDadgJwNjgtPQWvgcwwBnE7FKTXQpqAx2s8Bl9UElLjg3/mT7TcFum18f7z4/Y8tY
DRPQMJ1mrO/DexgDIIuoWYLZu7xTw8+NMRlPrQxMqKnB+fOp4vjT1rgpUJu9DwjaRFyjNFzkJ2nB
pu3bnOwtY8JBONWp5o1yKDr9XkTAsDPUZ6CTQLaSJEEN6/qp3HBkwY/dYS6IInlVrtw1+WDH/MH6
8Tve8fDMsNCXk29uF2m8vK3/uz895P/4hZpkG6m5qWdLdV6AL0e2KNAN3K9n5u/hzH6TLJT18kml
btYkHlu9KXmCiKhCXGF67voNvmTD5bty7PfSqEC0lRlQp59UFs0Wzc4+/rsqE9x7R8rtPgRJCyIb
JW4OQWgyluNb1BaPSKTjSdDOhpRYgbQOqtmvf5m2EQxsYOs4J2icybIywfw0TwXfZJabSDbn37a7
Nh9xIv+yZ0j2JRhxDU10YXdd0fQw2vWLjBsSAY+O5cYz95C0vjMJDQXK8swu9adKzzEvTtD8ADDM
RTDCrvesJ+5zn1DHuNYJ1b86+WNVLi4Vz24ZR5tcRtPbSRVQi95WLTdSodEhsZn6xTXQEEp/twNw
HNPcxb9f38cv7JAa2sVCJfgp49vAviaNedRye3wGo9k2qgqVYU5eIeCZpDsi0Hd36inqqkfLpT5R
itsvMxYiJoHx6rnFHOvf78CHsHk1N/8cF+XcKGcDutr+R9BgKeb+2Ohsangg/VKhhcZKfIY5EcP1
J3kaYr6B6JLEfIR4AtuBPPsYFuYfJQX0kID6805CJHlQB85qfcsdo0zTTtjKzRuXw9qXm0MbhkQx
zacPEXAxii6BBw045mkm8YgUoECJXhWljZAO5EtjKipr5x+21VRAFxIS56v72R/oyviay028Nxex
vahw/P7kIcg/LBf/OPxPhs/lA165GgF3JDN7WYLrwe74r2F6rk/6dS1MWFuoszZk47TmkHNVnp54
O/hY0kFfiZZd0Eap3hNWhTx32i2dTrmTXEUd15Ixa4TakBlUEse63/6u5B0S/kTZQokXiVLgEVk6
TYqj5R/uFNk3tek97KgwLxd8gB36IZ5a0qclfSVGce1ITLrSHxA8bin8gMhMwXk33itXqR2L+PUz
ZDvoBEKRq6VVksKPUbCnsylvxDlX6VCLmwGm/PmfeHrGq/zqhsXQzqRgxzljkDIbYV57rClAakF5
KRNWsDE+HXb6LIPFzAcTwbn6UE9Dos0WnaCZ5EP3pZS01sWR0t+Oa5Giz7fhF4lWsMGe9iAzdLC4
F/PYmDXcMU+pVHBvulY4FuBMYA6RcX5N0pFbA7/804aXSlbQOnfh96MEaafRpWQgDc+GqXWJZ5B3
Lm6lNiCkw95O2LBdlOVJc8Xb3nf1AkR5UgMKh0caFVR5CqXW3uCNMf0XBp43FkCNndtoydm7MCeb
8b1cpSpUhQBwjgJTiyor3vjm3bL7vVtFH5wBdymT2syjhZQp+8vK5UH1tUGB6AOhTMekch4lmQGT
Jb1/w7TOVMW5VH/dxxDrfG1J9yrw5rxCTUWb2wBkvyg+pEYCrqIIIXtlAaQvj55TuADgMspvL1PQ
fsJrOel2tRepNECx6fauTmeV0eNKRvl+ERyRMeYsOolXftyIPe9gzmdQPWf/ZDVluGRy3dkeD7Bc
VuqMhRw1bgz6s5rK1LiWJyrxyeYZ4rgIxP4qcMNLWju0acEWQ4t+crVaXwIEFL4x4aGxn3Al7Bx9
bbeGAcSyNNBS5armLBzZSIkAN2IIIEu+DnstbLlz0ltG1GR9ZjEAq8J5K7P7J28k/+Xy/sy5BIPD
vBKjUGxUBTyUnBJAml1T0mqof+CZYwaBlDYpEP5EFJP1Z7QcFjIgQWMK5i4NfoFrUtzLvkwuIaA6
ZWgcmri/gm7xAqz9s0SKsfgx9aKNBeU8YrxFI6z2+C7no1FaVC+AHw4nl8nTB3CIbXRYUWlmu9JA
reQFmuG/E2v7uxmsOSmEjjKPUd+L6oHT/uhkCM+q6q86IAM6FePwtvsv4ta9pPuWukJBmIPon0vS
Cd9CtUrudfWw5sS1tYQ+lMFeA+C67Islnd4MR6NkdUkERBkMp9UeXBkOYDzSoaw6OBPw69tzvMrF
jDjfEnhkP2nHZvOrrd0P2yNUW1mXg4qLuFbelg0fiSMjzwobOc6RH3aho8HUOXTVzj7+naQ5kHC2
c+jM78v9S+n+me5RtzTR88xpY9sDnD29gjvtOX4uX4AsaLPlXyIr34OICKa1yBR0aIrZrHa6IYvb
j42P612d9/+BnuVWxoNKirTLv9aTz+G97SzlkGr5+8Xfkbt8f4t3Zxc4txNL9eGBeZGuIPhayELW
QHQ+SwEmBxZvhqEWBN018bNSShC2KFwJ5Sj4qTfPqj+f5j09rERgvk2Wzng9aDcb9/G18UJDpSsV
IE+P61Ix92EMkh2PA3NS3ti0rUqNZ3ohXMZuM4BR1u4pc2ZFmZ5Szv1BSHnxSzQ2PwJTF8XDGQFd
Tt5wWVCbuahDlQ3AOzCtYiGf+13pQgB97xsgNhle5EE/TCSDWI6BQmqXcIejC69+lhVNoOOpqreJ
wrR4IufM4AJO/DF/RG2Vunou0W7gDS+PR5T+rzR7E5VZTa4XtLh+QTzQk80q96mTTEPb74/9xxVr
CFx88xAeFoUtxlzEFo72U1DZzDb/EQrQL/iPW74cg5ITVZUOmG3A2JsP2g+29/cxwqtuCt2faLwY
9APxpocSlr9uZshAemnO3GrKpKg7dMfOgwKVa08ISF1b/bCE2kzwb5iX0erahrdWS6UuYMmyq85H
QLjnsq1Fnt8T21UFML2H7XgpGn/hQS5IHTncd9QUAc/HE2l5AF7v3MoUAE2ViTKF60UdWAQUR7Fm
mRjsaY35tlz2YvWAwR+CAlEVrivyZfDhyuiDpJbxJiP1+/877KIA4z+IKg0XFw/erMrSnyrvni9x
Ri9Pdg7mJ8v0uFI7iJeKxujtU8Henu2Gtw+CkcMzxJ96tvzjEGN00+utPO3MiSwyLEtR98sSUGJ4
sns8IXOGDfHzDV4svRf381uYAG0ZnUjBtt0nbeLPXaneXAtqAeVrDMlac2ykshLuYiKWuD9e14//
ejal3PyiDxAJmOeKwbL4WzGyJADObJSZm5It53P9CG/D2Wg4fFFtjU+6Lm8mByv9eZvr575lgWM9
r7+NHAV3Cy+LRlNsNTdGyqIwcHTxTivNHrvY1I9CZ4VRwbpgMfvl7Vwc6rfGIr7PBUgomi6X/276
KC+wHq80MZk6QHjKCwvX4KfFzW+Y5XRl8g+tJd5xQ/+GpB3hKh8vwmM4pA0rZz9gov1tmO+eRDXw
43TnxIIhaIZI7XjkVbNlLIe+/b8hz4iNTZqNRJBqlmap7oIFdTWslB5h43JfBGbjHoCDzRoqKq19
Fbmlb2+HH3jg7gbynyvdWtFSJMuKpOTCkBuSbyBoDFW9lN1D8dV4R3hNRkz9gS2TXshfSl+n0eyS
o9MHHpdF8fWWL6k4klJuU6y5AASoIdMFGe2FkJ+H0yOakBWXhApJfNsu0Gymz2yB2Sjbh1XZb3CE
akeCFmv6tSTqfiiVkiV+uII38MvAW6gKB+6mzQIcsy8c9QM4dDni143iVXNzC0VqPhd/JIpMn23w
EsH7X/Oa3WkyCh1n8ZvPx9H3EEi8Inm54ArLf44gzjT8XU91p2JPf/0ByoM8I20t4c31w/JLHgS1
BgJrY8PFUU4tkZ2ae8VURqujYisAKybJ46Qy2H71GSiSMdzEva4/8xXMu3eq5aCojN05tdL2l71V
SZqddRStBHbUMLC6YktlcUELJltqNftfU+fwy/Y/6AOPE50il6U6SZcjq3eVtoVRLD+YYwxZFQGA
bhZj+AYvKLJuuv33TVhgNvUye0ikVOjyEUa9iFdwWyV0iIpW1HGiSOLy/eefPD6RlVHL6cO0hgl9
4NS2LETYsv724N26I4NxxPBOaz3412i9PQTpGRoMfhiLF/TTAJKHlxVLXwA3xAXN3VsuKOxQzYzD
VlcpIdw+73DeZ6MjylKW9DBH4sNC5JqtO/aoGygtT9xgcxNGzm7pPrtptKmgAqZHOzkatZLtv3BM
0kAzdOWF1YJGXu6EF4kGBNW9jWl8m6Jvu7uqCvhyFsHU2/tuSDNbO9yESYoZBDlVmEgrb4o99tCO
j6Px54GXzaojGOm2Xs8Vmuv00DF5v4aseg4xXNEKGm8nSpQwPPNR4p5STfIFQvYczGx9/XlLh8gk
o/0OlT/YNAZIepUgz7GYKl1O00oGzfYuCQEpnJppFQ5gvwC6H3NcKCgkHzIuctAgKAa9jOb35qma
SJBwoV0hAYoysl/k9PerlfL20j4o9SGglJa6hEAM03UFeFoc5QedkLB50csqN+RAHlkGvAPNXSXH
2+Jne1uq0E3281TW4E50uJqRPcXmXSuuO8qOG0K+wnmqg+MeD+Z2AbQnFNOoH+FLbKitj1ole5kv
mBO0rr3PN4e2WYEMFIgqZ11d9J540ivhXBPR18WeQrANczW/ya0BGy8TwOYchAAqSLCALygVnCDb
1uIeDD565co3j+HeHp/c86+c7ayKi50wbVz5VCOOwp26/v0cFa+jugg3mT2qR/9PfqQqCdGPSmub
kpFJwy6AeJFCAq7RKEpo88ZomiWZgWnLyU0Hm0RfRvYh9MbLm1iGuPqSF/cbKTMyktBuCUaDxQbH
8jViIc1IGhGEVoMNMOKOgOZ0xozDtM28is78TzuZmspWvDT3XxVcgOLV3wJwoKt8pOSRXnxe9i5e
YDsFxc3FndPEioMvuUeJAeGE+F4R0lb89057aA1b7qTelV/txM9x7eCtg6AnEfEFvjjo4bcM84ol
CbTylGgADtsfkJZ3nvRuuXXG7EYVj/WfwlaV4h5onHpbOk16sBK7Y9YNP2LKU2Xi2TQnkZnRRWaG
ZeCx+BAn1pWx2Y/x+8OZii0lqSl6rwmgx+fsvguSJvBk5SwluoHAg++6n2/hhF/BS3OOKHvdLj5L
Op22vj+BiZEaVFBoEPKPU+iCiCiUJq5HiTXwZoXtIxc1WWfQ+tIHF9yjJMlqMZ4BExBAEqZrOrGT
urDi9MqvZ+dmVMDw1GUTDmaYVZxYRPHtj9QolQ5Cw97F+KhmYoYSLbiSTVGiOwocbSkg9l/J8WNI
SPEpVsVey8kCJOv/vYD6xj++3qby0Es5i24yyH7NHZO1s9KjwGsy+dFIWnsKtes1kQteeRx2BWq9
A3xQz0EP5jmNJM/GVzmXLDkWVMLCVAY6qgEsqZF8+TjSFFB2oe12Fo6Btl35Orxe62yvLE2KQaxL
dEaWPPGOP4xkZwwCQiWNXmMz2wI53IIi5mFUBen4wxst2hOvkJn+XyS3oGYMg0nWpfXTYbjnkJRe
/SX9towzw4/Z7e3h6E85zC4tImIdVDy6Fyzakk60hTVYU/FzFckWBPy4Y1T0gXyjCTfMlp25efG/
EhsBNpiJ1mw2mviBGhwOcchi7EuwsRu7PmO6wltHeD64Q6KW+YQEnRNCnMkMXHag3acCVj0QUDLt
rBGfkv6hNS4YAAF1B7r08cuczG4uw3BwO3voXgSj+sw9m0jUAQEoGEmTiuzj/8AKmS0NrCfCgSNe
tUfxbyfw/qGPv3IzF4JhuvurvwmI3iQX7YMjzOo6osP2vD15qIfeQr7zo9QUF2HDPRfhWJ10MnrZ
GiGHYbwthUlYvwEXGAvAcuuwxeq8lJ4/8YwTetPsh8mE3dBYcKm+LVi+K0qn/OTRvNOlyEZMvnQX
IJLjvmplpWAnv1+KL9OzQqEsmvccA/Q/rUly1GUVZOPxhj5WUGBnW7JQil5rDZPXoSCTRlF2BGgv
/tThiKI+OyK+jh9T9Cm84UuzdYTywH/MkgoLL3rj8Qp4umJj2o2zOSO2PzHnY+r2NojHnoUliB9t
91+GMKzkpvh7JTaDKJcGHG0kZMkrRGWgRmk09nKtcdlirSrYO6w8JlQz+9wTZd7a4ar7zsij5zss
uraiXctgQf7GR4as50JnIRstioCZ9j818M0rXEiSfYgrvxq1rzctwXBBrNEsjMH6a6XWlNWKjElj
45oBc+9me5kken5382T1RhxCNnPllgU48ShDM9PlCCbJwQoXFpqT6S/bdT0Tr1Sljq775vaFYySr
PmlMWjUM6/L0ZEaT824Sp+ZbLeRaTm39McbssYry/F7XTHuTuEd59S5u2ecAjdyGrNdNmnCCjVby
Ck+/XaZ69o1y29RKkUexFEnThCACB4F4JXBbel4C1WqOsTTQ9v9IPC2iDRaroh65V82NkdVPwRLV
PY5M23Gukal+Q1gfurk8DZL9VRxQdJgfscNAuRHwW5eEVDf2wrHbpPOWa58gYlvcyNA43yruUDoi
auNWM+8+QCcxPCIMZu1HlqUZuFw9Opygw5dJExv9TLQ29f+BbYAjoABDopkGia37G/kt9LJPOe9R
/RbSb/60KfcZ0zJCQF4Jkz70+xkqJPPdXBwGHy9iSPsg/n3Noj0llKdmZ6OraJyPiD/R7UXTZ5eD
M3EiRYCaxH13HzOJoI6SXjeBkaeEscpMRFAOwLiSIZhcu4OhK3f0Wz5weT0QL7QUZrOzeYQcsl2q
348WjpupnywdWQRU3vlKrdhzD1GqVCmEVhVdImemjiKmvOA1iqsCrYkS+NuQDC6Ca7s4Hvf5Y1PW
DvHgYF2iWCQfSEXY3iphose1IZBLSaOtFcBvuDzDJgP+QiY2sx3iDNgdIruyHZT0H3rAnEkl3zxU
f0u5HRq0SFHgGcneJMhNj4m7qLzcI1x8Z6RKmf6mwG3jusoAmLjAOoDIrZTeBCD3NrOMuRtYcTG5
qcFwdnEoDhHtFyLtFuQbbcw9gE29se9rn/ME3PDJw0IW+7WbJEDq7gJ4+NDZM4k7HDg/avXGJ/I+
ioyjW0jq2SmIZIp1xxQozbRn8NkY76DGRIVOjkxRmjdUdPvhIDC4C9mY0ZDmi1kJdCGkg0fyvYN9
ia7oBrBB9dk0vAON5rDvA5PhWxdPUUk6YsiK8eDcYyhXpXTxt//z31AwMT0SmG8lGlOD1+yr3/kK
G6gNJeEJt1FsuegSkhsDaEUTX6+isiRrjcoWlEqSLSud7PlENcXwTfcB7VqyNG7WBgiEAU72IH9S
+7vIPniVk7NMBKBJP7T2Pv+SpZrdwFbgYjZnJHsun5Sh6uxGooMmj8MvFrw0gdFL2ghHkbzhuOOt
tyXi1ZnyIgNhyjeV6Fk9DBKuDq5iF09tRJnE7du/F6PIQLb0j3zM/Qy/v4MZ1YT2iOOTq2nbNYyj
Xd/T7xhkQP3YvcLkRA51i8umzZeYq3PMgV+EVyPs2ouwqXAqJeyyRGP01PVug0CnHb4IsqoB2tb3
rbF7GrOmchnAUEYzRaMevj+jAZ20TAy5dDHu5z/VGickvOWG6U5bdRr+lKQrGLIZiedEYVCW02x9
kCVpvAoWtF6e2txyQ7psN/fouOb7WJsGqxQqEc3QCPklY8v7oV62dVDeFjVpii2BB0sU1FThmC6b
oyyECl3wLua1SrGoV4v8yb4aJXGpOs6Kr8b9diTN4861P7UU0kzAByEnuSgCE6r4qZKoHpxAFVj7
2UdmVXStM4br04PGzC9JK8L35NN0uz5DhNKlo7z0ORQbHW6HGsoCaERQfbU+aLPUe0Ucg3saGtfD
HxnXf1BjAyrO2qkOQVAUIeQxOAD9nWjJd5yjMMhB/gmhUdSjloZ7YJrwO5ckT2/0iQVa0mvn2mEI
vDc7uvPedeth4URd2LfqO6hkAX6P+pLiWauTm2GPKu3dpkiFb1pSWnyVQ9H9843O9zkSqOHtFe01
56L7tsHpxaSUd4fjxVyUZZNVwOkWPR//W4HnDZVjfHxcGhtsxpGYqt81RAr8BGMY3oVqLVqRVNTY
dt+oRD7KiJSCn9M8rTJ84AOEch2dtH8s4Re9h7sK5XiTIUbMEqHYP7uyqKFogMySe/YqHl7Y9XfJ
XxSmBk3XwLklWan0TCHZbcR8sBl8JeHxkRwfB1CDiMIVR7HlVOXkwlp33ebch7ciitbIIyj9U9rZ
JWYrTmQBnmX8N+FmhNerQo6m6ieOpowPAqPa9JYcnvRCEGM1B9sIc7POj85PLS6emRxxXi1RjTPW
8rjY2hJ1D9klhQVCetNKEUBRwYm9MgMdWn+nqxpYc+c5IH3Kfd6ZLvILUXDwlYvV6I/rmcs+8j28
UCZHrrS6PHrz4a2s+6KcEtK2T1oXuNdOSTQoyBuGu7CD/ik1lu2kuVaylv+FBepDg8k+BY5S4ZN1
LXnPT0y/BfC6HEv8afYfMy6RbkELxwFoYlPq53zCHrd0wIw2u9F4a7GAbemYDgeqZUWC/rT1kae1
rQadh+VcYWDZE0Ija5SVT8W+pHkya0m8dgQlpkbtgw3dyOxkQRuDm3F5po7ItqjsGA4JZJ6pFCSP
4orAl1Y4jNtxtBsAqaxa3e9/sez1Ck+R/IVGRVRy1WGO7caEv6/GwitP9uexi526lOVgZHW+NNve
GHfw366OnRAa5Kok081fAA6kCpzuhiujKa0xdkOFASCTocVFYK4KXaG6Mj4pYr4T2jWb0nWhfhmc
j6Bzw6wKWryqizXBNXTMSdcYnTnVhwAPaCFSjH5jj6f2wZAJ7TGg5BJpzfNpHZRsQm7Rcij3Rk35
RJ9gWVIbvmhk1BKeGlTeVqOtVUqJZz5rpfJnVTGHcNfNcQiFYiiJkIKEuD18oHlnhghzbhEXVQlS
2TbeIlypEXeHgvHlznQAL2CijzI4Ao916dzzcayjwJYudHKPlB2zERz8jRY/4sWFAuCbp9m2E7Ud
YrtXth+3JQM3hXVqhqs76+JH/FPvTO2jhXtSR0rVeLmJOKf1JFN8T1iUhNXxAlKxyr0zpgJAYXfo
hc/DdsScsvq32V+//ARGTd9xvw1yZeMWGwlci5IpF9ljSfLm5dvQ4NxKm8aUpx4u5zduqXTBe1mS
bHAU0jpl4YdHsH9w5geE3IwiiIZITaQLPTi043UUD2/eEbce0pNJ4/SrFnavGb2zTfTq8rcPr/0v
XUsYRjjVE04XsaPGIYqZcpgiv2H3YXKg0p4P9o+0i4Vaep3X6OKy77XZSRA9fXjb9B8xyjSCc+E1
6blX7VqkhGodFLsynYpRNWIjIl6yb4WGOrwW6v4JD5YDIRl6G0LhqEMvxm0IOIAZAYayUyBFaRU1
SqdT/m+m6jUdpMPvsovVxD5jGPinrycSj3k24xCzoqO3fGbJUQSQcq4ZlH+5OaYKsAh929gICR+R
oRkCGQZaTJGNr9IvMMgo1rUcADVCLyiiCPnkDesi0cQakBe28biEEz/zED2gJhQaBkT4iH3VRC/2
vYnAfktVtkd5xHUyMVsn0ZaLFjJQhScgrvGUj3oTFnnFdnwvP0eqyG6y1vLpQapFouDaojL8K0uJ
2VK6OEi4yNGISUlNtMP/QyvPm8T9VYD5BE+7i+0qPn+nUVLfhLbw4ABXZhApM3Lv4sazpYJieCSs
mfe1+J8NoFApSxvEtz3r+I7huxTazDwHU7kwyP3PrjhMGG4CRc/YPA/7IHHxClR6i150oMk4hwPg
YPee9DWh13hD9XOP9uBbJfEQxFbsKH/7kxMEQknuu9uK7+ILIvxXrnuXba7HDpDLfbBQc+PA579d
kyKeYJdZ9o1AA3DTjqeWxqM05VDA4ppycsONi5mrw+nHVuF7dKEHAy3qLvklrt3x4oBTtOGF2fSa
mqxVgiabiihuz1Lg4Ig45wHPS8Csm5WqPv9p/5dHZticNACut+za2ebLL4ZFPCDc5/Oq+CIS1j/C
uImd8Xh8fOcRCBqA+zvTit51QxB6gccUlpk7C5Ja/lVEQPk0IfugYP50lZmqWBqll8XQtSpPhxZ9
HjLK0hnqyFoeGFA4ehe+fBFnBmziEKKMy6QySXN8W4jU0QKfF+SqMv3V06ZYWUHgQ6U/sxnG/8xq
VRZjTcq8kM3hUW4p+oXEKAePmh8UAOvui4ufTihlju30OfiHRfRr+GAO8DTYTuAbaFSlnIUv48Jb
o+ai+V+Dj4FVoBL7o7GRDEj25y/O9h0qlb/OLKFFiQ3w6H/2zulP9HY+z8eidfh7Ied/WFqbI95z
fNA4peMul5v/D9xDxLw298lCcMxQxfzEiI/qlSZQNU5OKtM/+SQ7zpqiTx2r7jVwFMF5FWDsjFPJ
a6YpeaiglCiEy43Mh3sdPyOPqHvS1QAZlqvOrEVoemVJzBLE6OQatQEyzhQib2gfOYUdZRlOIC2e
7WAfYiSc4rZtEZQdpZNLvX3XSg9tJCpq0DXbgeaOYzeLP3dBie4oCcsaDJnBXtqxciZ7GYOyv3qX
aeqAhzyOSvrqKZY6cSoNrl8RJIAMxfU7itkOuCqBtsYDgYQjcn6e+MOVyAiAK1qBP9tetY3ZnZNf
Kr0vv1Zdxc9qRe4kc4EvWEOWRL0FC7vcvTqzRQragH4u8BaLg9fZnvvn5gfaeZ47TzHF/nvQtNw6
0XSp/kZkDDHxskqbL/KalctJak8XSTDWJTVPk/RT1HS7oMGMlUQhc9HxGJaGQ3OMKlAtF+8MWa0o
5HwHTLxVzaZfKT4KVUz8g2zExl5TU4ZfIwxNz4M4f2GrjU8y7D+CiD+GhDA35TUiU+AEXqLSmIjK
WBnuXdaofRhx4uIYaYVtHIZJomPXB9Ng9i6TVx79CuKR/pOmqmJQxPG7FhdeCVPFmq0LxNXE2Bc9
k7OSej6eUSbWEoPNvcdcidVE/pDLQf7uyAJ0nXsaYtvByAPeS2rRISmjbdy3nfjVaKnEH7tS2NM8
NnJ5QmgirGWbBQ0OP+FvGGWEkGqMwtR1WpOCEIUxC7+xrOh4QDlz8DqibuxfUfhdjx5a4bRu01ny
fu75XtL3NOtPNQJexWRz7QGR6OEFaM2B7kPay8kBGBKGOU98d7Ff5qrscSwwEMoTAaTWY5CRq7hm
q37K/QqYSOl7tpmDghHG5ZiWCTBv5djcch8O++xSOAZjW5VPWbtQG7W9dmepOV9NTaz0LTamsVEC
byW5YAmrP/eGrbwrI2tKgmc7VYRMxiT7SQg+QtfKnSSt7MInbNRYeIrfu70KohiC1/lNytzu1sju
B2JvDEJ/NVsMsBv5Fb11hcV++VvqSMLIYJ5de3WZIsiPKPiBnjFRWwcCgmkoqtsSNb+F0AWs6ChA
RTQ/J/1A+/xEfxcS0EQB3VLgu3McMXlSFAQQJYFI9CLtOIvybhhp1QCwSk1j/iX+0/DXefIyNw6Z
uKZuPBtdb24pPrRks6XjLoSTB2rf4nPPC3TAw5vRrqoWt0shMRCLaTeraUAlLkFmrSVMJrrAb2Yv
fnZi7qwM0jAAkSru/QWDrsrixVyrqZtYmy8ouhaOnhlK0vHxRgAi5iHuPjKZJWiEWcTCxh3GYRmX
mBp2ma+IdpWzELtfwrWuXEGfbYwYyY0TWS6EPYSMYJhcAIAR5tRn1NyKJzQz0U/qGj+awCNGd0mq
4zPwdNUjwEewSE3zGJ/GX7g6sefqaATW8QcIHQS6BnupVkiW0Eee4dPzoWq91UaO1w17vru6lQAb
rKpd7Piq7mYpI5ffg2d8Xw1iEp4ZeulC9iYmOEZr49GNcDw7pzIvpJgiPP3UNWZhPrbAY6M5Mzpj
4SN7fiI0kGwgf+k7Hx7o/onGxh7Ao8GsSvaXn5em1DdwIDjNgktgC8VtbmIQDdXF/+aovRAXgiVT
xTYXLb+9x5uxIEiM6dyAvzZFsMhCL3LcZrsPYF5LGVb/RO2XaQPDGsskTuKRu6sB7CTn+TSooDHS
nbRD8Ua+cJ5GKAg9HieZVO0is7fNxQZQ42FB/n0hQP7pWFhmlvzRjX5YdxRbqa7Cy+dloXDTiIb2
25DxCoJ9KCAhds4W607/PwN1qtqfEIm7LwqWwXEZEbCHI5Fx/rrSlIibyBPn72PmsLp5gJAU5haj
PN2AaHxIRnsFjZu9YXye3qXCLgWknEXdEVxVmTB+mmoZqJ0t7Nxj78j4P70zDgZH25fQeSdb9BTr
aeNvGG87X//9P+rkBfJsni9tZiA417k8HfNUlEDhj4Uss7gpN4xVEhWMsRx36mJesWIHPNLeVYzb
gbsHX6j9ggDYFfTiRLRIZQ8oU+oOaNpWTNCqVzIuz1YVXplwhqj8ehyLQFzGEgIkbGG83xyAglh0
LlaZ3azyRoRl8Mvmx9EB4yj9o6gu20ppzfLtzpumhJuutGSkBECJUAIwIy2a8f9Nke3PPVA9m07Z
J/7NPAIjir30xBJ06oY1QPzVH5TAYWhYP12hO69oeEyT8AviPiWj+vl3Ewx3g7vO1mXYw5py6/YC
lMqu+Fiv7qLgE9qknYZBR7huwO9xOoUb6Agyt3prhbo8Fz5IwbA8Kp14QxowUykuZiBA9YI81yzL
38qbWlEJ7Ok61aatQtpvdvQ1EI8DImKyWZ7MHU0QArkGVnedSop/zOVS6JpbQm65Un+Z/eiULIdx
Vpp9rcEG4LeVhOYZ7bWH4U7wNipW2aUZVOZ3S0WDcagAwKWV311Qja5Gfj4z0zS95kOvwc0iyXL5
6vLgcjwCg2lCK4QhPsBSDuDEcHNfrLHfF0CpW0O3BFOqxoOJxPNBb2Sf530vCakP5WXqtmgvLn+S
PkTaUb8P54Ah7vbkPqAy6giCBOQrEG70aReOw0wHZ55f8etURiBh/076WN4vkIhP+1gA47p6fwhd
qVy5k6e2XzVxpMVGc5W3alkIDj09swtV2yoLnAIpIUZ+jEGvJLL5Wnr7zPmR2yA22wrGRK8soV/+
hBHgQ6CCbISqh00pXmkh9GRTmzQwhh6oyWwP/rKCOSp/QZaT3Exp1t+8vijxBwKy003d+lxjzrVj
VTt8IbDO7HUhpFGQNKfWyNwEZLbebXObRkCRfWLerQCEHBjgbdqrbpikOJd1nQXmni6CQchj6wdp
+5aTdJ8DsFbUEdDgR19k5xWZZWa2TNYHNpH4PaozL3+UswshpaOL9Tl+SbUw+sEaKS6oCoLJ8q2e
9aAWtieYxhvf3OXvkRswyoYj4K8zYi41XKpHviu66J3Zk0SlgxHqrsM+eHNxQDnXBz38nW+y72pp
RDlduEE/IRvj73Gn6MJuLBHN2GP3I1/ivDNN+V1q5Bx5pFIAG7kSeCF3M5Lo7bsnniu7tWycaq0D
bgkPL1q5LkzFWtjc7HWU61LUHTR1kMP+bSfp2lfkCyFO/Bn47xCKcGXNVEOIy5TdPF+E3NT9n/8O
PJhFAqzgWrlvdcwNPyRM0p6P22yutd1OjfcjeQ5ujulLdd17Ts9ITP8gI8es5tBl4PVGkgHKt9Zc
evaOwpfH1pwP4PSvKBjBQTKJPvK7TVjGJDp/hIGc6EeaoAUXlU0V20eiAOsQBqwcoj1oIG7JHCDW
TUV0M5NOxZQ7Y0cvtJ1V+htw5MjlL5eYcQItZQHipcQKMRVuzfesbiqh5yITDwfVCDqwXhDOEDmt
TA/yVAtLzSKBwWbqSNGz2eHlnfDCZ7ESP+cBEiCd9DSdmKvQV4ITgTBneA8X337tXe7hR8VzDoG8
UdC3DLazfeInhFJthw15bSUsJr9RaC92eLXbYPT0nhg6Y26YxPqJL4TNs1/a2rWz5idajDDXraxk
74+ag/MtFFkpLQ8tZMKHO19ZB41UnkEAD5qcPNCW4d8kyF51Z8WKJqj+rxvJp5rX1yEa+qZ9GYzA
aExtf/elJZZ/wddu10CZVhImwULuhIxzrz98cywtT86bp0rZt6zIJptwbgqzH7QLdcyoUa3eDfbA
gzQvJROleNVfUprAZsFgDqO7it+7le5bOrJH8iwjj7R0XGiW06uUwHXhrKjHfIPrYWlLDFKl5PuK
mH2eaqSvrVSSqciKYBXzwg4/vcpbR37Bh6nZbEi4AIjWanaVZILLU2sUXfp2/4CFiSq0T7r9mL/C
MHWCsRorLHVg3rGwk6xDKLI9o1uBsuYWHm4lt+ye+WQkOq6AzYjFx3Sp0hOtFtdnfcIRPyaC9Bs/
Fb9vDs9kYe3pVwLSx6yx1eQxv2DuO49qiqexY4wmnPQJUSHSepKZXInrA8h3PT+hqmV0YrvtWLFO
wof2RXy4XSY/TlAyMDmJuj2tP2IIfDLZkYTeIB4HhWJexqXi8alSIa2JYx2+T2BJIQpp5Jx4XUao
q4ZuOAwt6ztymNgOO6FS9hZn/swevEoBqjWY32BQbk3zAiuD1FQOBV/vBEZzCKILDf+cXOosuHV1
N3ddtHq3LKv592YbDYYT0XENQgQCW6i1Wp/PbPKq2ayHbGX/1c44agbsfSgzrx2jtymFzpj6cfrU
wwmG0ZWYrXa/obFXRw3J3R5sW7NU5QUPvc/NMFhbvjh72UJxX073IQG2Yi6wa+Im8Jw3RrDD9j0x
FSlpcHJN6iuTBIEiX7Bsf+eVUw+Jmp8HzjzHpqDvmMur/wW+oKkHuJVBilmCkohimBDzez6ds/Xl
9NLncFZLhqmG9x8j8ysY0eeEPw9G1l+U0F+ypGnup89uEMymB8lbTyCgbv4w2mHrO8LGmL71sPZO
Ag+f6m/AHOJqkuDuzQzQ0TFiJRHnKC8dyS44UHLZAkeTjbD7KNj3De7ocImUZZkh2E4JOD0HGIM3
TJ3s7/uvxoSTP5pexTm/o83cYzgJR/yMz72ve6lD5l3i2vkkDj8PD2mD3bERSj/VzcnLux9mtZds
gQ+cFdYN9D0gMV8d8ucwJGQOjJplz4Y7F1sSE2adiMM19KiexBdLY+QzsGRplEmNcsxHjYcLGxMh
3dcbJxlbh1ZIMajDVSFKDzAEx1JOFw+kLvt/WcpDF2LnYkvA+OoKwnj6Y+K9YzPY3cJm/8KWWI6o
ZNpTonNq2UmhGlBP15zUr0YBk9j7PakqvbXxInmE6v+Q9sxjA12P2fxfD0C/NsS3307fZ0CTrpOl
YXeAAeIEgKHK6X25QkKJvIrGds/LHC+LpLERyX2fUXM7soi+QeK+962FekW7Jv6BMFiipUcmxM9g
ePLEzLNBlj9mEVhjfSyoBgN2pjJWDqPHG49APjYaztYWfzF/T7bOchM+w6ZZmHX9AibVhERAe8My
ykBmGuq2WQw25hOOTwcxx68vr1dQUcY87qAUb8+6gAwKvccpQbo6Xb1GVJed1vUaM4m26NOmdFFI
YZgv600aKOoDquBIqzTHRLrEZDp+zBidZ+q/E8XQVxFKMSrFqOtZWZeRaBbW48dW8+nmHpZLpaZA
CV+HtcArGeVd63XJbH8itL1QL7nCwKFcNVM5L5LK2v5Gh2GnqOHSs+KR3JprwF84RtcBCwcliJe8
rcAJHlKHum0swVe3+Yv8CT+2s5xE4eELUmE7srBNIITRdndtCsu6wA6nn/ZugZ6ekdBwtfp5ka2I
lfnAokdJkbVa5ZrSisbWPfNZKlomb9exsOsV71CzfjAwTNsMWY2xICnaYowGl7HPTnGzORIl+x4n
vNLpkC85iIaq7CnKLJ+h7qRul7NrW+XdSBoq3FgcFjWw6/9Fcr60O7mLJSPeZkIJNLop4NF1p+dg
cvC0kcfdISKUPitdo5ZDqh/n35hzAOXjtfWduNp/PO8N7oHNO9ckulgJC5oKwOe08LiQdzJGrPit
2XYuuy+R7p/6FjTczqvp0/GBaALvX1hpi3l0bq8dRtVnK0cPLKLx+u+9ddHog96rJf+g/kvKNuXm
K4mQSfv4TeDN4h2wxLgHrgZ/llnQqT10digHua/aopcMyD7QqoCkSdHvEZECapcDQH+IFVYz6ZCK
cCaxpuAHlVFR1VU/gljG05skXDdh/84brvItmIRd2mQ7pKVuspaL7N4QjK7mY3YPrzA5Qopuum9+
XVyS4kbLLwpLO8hJqguVwn3uIBIOG1ubkXtgmXfXQngss5WUS+DkLelDX7E+4cVJbPZUQkgMe+cm
+WegIlmCltD+Mq2de1NxbzfPLM3XE7CTm3+DXhZlb6rh0EHdg8BJdx8+vD/T2xv03s5tQ2dqqeGz
dH2pt1sbwIedZr6bqrmeB96faxopYMNk2O2hnxfahvlKncqzxVLMpQcbG4YYrtPvZi/NSPn0qu3d
O9r5sEmZJTUeornlH02krBwubHASKuf5CI2/gwOcw5sbVYPTEWTSz0+5RBy5OjlcgXU6y/o55VEJ
xRB+5VLj8O7d4BomNcYV8Zbouf0FYVe3z1LFi1Qq/bzJBP3hzUq/NPO2obp2TCsgxrVCVV0ywuv5
LLjNigaBzWf7R+sc3vURlPHcIbySdOpN8/kE8E9goyx/ZH31zbowvpb+xmHsOzaCgYVbUlpzg5sB
Z/qFTEuyXVAlFLpFsgLZTUsebeGvorm0RMx+t+WU8tbo+GRHNdGFrwSD8fThFbVlLn77SPPEn5WE
sIkhFs7AQa4+9ikVZOo5xXHInbNy54NuZ+TsyxEtCtamPm2TOLrxTIwWExhmowUjQMZ4c5PEP246
oTeSIKf/MTWqrSUWhb+Zcavp1apFmpYEVQ9l3PSkWeIcki1aOXZitEi67DcdYaMPx2GKzrM2Tae8
XuYsN37hEUFfC5GoJguNMqa39HWR6SWHTDmLiuqgspULauL6mkxrNvcBTLUOLSphrcSgXQSfKAXr
DOTxxREMlPGz2YEyHCyFD4DgjiUtvMpV2bVcDYa0kDe5l986Omep/JDaruZSU05jyFfPnJIF+lbx
7Mgs32z56r4Og0CR5BQVyfefgI4t1RpuEt1+nuvHNM845vTcGUgW7JGyiQCwJvDmBBp5KJmRMA3L
D90Un3vYWzYwtkjnxPRyJqPmqqaZ2iJEyhhO6Pz0AmGm1C89Htd/fDJvtd5fJxV9JLcJUeASS1r9
pYmjqBwzDaz06soj27uFMwPj2D9MMKv7NiftiQ4vALwKx/tzT9WIS37JylLBv9kaEjHUX3eVY628
4iliSaVPWqDrtUc2Cp63BEMN5epxCIrnpsyHSPzi+Y5Mx+lPeU3rSp6dON7iLnutHn59JRTEDk2K
xSwXdLzlrX6pNHNKBDZJoPn+dmesOTzXH29IN2YwTVI1HA6kfs7DyD97HWTSI9FGOfuOtYAYA5kS
hlhVuC3XntgVRKfa9dauCH2qX7Vgl/gxu/9vzyaemtU7pJmaJ1eT3uMZXrFcMBtqhcIMZPaHCNFv
hrQDtp5eJQoUsD03LXJXfvCv4t4DVv+SgKp126KdaTzYrs37Z7yWwtvUBQlL7CzVMrdYNLil0rWX
yGfwl6ms3FlKvRoI6Jg0AECLX3iP27OIPWNHNEcbOoT0o+FI5p6PVcR+o06mkHZFRGL8EVCbhX/i
YlYarn+mnb0kVwv9GisMUZS0Hq87+6IGGPjr94AgJPEgbj2+YhuzvPsFZhzz5OnmhKI45nsD5mkG
9DKwx3dqTIbNHQps3bvpOkVa76uqmUPRYHhWLXaPfW/cwYilDFSlHfkCEzn0EdSdGvGXB0pYThb+
VEfKAyFNYUNZMJw0Yr6+yhZmapuUL0OWrY8rbOgRpSw/Z95pF2ceAedxPOWEAemiiw8Q4PSajPxj
LFfqxzALe/xOhBN9lYw0mWK87ri9uHTZkzzBFisKUA5U3K+aJ/I4NMhj7NIRxtg3fIhEwcJDArcn
Za+1RSlvuyRsy6GHBrpNVjDpxH3OV8NMIetRofG8gWr/cyg6VBAEitoAyH3r4vK+aRwGiFIJ57Qg
+aNHtBR3i4Z0HQrwFgGA1jG4YTp7v8PhWqlURivVK3S78FALrZK1nhoFf2Kt2yMkCQWMQg51b9Gy
Ootlt1ABpq2hcS5Og4XbOZP6kQA6dNZZL1Gvv3fDzV8CqMBh2wPGG1BTfofHcL+nGDjtBFKs5YtY
v4kDFgh1JjDb55h2Qm0AXGF8glOheKq6e93H0mgdUFM7L59c/o0yPN1DwSJjWHztm0KSx7fVPi8f
ydMAQD7D+ARjyr+BpGkool7m37SOmB0ZO4gFyYmd0YGNGIkUEqCCq3h8rD4MUlBsszdbN7kvzM5J
8fRGXdtg3kEuTZbwU96/GHkGYA6wbBffPLl+hJ2k0nbqS5MgcJEewK3Yn8ElYnSVQiSCsOvxEZy+
9Are9YmzGxAmUA/uEfV/QyBGshK9BN0pLFh9DuFhp5T1SFdc08COgD4lDPAsNBEOqM8gaaxwB/VU
k+2EWKnGddrAc85IFEXS3Lou1Jj2Kt4VVAGWZERCuSiGA0Y6KGYaOAYlIicwU9qDV78T/jHg2V1M
Hd8StI4weLYlbfIdFg+m9Dvg58Sz1P65q36AyGbEICYz/UVUG3vQzBFpvyuedSPdUb+k25RtcMOR
WyxkjSVjRHlo8lu5EQM8/kW5GyeGu7QJvvrbm7oBgnvIBtzIji1sYADZljKEg4spffU7aU0ltubV
SO3+MuSXBKQ/MBwH//+hdLZ/DMY612PG3sVrw9n3s8euBXH7WxORyQ4kd3Wa1CZ1qca6lqrIsw2e
gK/4TnINtO4ZKqnBEYU66lKvA9IEGFIUZMNJ67bHzJia/g5kVWIlkCQDsTTfzYndQVV+xgtsn7A8
davzLFSLXYwTEGlldRTA5TREeR6nDUQt4L1JpcSa2tc3FbWHLVsGsAoTxOpfYJ6buLH1s5iTRgS1
AbJkWGx+Gzha3J1473lGz9mV6Q6qfRufO8zvbFLCp3dbuSAwNTerfhZUdU6FHyGR3uMWp3mTWh1/
naAgq+WR2I6SRYum1g+SFVs8/vCMACmYHSx/1VmkFfajWm7JM/tDi7YGibzmwaNq/iGEq51cxIVJ
AY3PVFNLonaw9EjHDjZ5NFy5eXCxE+0lPwIUw0tApVGZN8+RFOp4B6Mp7EOcpEvT/P9PJkivC06q
PAmvzqWaWuCBTl8utsRSzU9LLHpC4tdELDrEqQlZDbNp1vweyoC2Uaexk+FT16w7r7IlE9rAOgCN
C6oL1l6m/sU/4IrvP/AQmudvFu5SPNDEtzf6pgc+UMzMbZwvQlA3E1068e1amD1mPNcdwpKAddLA
lZuOH5dG/UgYi4CHkh9tYPfpWFVbTacYDhOFN2J5gW2wZ6pn+XK87sxhh2qe7Zmj2y+0AFgJ1X5v
D8ZIl909D11GzodonEVdiQ26Fw52N05mY7uuhQORvaq7/4+GKtSucKunLJQkPKDDu0uaCnQoAZbw
IRWb53Yn2E4K5X8SBJ8R3uiHP0OdW3YGbWEMb/zi8Vq/KSx7MpJXHDM4GM2HSnNGvUoHH3A+HKek
yDBrBJ1KRn40viu2DRXmiA+eKm+/2I5QJ5Ge8F9cGjkLOjn/5AUzUvWfShQYrJ2Sd6MVeCe1vw/F
6CGtC/fS1DJa/0sf5+Nd3o0R+OsIUgcSPHVzbRJAfGkuS/3kPdpLLRMZ+YA4eeVEP+21a6XbReuj
lyvRJegjV+NJoxcTB/i+sOpw4HxtCrC+kFcRFGIRSG+ONnlBe0X2ZEYCdgzw+bgMlsUvH7RNRQkV
CypNhTtJOJvuc8PwyB8CozQmGPoM+7T2DdOzl7fadKopY6RuPF3tewDNGY2oxP7k2vEmUojuryvE
IN75/EzbsIVGzMilOmpzys0SdHabYLWTLWfTpOHlsYYAu4ceB6BvyBuzy1VPwlwEq0QMtTYKokzI
tCGljzH9tC6njYGVAmafRJ1PBMC7exne5cKRnbGkzwO09K4p9XJgqcQuY+m/UF++ajYRPr5iTt57
IC1/3d1kDoFXWo189UjZ18ISz0wHwkidU4RRqlyKckWWt3H6QHSxanOlpuLKi6LRwiLhGlNta/A3
zK7nJI9mbB60QY7qciYLhyPn9yBr4IBbOijbmI7fvLoGWnzi3EAPrqoAHKqui2TjWAw3noYHyaZ2
sBWCvMPsCKl7BP0ZCTo8qN6fuGiyQ8uqYEHYeTgg0m6tDj0Gq8pWKWk45g83y4ewUc/+l0c4OXVX
iajZJjGzSuaF/3migxMHoMRdVi1plB800Y9Y9emcV3iEhYZoZO2Gv7Z5mJuAeR/2M05Iqx1fs4Tf
t8sBpqUWJ5MngQBc1F84EvSXaYs7jhmA23YilCNK8ftor1NlNLjlSIntmitc+p9BEItB5Jj4BcL7
Xyade8fFrp28Fyi3lEYzLpJbQN0jLaf1cKYO77qjA9cXztFHAq06IXfwdi7NF1nIPQNrRZh9iLHt
9FIJAgJ9DSL6/Jelkg3uQRlldWbjT6pEBcbMzTpwJC+qSPZlbLH8y8sp2iKl3+diOpC5sbBxusiH
V3Ve8yHCxeNfaw9NJ2+IJ9Av8ymJYMd+lQ3Z1eNhCMzh1RlrQXMBt6fAJwGgN0ZRH8w0igjU51Xz
MfkajX/2ERXzvjXjtjg6OlPW3voUyH3Jge6XuWJ8nWl6s47efxKes26dB9T7CxkqI1Z46Zpe5ZXN
NMdYCU/jUXg7v5ie8f3rjvUUy1h5vrnvtZZW6lz1zZViE43mBgNEo1VgmDwKoZS5kn9GRPE2GXf0
ZTnzvR3FtMwBeKh7ODk4sVHZgtjVv/xqvKG7qnuu74sM3Wq0RA4Lj7FDNDfer+4jrnzoJYBdD9Kw
7B/puyM8mSE+Tm5DN4lLT66uy3KVGD3PvshNiISLJ1/hnlWm+whCDEps10WvQ4i2/vn8F93kZ3Zj
YvRVV58mF2OL9WqltVFcgiFVJ+wgaNtZNDNKXiwaCdlpRl277pHUUxdC7sYcgMQMk0wx4oXuahX9
4UnXniTS1VhljaQZ3aAbOJcPgunGLYq/gBy4l+kULqINqzW91hqIKtRLabS6TGWtoGTyFhRP3bmV
oaJqGgl0zwUZTjmgKigaSmuwcUYyHFocJCNwATyup6JJQ6I3KW7Reqvq82ubC0FV98r+x03d+HWE
C4fp4O7UwFofpEHMa2MIQ1cedKtcdye+693laV156mTsXazXZ05EUOGHlcYKHdc39rt4yHcTkX1V
XIuEEyoDqEmq5YuQWeoHI7q6aZ8+/UsfXlr2wf2YM5HuhkNwUgjaCiRYsQotj+R4EnHWYWYoJDgf
OEjRQWsQkhIF8l+Ziif7IcyT+BvJ5aQ7OhmMt+zDyOvLtVj1QUBr8q5r9UoIrV8l2tQNlvCCwl+s
JLDwAiVkJMrg/Xxd9lNqaKO0us+hmTO/WyURheiq55GPzs4A82oTHS7x1Rb2qGkh7ZtHDLeRDzNu
FH7ujOSpyUjLssKoHaZyM92Yz6VwcKkITxKApu/3G9JRVW1Zih5dJwKW3/+OxxblS7qiVDoxtF5m
tresx9URpvljNS5f+IMi73FWsJCPmUnSe6YjUrdk+QpLydcE2C5zd/6SFMz9oXXF1ezC+XV132+X
aYts9OplWFT1vSbHCR904afKd1yoM7OT0kkOhmVMdxymH+nBc2noXiEXAesi02fiFSmCBkEUa6ih
hU0EO5swwSkIGaTw48WdlCDcn5+DxbHRYLgpC/SvXDjipUntx+dfb2g7NUMbwOehGhegzyGwWbpU
MIVmUKqmOqqdBxuiZF+wCCrWq/vF1GmgZF+bf4d+ed4lAL1VoD7mDE24HTWl49wStBoDsfN8dciR
qThD+XAJFVM0oyMNwQOuCMDWKFFchXk2v3Ce/UhThBPimYZ3DFs//iAPLYi1iLDqgE1PEgUdQoN1
qi8uOgUPgqXGli/LFOX27/e39fOK/QYiNAWVNNfRvU7P3gvdEWuD3ZL9qtyfL/iFMNJJjpAkDeCh
imCsqP3ns9kCIdWIp2dancGVaCHNy/xh8NC7cqHEh8YsmRCsEIqfyhn9vR6Uj93fhuRmWlc1xb6C
GFxDyvm3kNqGOW/R+ljtnr79LnCtzGUWs45IzCzhPgKvldLwZx2H8SnCYJ3jgt+QrCw790WB6oPl
cQJzj2EatUyvbxlazJ790n8gNKPQrH+WvN3XCI8kf1lNZ8i1QRFedFxRrOufb665DDQyZ8AvGciC
VoWP9Hv7iIYyiRmCZvZtnXZ98h+9m8/zoPfbk7XPuSOAzxwfhway4Fe1/o98NqBgjoelTHEKzkVn
1YFhp5/ZufZ/lcMEphOkMVT54z9/+Pp7MpCHsNA1KwXe9qUJsWsbQJZilD279BMIbBuqCNSCZIOU
aB4Wo2sQoMxBMPvEp2J9KRbKvx8zmFwTvEABfneKAd1g3cTwzUL2dTOuLQExE2qpaK/hjR12DwOA
JiiT0wj0JqfdsiORhqIWSX+1UnVti6GGhSLa5bhyJmVdj0j5HOxdqJRJsgTCfIjnXOgqoietxwxs
YCK+/QXDJE/4xnFVyA9mUiUrlh90uShLaeJtdduU4IQwgIRGGEJrklZZJghVhXEYTc49hAMSppdM
6fCkchQwN8QgBFGcFsC+nedhSAOzVraHcOYyrekMS5f+mvSAKpMCIalvzVwSwz1QPKqjWhoaZGf0
t6FSWp8lRWITD/tNDN80tdN5kTJuemT3LGu0YuIMTyKs/JiRRDp016vnOXcmdT9paCK/xYVQjNfE
Ra86SgoytuXZKBFFL+6H3fis7aM0Fb9Bn88XMwQxyfzX88yxPvIwmFFYYwpbFpEQZQflQhk8xUmi
YtzNUj2ZojmVWpWNsCXDeU9TZy6jtW0/H6ci5mh6ep/b+HyssFDg0Y3lgeg52xKt0UqIlrCgQLXR
HBvuGRmDiLrZLs+R3dergjNRw0n/p2FeaSxEN9dWb/OfogHwgUgf7PpJwfrKH+jb5XIVJ2rMXA4u
UmeOPVG33OhK0SIVD2XqdcGMcdETmN7nbDNXfxxvne0FOyUR57CYbuvbMtUzoBS65BzlXfw64mKJ
mlfJAEUarBxBlAofGztfa4Bqvry9KcX258GxGMroB7Hbqzbe6mkieeamY1c2Pj1C/aKrvPkgfSpx
JGfl4zjoHdlzgiDZxbzBzpnTqVVZpieCm/x25EyCzRdo0hKhT2QTXKef3D7duUrd2Pel8aR9MXvB
XaKFql4SpGTS61SwTgZHO7jxn5Ax6rNljzqWvJAPh/F8sRrJtPj59IORj2C2EveFJaP4EfixzeYm
vpWdJuwGg9xg1xwDPt8U/GKWaBMfDXu4Bc6EQx1PUbzQq6SCNGELiH0+gWXsMM4OLnkMIafbpc0e
0CTwaZF2nmq7xZ845ba5wPzM5GDF2IlYC2D2TN0kyY+y0zTsJGLzGx/7BiUQKN0aoJwGQM3lzRF0
jxTgGVyhYv5WZ29nxlRa9AQLz3vuffDpzoH1ehD5N7f/CF/JiQrpjmnC9eW45L0eMNzZQahudJWc
ZBEmYGHYOKlhfhwD4KemseusX2QkqxM7OrvU25/VEXoXr0l9QH2HkeKevrxUIMHW7jmLiLXkaRFi
0vxhMXZ8ul0i1uOYE7Enp8Ucp1QCWH+2q/j5iNxIUJS6dat19lYTK9PpJ7N+yGTas8Jaj4/pREtk
aUKC86H9ZHJAqJ/244uDPcplmWOLjVGa+Sf7VqpjkvBu5La/vW2LiIeAac2QGnj5K1OyFbTgAZO3
Ya+Uv8Sya3caCsvNdszUJn5BN4mD+9sYn3gSYdp0PzCD8dx3rwCWgphB2oDqXwynBNAbLgS+daxH
FO0XQ2glucqJs8cUiPJrX+r9TaIHFbEgxrQA1iOU/uas9DHzcorl8wSxbi4EQXBBAIqJjX29eXar
deyo0dY8WSqcIElsY5XjUZD0Gi+voSb6ZCr7jk+WXp6W6wYit4U9tTLeEOJBGU9tjHfKapRGm2BM
2Qk8aBGGRWXsmpv3qtCBctIXwW/Tzeg56olvj06hUonrOdWW9N1QAmXZ4Le/TQzIrQOXl/46CZtb
F9rLCd8T3YTrpa2vI+14kE4NzxK/du44+/1VYO8Nsx4mkMEKyM8SX6UNNw5LujH4BrTGR5ce3Phy
vKM9Kw1qBQXLry0+i0Zsa8Gi8UepqAws4TmSKZRENZgRgf1eHfF861LZTkJ9slrLuMf912X2d8Mx
71bBYe53BYiyt58PbXr38+LQ5kVxvPpYLgcNaeyKtmG4k4fNzhBihIcWDEaqeOMi8gWSpLwPEjPR
lvdIFvNF+aWoJbEi4jX+qiH7bV8Jsx4N/fzWJ3F/odgSDMvPD2/tvyvrJJrFgdBbjdArd49ofi7E
pP/e9og2UpNIS82andGFw3cueTeexrn/x50lxTmHbHNfFvws3iZMx9DxRDE1rVdAZ7IUwVslLpzH
EpS5ykk/ACoHlMa1LUPtuvx9XGf2cWpEE7coSD3tUZd440X5xjpqN5Z05+uTlDzbVPS8bcl1tpf7
5+UWlViI5Kpz6L5t9Y3jGfEW58DDqI3RUw19NTcgMlW7MQWDtdnNmMpVJWam3/zJussbV0/0qeOb
/9ITEKYx02zOF3VsVNGXddNQhmV2GcojbJ4/v+uiPtd0iXWvvuf431c7IQEUjCOAudFiZUr6cIcs
axU2HupfQ8d1tKsxX/630tX/yu7qeMdWTaC6O6hDwXzqt/d3YeO1D1qCnJrROnr/gMHh74K0Y5Wc
H0jtqj8bnkyKlUxLKZh1JSWWCGtrYlCFA/WGmACukoe3DQuGEZBQ0mnQGtPsOWex+oJIYZ/MeEXV
mLXwhmo8ie6v81GvVEkhvmzV/bcTdr7qyAg1+UHob9b8wWu/eaphDDfryZwY+MO4YHoRMnzXhosr
YuvbYMJ8AVkNe1nELOkKI2vT4Fdseo8NCL3PT2PrtNip5zx4o72INpOgmSpb4IvaBSboaFE1CvyK
hfHF58dND7wgvhUEFEgKfUzlgnMVXhXqbyGGQ+NhVao+jJS+uIPXYIcQI16ookPMSWE1gavp25NY
DJKXxlmRmWnkoyTZ+WNiEOP7xZi3LcqeTW/aA+am/Gp8ArW8HonANIZ8Hm3EJWFBXSzzYLWzzqJ5
pJ9q9igjq+529HKvmr1uYn8kfCYeUrcQNCXQ9/QBDD1m2Y5Gkr3b2U2ae4v/utp8CnETa5CtUx1k
RK6v4bZZOI95YDmcS7zLVj5iGWDjOxpJ6wxtROLGUU4Zh1M3VIqkesOGHWC+bjtpmpUR8xL32pbE
5KXoRYOK1CoxqBmD2c5S715PLKWkCizo6BdqTxeoS154xONH3birvyG0NNCeXaQRsNorQxwahEZI
XlTh+ij5SyMOcaTUeUNdTKCzWWEr6qtbRkEWkBgj4giMKX3cy/B6aYFckI6db/R/ELVV/OeJiDMf
PqpunZxqWzrh1GjH2EpRq7hmboFiHPwGLmjplOx+AJaaQVtrQRCAb9rduRoEYdQ4ptAXZgLhahQ9
rIJ35qXbT4FfAK0NI4iFAFcW6m927ymR820Fjl22LNRJ8FLFUzrhR6nUdH+EAqYFPfH+aSAOJs1V
va5G+expLlHmBfdU0yNv5HdHMWlamMS6apLw27MF6XtUWN7fqPe2Dng11b69RtJxtI0KWsycdrdr
tP7hA/EY/lu8eAvfzOTmIwK5O/NbAgucQBAepFNEjnTytcxEkaIbmDCMdWbgOCP/t3R4+O7ySj0D
BDis4oa6oO9FDDGCBAb2lo2XeOrSlREUEtX0vPmpyhJF1Fy9yncjFieZ1KpUXYu4IQGX0pWWP9BL
giNPdAMNQcX5CPZu4uEAnhNV+Mx8rMFOyi+veFBrh37h1I1/vvuBj2yKPapzSWX3WFGkM6cKmJuo
eEm5HN5tzrm+yUauLAbKcTpMCQOESlGNiBRZALx/yy0j1XGxEVsVuLsuvpVgGn19jfjreA20K2jP
1xpLxY9GMlIlOTWNDJ18ntqMnliR2GG6CunjYGQKhnWQBR0uo8cSnwnzhd9SRQb37iu5464y/0z4
JC0Z07zuqszwmYsRsf20cTctG+rcB+vcVw4jPlX8yOCrWThtGCAHxdspIfRMghuGXHMmHToA+Dhu
CKt7EfKSEe+UG/AOVnDbiYNam8qKQ6lTGOBkZTUIdUiD/N2YMKHBb8r0GFtW/eo7tuSTNFifGRxH
3QuRx8ZjO3Wmvlu5VHo48K/NCZENuXs8twss+1NRkVK+HktvdASjbM6iot8+icwZal9PddHkC3SK
BJykVBaNGXjoMHeNBRyLWIB4Ek9sFmcDEKG0MAC/6hOb44EAWrQAeYrY9yyp0mCV1N8cij/piyKk
0bcwwj1dLMoJABIuGQHLrlCqeSzF9nRMATqxzFGULaEW6vC6b5MvZ1cFkKRoSQRZ61vZjrc0TqVq
YnNNl0jWLjW7zOP1AYy9wKtteo5zKHUSURQVIYNHEgPLTNU6lO8/uymaqQHQdVA4qYNvo8TylgJ2
8aGxiX4r9dM/7dh+TpvtXgBYkHn+ymDnzlmkkiDS/OhIeAqP3eD2GrSxPeHPhXNCOV4exJaac8x7
oyqsXxQgnKKaUj1l6gPvq8PiLJ9dQ/mQhM5AnKoup7+nOTGww8uicp1peUnvEB6GVC9xiVPn/Wk+
fbO1l7Pvcjfsw5zzzwU3rqLJJ9OuXQ/u+B1S6/uianHnLFPaM3BDDzjs/i3KmUDca65UkLde/+rG
X4S00dWjaA34/dNZFsUuFst2agrX6poxNp98RiCk7q030Dx4JG+5jRC5c+IzJr4aCoWANncXcORF
OOkiSa0XjkVIp8JcxcGcdZpKeNeKqA8h+un3PJRdsJhcGjYHoddZQS6JlY5Qtf1X8BO93hq3nSuR
jnXmzonrEZAHWIjUbTpewq75tq6Et4zai4m6+I0iwteh4iqgBe3qWSI9bW69EtDYovoyPks2hTNP
CcRDNBAgpnEz6dX2q0kykQNg0Ggzs8KDR/X3GdQ5CVtJsowRdcDjo5K34YMZhlIg4uy6Ei4BVUqa
/RJpOQs2spXSZC6Ak2FtMZhFA2QC3QqjVyXlNdyG2pMd2kV0xGQvAZujhTslMIWnmSOeoNDEEVs3
aT8vk+bzp3zc1X0Fp2TccCdhwkrWWjB03BpY3jqw9/J4uGguFalfQWxtZt1aMUjTolaIKiuImiDO
Wcw2GDDbVadc+yh24BBnirPqw7hLu9dW8blqLcWfmlJHu5VFrUKksoMANn1ilnh04652P39kodS1
qNWtdNt9/3vXQZqTExu7ZfaCcl+r2ed3aKoa8whLBqWuMuyEyxvmYL0GKOdl5PbRLhqiIrTDAuTk
ofjV1eh5Alo2L6AE9tEDv9YeABdxkZ1OL5XxktE9d4i4of20KDbH2NhEZtFuFCzVWcdJS24QX0EB
Kb3KyCDDXPx87V05aSgzFuWQQCLSgRqu/9Cw2VqPSFTSUJ9QKwKtN43QMeYs/x95YoKKg2lCEoq8
Lk//yp1ToxCjwfX8hcuGNIYYwbCSVPjPOMm3kvcTvk1olxxeubH0sBq/63ngvsvyU7vzdYgziQYZ
/uv+DvIfe+oyL+86q+tEjuXPHsp1ar256ywPq5eetjuGGt08VB6pCCZPJmf6D5PlrLsVIKzmkHfX
paLc0Af2ZiGFV1OobvH5BYXDn8MnJauUygSTKfRQkflMQ0CzqikTFN5+/jm+yQHmv2fs9Jlbcu+H
VmHdtbXkUGqtmdfS8auH/1W3WcSxLxtw3yPGdCRSFX9vM8clXsw0xXolDcerxLzBR8LAxRp6ahnv
sqLjlD4iVq3hOlG97K5p/6vMNQC3j/3XzwtpHHoUJMMi0lGa4/eBNtRI5oXU5GAcRuhBWuCM6Rr9
mQhTBCQ95lDPkDbgQXAfnknvTiienlNemGW/1XaX/P9621e4CO9D+Nr1t2WfzfEOmTO8p7VAoEPG
c7Jqi+EGMfAyv20DOHtXBkp5bx3bavYjTYifa/TvQXtq6BctHdbolELvc3ZUkp2OtkZmudg5sEmQ
wRGT++4cL6A/4ftOVaKOr1vig7Jt15zmo3Gc/tPOwrVDT4VP3V3MRFKSk9ZAa9h6iqpFL6s1gENn
J2o+6rU188u+sU6MpsDNOqB/s7w6IITxVFEXygjc8Vd7rSHZRfnbnu7ZgzR5qnw6ACk1Ofd1NZp0
KfwLKy/4JMiBjT4BAM7xyD7fm5Rlgf4dhkL8KwuRQg+nrgadL/KtH2JADhlofxd9JfOeP4ft+3K1
VBaMz0Fbu3XZ77LGy0hOmX5JhaPN4GbKLtT7bAFcOGxTRgFi0MMLg2eQ43KK2rsxUsaJuxPWufRm
N7q5i2KElX6WCHCASxwtCVlyhMzy+Pf7uvcuhCFYixW0RcNk0pl+VzFk98hjA6lQ6osxx7go1otq
0DCLl5J6koGNeer4q6MfOwOTH5wT+ieNNqp7m0eGmtRiktHYmfVdjE67Scp3ljIfl8jYqi+Sb1Au
K8QY4+6g06iZOgMiq6CPaqfiJ9wcRqOjPq6jsTr6MjbcIcSHDfl/0TjQUXAgWA7Djhw8uOLsgUbk
NufCqVNe05PQl6JFflwxUvS9rRxdSe3856G8JKgUQZeOfwCWxg0hAqS1jAHzxguy0WcTe8O7a9JB
aVxk8xZXiG5xJzgKcvGrCal79jSVwsy7s1PPk/qd7sl8QsmFhsRntsgMPmjVbZIp4uDb3Blj08m9
JppFK423GkPp9w46G3P2Ig1b9nwb/ytMKC/j0/McKI67y4PbFrSrBs42OhEGEWPzsH4lETt9CbTp
UB3hd73VLV77l7ehTvs6/srHjgoxNfNj4Jieo38qsYlDjUr2tDbAfigFTCjCXaHRwdJGa5omIXo/
jCec3urGPFo24eLcW1JdV/nUNhvoYAWMw5RgsP0FqborM051orsHAC/KvJgAgC9nQ2EZ5ZAAsYL2
pFdhRiVfypcIOxl4D9CKLy7YKtbKBppn7i+F6a0vh7iyhqS2vTDWgtbk/+Xct+sV3Pqfjtz6hJEb
pVFIuqgYu0dA9LxsUy4aI43vIY2d9F0ZBe4H9ulvq7KySVwg8Mm1O9O6Q2iw+tNmWCx5o/1nGW5d
djdWazRGPMORdzyaFAgcZy1k8P0NCb8qz9wh4Tu5IFDwJB0g6VjFfEqKS8ziUbG5Bh0ivRZ0wdRA
ZflPDiKWEDDMN9yoaYzZPvkg1/0gx9L6zpBgGpIA+Nz0xAveGgtt50XpbN0dc/mihsX6fjF64kPt
bnzUhVAs2SMZFjLCegFtTOGbzxNW/MkXLaKVS58/OjSHtUJqxjiR0smmcmDb4cahBK0484WVc1t4
hIwWBLpw1TSorJYgXbDEYsSuWl2dJH1sXfifcIFF3K82cHH6h05zfQu2ydgb9xBMVmR22/XpsMXn
Mbdwl5fFUB5BZZlbqCm4Tk6VQAtZgIOIkIMbXe2dvaIzTw7ewTib4oLUTr3tzuUETTrk1m/K6BYn
ihAcg1vAv2lT8NBKdrelI/YK8E0O0kQwdQORwfUYTgfmueaDtQIpg2Tn1/rt/nABRwiKvntENQvD
Vu2HMBkpwf1lPbmuaIH7/BGuojZ9PAWgi81hFrbwgaXP6AhU63IyhRoYEcQ+sQ9qV3Tb43B7yFrX
nZs9plbeo5WuOqo36rNT26XJ5ShJVCu4TDdXt7j4+8ABoYEEc5hcxS8MHCwC7yk9tOT0flyle6en
8PmUV/Lpr7nblyuxIh/frxcP9UAlG4jZslE8fXYS3H9knREtLGxisp6rd4t2AEHFTKaoFLZysf6K
oIIACneXaetuRO40lfmp/mpxfdKHRigOh9qeEmSj4cxKwsEmN3rAhGNe23uOzBeFWON0t8s21hup
FEkKkPom53Ht8O7QgX20eH3GM0GsJZkCRlZ28CoqM7zfgnVCH8GOrntWOGONY2VyWKwJtAU9C1f9
zSdI6sLc03XkDw9HMiZ8RmyFZF3Kt5j3bJFW8Rx2L6Zv1aM1pFodu+BNebeSEJ5an3RX0isLDlNj
qxErPvCM0cJIAVcGjmHhzDpQmYP2pYmvWIfLW2DY+KpvCnA431WRG8ujOLN/OlLjuWovMoJkCJxy
k0MWHJC9H9fDZ4bcz/kn+6I12Le4OxL1NxudianTMx26/a7omJnb4kpXQtDK03EZniXFxdsAS25e
w22kfCB+6S9s9FRAWkwMDMo1veCRoNDptev8RMWq+sxJ1siRJN4ABFMkHfCGpGpwIgAPQD3jZnb6
KgYKAou9JZnvfFsCAiaU0P+UoB5De740Ui5TQ25JCgnuYatU4eycWt2wx5dSfNy6QtmYTi+1swBR
h2gDHHCD6iuEeYmC76uGgxgS+Zgca5K8fPa2qvpfKX0jgqF2+ZKL2Nyx5nVIFEE/wMOR4aaFYI9C
RWxqS4J0jzB560ssfJ9bwXo0DCgOyVHacUZf+7oQYgbr5n0vnRiT+UJXsAG1raCKwg3yhIbQxDfh
jLFlskGoYaL7DkbxzeoRAa701Bc9/t5I0tvUEHhhqOFmnJ+MlA+KxtzV9JGF1trrttHMrEKfRZc/
hxXTUliCHjECKvPrcoHNxN4U138Ir57sua+mkZ7688GmgLf2r66QFNO8Odb4UxmPPPj5wFJErNDt
ry6qXtfTWosmHudgrBwWtmH4wmvsFypnJcqF81pJP5pnDJy3BweHLC/ZogwJLbkXxV+p7SPvKrgz
LxEaaQsswZJNZp9PjSBSThaemwX24XHzlJo1oMvTjRh8Hrl48kAFtYJNTYqLuaxZa3KU/FdHTn2D
YH9fUJA9eVq2Uc9GsU+67eFo/zR7CjCiXmhKAbcJzqzgXth6Zlj+rNQ2wScyC9GycV1S20C5uCZ7
i1ioTGvH4XPQ4hfzrFj8ifSSgDpT19THYj44yW+ZQmnKjc0AslgFJ+cm1+SmbOgXIWY8xYoHvliO
AyaKECQ31od6Jcnuq+fUiDqmgZV4FLcVa+Nr/2d1I2nRG5ed/ZiwP6sB49iJ7BQhzQvPbFIricYu
t+w2N4E0ULjficx9pI+fzFoSbK7knUKGX8gn/BhPRzTCkNZMnIIM7HoRmINmIjTTQkbJarGZNv7M
5wtkBb5yQIbySjOpXnLbdAmkgw7Iywgqa7Nfo+w8Qa+Pfz+3DvmIy5gjzMXjF6wZu3ydkFvkpNOh
oDdG+a0xkd13683WZSYVWJvK+g8UmPqKKprGlJlXo5WA3rMFXpUeASXupD5EkUrMACpDwfauvDP6
hTtTRSvxpjmJ0sUi73gPjerQ5B1NzvgtbcXgWGcpemkpzrJXzaaTkaNrxsHDg+RJzS2AwbWrYJ2U
+d0zYVAALLM26hDMaoQYElXqykh8uOKvjFcoUsJCV0GyRZlWZmCY0rH1fgp8IfJbnjRee/IaUCuI
u4V9ovE5dA/KkwycSR4H9Rh+5pzjKcxcBdqEWqwvp+SniwNeASvL7PwVjSLrCe5WEh/jsRmyWTAi
iOoiB0qL8THJcqMY84O5SdWOqwQ7Ie29QP1qXHJjMkr2UUA1S0bs+Hurk1vOSLkIIrIC+1MpuBnz
/GKkrn+X7a/3C1GLS2JxsYR5cl7eI9pSlGKuUsZQ9LiAQi5Nve/LvKahZ3KctdgpKC71ue+WIlXc
+NsvfDzw5Rycj1LXqkXGXmnbMIkQhQDvBtyqPVgJeP0cwTizACIKvsfWRw/FvCzI2yZcvEK6DHkH
pc9yrECRkip5s+CQHQ5vnRqnoGA1RqNIRYP5sRnj4kX84WhVrFjVTLuSCiyLQlvf/78/oDtROjYG
LsDALreUIBmNwnGEBgadeNdC0HzCJJsccG/1NIq36dPmY5VEuky2SMm0eqmgzjXjUEFrSeS6yUK3
7nUeCszZuZxVqPdhDoevA58eWdCIpqyDA0fmJBTdJ5bQMVKU4M2naux4J4ZxdolG/MSmP4unXUzg
l4e89mTmDmQMyLCjwH66YacdVv36c4MZ8yz/iA6Z8XTWwwmG1xPjZehWsVe7AV1LCs1/Miq1Zi1O
fMT5vjGPKLn4K2NNjxyh4I7reHF4ijC585cFB/Mlay98hpRZ3E5InmMaGyiM7U3Nfhx8VzKaS/iY
PIE5Ysz2oopHlw5sYV8+ILGzOqYGBMa64tDcr6ALlgarnv+rk5y6bCrInj5F9l/TEGCs3dJMOguL
+wk/yTrGrsYQ+kVSTOOe+7GGEK/f1hZ8z6ooAERjsEpwYBhJcLqiy9fKbxS1X+wWz671knuVgsYc
rx7RwIJUBiQ7K4kKlPGO2Bc/T/+hoENOrt+aPcNePTYII6qroVwpvaOQMMYaycJmLAmRikP92+4z
ycUmKIhc8zaUcVRHXbcujJN2YXU2lXA+xXzl5Etl3/RGKC0Ci0Ec2OcEzsR4RGJYFXgX3jLUZ5N+
ql/XiVQO40t+t+cSjsqT6hrolGtgRBwDELGyNJNgkhglxS13sS3orEKu8ThaIZm+iEy48HTvK2Dx
TsDs56mOg2VrPdoeByZMQtjzuuRlxsym9bdw4Nkcv6nk8YZ3tvpIIVL1EtS0cnTE2LgxybC9SWUS
bTBarGtc2rMyXJ4WTKTcIPCbINWy+RYUYYcxmwN9s13suX82XISNu5YPrgfqf3/7DJX+0EFTcT4E
Olz2TpSX9z0OUHXEGBJvMAd3jlJLPbfuR9Kx2Gj/tcJEQffA5/Cp8SRrbjhOaNkhznPXHVG9zr8u
rwisebtvKyz+EItMorE9ETWHqsvdbcNR8bdqpGq4JWGUUlYV8pjVdlqS0bhaAqQJinjvJoPurvrY
CWsIn08/vQNWJxvaH/3W5t/ww/vyurzsHGTy0JCifIMADMKm0QYbe97Ax0pc+2icFmn2QqRzI0G0
/rehaKnpzH9LJnFeyniqtvxExbAJxbW0GKeyVXrc8BG0M5Tmolq1MqojAnKx0FH9URMmwmhjOqWm
1exb8SY5hRZLpiExiNfgrgh+ewWQqT7DIICBzKB3D4+n3msX3OSobBhoLQxC7Ri3/j+AQMgCndT+
rSUGyq3qxz8q8rgplK2YriadV45BQyK/jd2mKKlEQ9qfgWQwb3pAJ+1bR47FUrXUiVovEVanqeEc
P8zs1y8ZDbgvIJ4fzQY/4lHfD+3B4l3Q1/PkboLbJNMoTGQZ4ww5xbYX8bUKb8eqSGFxJtnW+4O8
kyNuyG6RckkohIwa6Inbx5Q9HxZzRxDi+U81YiuqLXwzPCfD5QJPU1188+Rrl73cikN0jY2XFMJQ
1IHVj1/r2PEwlOyrRqjkZPLvSuM2diMOvZ3+66LWaQ3LalOl6vT23AE1IetpqPFK9l0wpqlUCFHO
n/6tiP3/GgNVOmEm4up0AY+MaSKFrLnxrkMIx25t+O6fArhGC97xLkGIDG23EKga+9x5UthQmbht
5QiHAVZ2WRZ3vNcoebtwf9wiY8jyX7m22akqOBD8kxSxaE4oxVzFTeVz1v6CqEHQF6ql+cUf1PhK
VDiGneX5F/HjcdbpfIPF0/e1g9ZZIVxOJknAoopiriwCr6oTbuMY8T8MFMLYWuWWIlYnJSb2PuV8
rulG5ya0HNaqGv6DHMopND226Amdz6uiwRyI2ufOfe+BK1/hIXkQreADejgWm0JHStwlDPtDO/mi
iFqTqGCNlJdpprxgPgnoSrfF2XK1zUWhEGfbm3j9IIC3iYzgELMCeSwtgUfJ3nB+68aV8r6F8vO3
cIf98LwZy/8iCbS7zBWrNQ728AuI3DhyscfB+AaT4T43ZZ5+ZMr0x+/DU7qfIgXhBiW9Tx5azUQw
PmbH9cgUUhB3DJAydk25wa9C9lkxEIC2oi+mqNsQfm2Az7f/8P1LPP/WKrjTNHaXxLyGcqIUoaVX
ohpHGjerds8DmgXYI7WCnDpqyQB/xvXlJwI1Tf2fm2U1U+x4rh5f03g8SYl3PIJP75EdB4EZNjvk
V6JweRFkuxTX0tWWmn5KjX2eYXCV8eV0cBC4e0khXgqVUm8a2PmFD6mjH+0bNPj18cmtelTiMtTa
cmbinN6WgCEHI0DX4psRGWWoEhwh8sqEQLu9ciWcCFYIXWZo82peGKl4gNnxKH+rlH5xu+Y4lej1
lkN128zxP7GPnQpnD52hyb4ekdv6yJJ0v4zuMxckuADJLiVt3Bk81myBcsV0LnGTAGjIDHi21HXt
vyy4o9iqVlukIFmSXwNYoG6JXW7RtGQA0Qcgm7FdO8U4IQ3B2/AJJxOiqVslTZ4eLI4yED3ozE4j
N/l+OtkkuRecdD3CT0dU+/hkhIDMjYxwYjPD6E+/g4eFUnADC9k9Yp1n+famgD16kjmYJ7CLbQYu
g0dvVi6zqbC0KljVCeScmFLisqqQ2R4ERyE6b3A3gnKeVh5N5YOCLLd9d4KI8qjjJY/tpVtFy2cK
F7uCk0DLRS28e37XWDrNSKVtqkFsSZBdWcgMzZmuKaT9OGHin377znk+x2Szf0I4mHzGTnXl9aVU
iUgOCH6BkBTfl6SjVmfOmn2UpLO/TxE86LCZcfNxlVttxksCehrwMeTe92LNQqrIbIBf/qVD7EdJ
cO7YwrMyw3364yAuUKmGr/b9mVVJAumltiUEXrwk8IxSwlegUfuQfUNoqXnJyjNyI996l0g28qE0
Djk4UFmBMQ0Q3LkfXAOkj9/nK4UOFQxiNbpeoFMp8GwrqS5rUPRb4nmji6z1Dofkdk8TllfDFgmi
uJA4XwAH9VU/9DvcesURUyofOgO2eXf90XDqocPqUg/nd7BXMXCxryeXLx/0fmHCoarrd4Xb3lJ7
9ZBRL4a9YnRcz4VS1fxOuvxIxogEl8O3/jP3YU1KgOzaB3rPoAhP+0/nMdr3DOIEZW4OV2afvBOL
srng8OI0Q9VzCm4qVVOY8PPRwpYVoB0huWSgblThZ8jnuj3x4sw+CMHKqnWK++sf2ltLdyRDdp98
cHELUa9MQZm2pKCCoe6PZO9ScuLcupYwLzCdanbMYZpQDMR49ak2hYpKwV7nDdfLPgralf4DXJYN
RBZ4gapfCN4QLv7ZgeSO8Yi15zyHnFcfDnSWhNhvQXdpedYBh8sITLxe3a2FL0NfVIIm0r6fkmpg
axYMMQKT41cNMEaAYQsdiBXUYWFe4PAAutrQIAEix46559Dywzr5TKtf/TIpFZQTNfU/BGavaeBj
+Mjzggk6tMubeJfV0FPa9zRtO/mgmpx2Sfm1dPXSJYbfpwuHQPXM2H+dcTD/Z9sZ8K+zS5bBhaT1
uQYyboa5xpgSU9TAVMKR1xnED1d2i9xZupeZOLXpR+F8dUrxDDSV4CcHVYm9xZfYWIf9q/OaBuR+
Ql+g6bbTSBIqagkMsTTlIaGIxdc3ZzavZ+Yh842HRkXxArMdXkec/M19kbK+B1bSe/QWDq+mBPs9
QaDSujltnXz6nsAekLD4/HLfQPSwO24EV0m5ZROY8A/lm4ZpKiZjMVOAK8OIy6Ylw7WwfjMuzHzx
qLFK5uZAKjUjmVdFFS2Oq5SvjnB0serkCDO/vkttJOefX1TDQjg0YIGNe2zO9u1deeaAeCNwY0JB
DdJJqEj+Nwt4Q5xSJ6BMlZl6rGS44JTuEpX8jAJ4o1ttm4vV4qSM8Ey3qkgvcQoP4LtitKPiBhyf
FTut4XCBcaIylUr9I33tcSkUKlalKEBONqz9WY4DIZ27oyAAV/qHTpNsHM/zuAzKyxSOfzpAQ+Nz
Jzd1so1KiwZYN9g8WZu/U0cJgRjc8j6Z4BvrPSRZt0f0/8YROlRYrSYiWHpuQaTjrie5jSIYIhwC
yNbhd2j5EswYOljykhv23HBSpyLNzPUS4QXlXUGeklqp+FFg3GQkbjZls6laGgBBz91PpEuSSCtT
1sx2MknoGiJX4lKsgco//qwOJSbJN0Q36OKBgIjTyD4WCYng7a1VG7Yuq0TWF7GY5FU6mJkvJQgv
P2NTHwkRxnOY1zTEV55ti639ELLJgNQK2lLtIB9+v41Zhl1gr3cQLfUX1adjAd+X3HzPkcXeTnJj
+8UfqWRvQ32/5EJ7Chrg4FAttWsyhcFEBck6TkgUlbc2T0ycciPacNSzm9trQuT3kVx14MJIOuUr
4Dg4b3kOBugJJfE9TFYK3meVma0reeBjsaIQQKK6v/v4l1ApzYT6O8IR2AOzJBWa3lmb0lfqEEMx
yQt/9x/InJ1TbDfMK+DZcpecEVfmAmP776R5vi2vACjBWVhtPNClzKA+9u8oPM98zRKPlDwzyZ+4
aIf3/I4+UKPHn8dKZ620LGDf7x4uPTGRt6s1vyV8KWGifOgWXMbhPoYn4fv/GDzIMjQgyIYtUUHg
3CvF7atD2lyfu2PpO2k6vQtmf3e7Z9y26eSOfjnUs5xb6FkaDr6vZW//vmZfErXNnALPepu5oZyt
djOvgxi1x3+EGr35bebzhuTBmSf+peqzWF3shHnj//OA5JW4oRBNY48lkkoP9vnwXh4IX/ytKicx
wLXlkKx6JAX9iSpsfn/3qtjJaXZyXFWj41FQjhKlOagLuGAed1oLFIvFK2cIawkNCWUOJlL6QIZN
dk/6EPjQa3r2b3DUtGv4JaeFAU+PKg40AlrqlBD8MV7S6P4BW1xmDGnQU0F9EB5unvfRobr4MMJz
tGH5EQFDz1HU9F7WXAmaBOfUVTsZgWToFnqewN5il7vlIAu0bFlftNd7VJJFc4Evrd4AhWMpYwK9
1Dgan8hL0UYZHsbFWIfQbqeONI2grFqPWhQXouMYQgkUpqxn4oGYV0K0QAWQFmfXQFGSf9INlsvL
KBXbFh6bp7K8Q1y7Bn2dyr9kS93TNqIT6eiRD+nZBqD0JvjJmng7EaGNGpXWIVjWVgvto72LINW5
JVijEj3tD34Bky5FQq+3UbCZSFrDuV1EEifbv3ImfCYv+smpNiBAVIMMaTrBr7AJclLCYa3MQ8Qy
SdRvtbm5//fQ69q3KC1LAyn718dpuzO2K7yu/AFXzAZ1mtlsdc3VCZwqp5tqT+ZFVJzffNGObwCf
/ULNIwhtnPI8ehTHTMqXAR6/ir2zzB5zVg95NyrRj7oEY1XDLKpnXuPqzBeu9PbMzI36HTgMy8CC
n/XISZmlfx2PWeuiasGmQVfUJBgPHX7/YA7s1wP4SfW7xC/CLyT+jYq0Hz9z+YKv+4dsQwvTP7/k
8fu09JvIGJtMXfLaFF2i6HZzPDEx3defKHq/NgdvgS2F9L9AGeMaIus4JPSi6J8OvFqx/QMEl4L3
/snfyAU5BZD/dFRCs280FlyatO4dd9awJDb22v83nQUt5GNMJeyhMVpXKnd0GaRusi/QU8iYTzxS
SAyh7T7I0OeVp2GRn4WDMeGlfoE9ElICRGO8iTiERXBC2CfxxNnQRQW1N8k8zY8QzL0Rin6GXOju
cEb7NwpEp2c6277C1k6iSb+VexAcvffNzDpont34UCjB/i70DJyhVQYHc7d7MC8JxN5coHzE+EK2
p+/sDA2IiNT7HHnXwp0eOg2yWAtMtVd2fqy2wRxTTMJo7YX6/1HhbdVnB80oFHNj+YL67zV5Zymo
D5EXLU44N6DIJYqmnRSyq2Z0R/Z5/giZeHwc6+7PpI1QmZcUkzoeg7AyophXDXkAQ29dR2w7K1EI
uJBfDDzXG9LZG5PSLX6m2cjLHnY2/zdgg4yOY/iFQPB5FhRV6+934h7HLsnkYgegaUfbe+AC5Pa4
HJpV5pMVjgP4D553LgOdqrrtZdhTuKOqPtPi8EPXEWddD4wgt8lPXMfARGSJAKIhDN/sTVsbDZ5R
INQFwBoQllrS6C0+3d21057euBXGlnOJNljt+fUmFDEwbIPuX4TP0EeOL83sKlPPGw2/WHJEFm8u
HKqHV1+L7gunaMlCd2UIHnMZ3nr1unn/LvODJt9Wc+CCTKEWGdviDzAdHCPJI5XFj9dqBA8iqkdH
s+lYOi9Q/Cwgb+rEKHc5oJNkY4pj4VJrBs4vp/H73NBP0hM6OwGrkpXGccQsf10OY0Oomgl+oetd
oHlAUtIUOc5409w+tjuacv4QY2d7ZCI7aqs0NOK8dro6DFhWGRFy7ZYwGW4hKje7jNWYD4ol+sUx
d7eKNJnhZL6a2EOA8BSsOYqPt+HPlyCGcL4MVgIVZ5luozHVM+wuoZQQJJXh4yFejwE60ks0fLGE
zzU7zk+SbfWnnllClUjqg2Z0RmVBHlXxaAYROjNFLZR9ErnmxGbql6PvUdk2Qz1EbGetKg6FGtIR
NbFWaUB/akDhJOpxj3FGSk6K4f8CCMu1cFltXoKPI/DTPiKa/+McJg4tLbM0a4RiRky5xzc8/cnX
spjEagTVxQIQlaNfPmJ84kLm/xOEPDk+r5wqwlJ/Nd8knt+rn1XzIwwoJ/2+Gf6bWPsyaRXapDnZ
Y/MfmRFWTBiuaT50n45hTVT1ZuCh2mQzUIORYIvgnWvb7JsJ58exvIJsYPFbfQZGLVunGkM1BmbK
wO3j2YujjPneQAMLY3SAzXcU5HBmKb5/I1vCvUHck6hguwwyFRIvsWGjZdO7XNUq9frcuCuU873O
adGmXFWI6ww9t3Ntb47QPyGhXB2IIf/Q7hxwzNoCINQBBdz1rEEqzytvLVTcUcrnoPWbmCG4BIxP
KCP0S8EjjK2PCLKaY6XSO/QDgpdgsZfzToqfg68Vz3oc1z5ty6f95agpeKidW9xi3gRMgTUPuBe0
AYRkv4Emv4cBGZvdwYI/rFHOodf2MqT+gATQ0dhJKa2yg7bUYYd005TGg6NZBd6SW47NRYKBx8R+
rriETLtjx0K2cyVX3jwjocSwIFq8ygiHM92p9mUUEMUEYKweYxvJdGm2GMScVydHwKqd0CF+cI/W
afcYYtCAgggOtPkkjQ1/AC8sOkf6ftAfmDsdvuAZdZt87oataXHNStIYbeoP+m+FX6INU9m5uoAL
zM+tQOE9aXSMLGxqGVRZJ9FAAJymgQ65duyu3b+sfKbaij8J6Cjx9ogIKZgf4gKDjKoTNHgSIl/2
Y3HiotwRoxtYJb5J005lJggcngTaSCpqZ1YEL/jAvZAJ4yK0OLCC8KqTwftr85UV82kBEkUXRzjb
X2S1cKEEx0SFin7yca+NTN38Jz3YR/Xrl4f96G8wJfukWCU5U8eh8fd7iyrPXwgvJmslaxk9dr/r
jZqc0NeKuMCHFZn+GOFJF3riEKQOcyk7D7GV3qTS20l1wSd3x7AaHouCdAXYGKBLkZKrKiofszLb
goKWq+For9J+23m3cfeo7HCQNnVj+bxTHaT9MCv6IWDGbMxjlCtIYDMhcQx7GJTsiTJOmAfs1AW3
5U7lcQuVA6GogJb0F4W/GgPwTYO8UwuNzHFeHjxy0vLUmf754Jjs7/uoDiPD4KiWHey0SOJtKCLQ
NZzDKlNXpdugLjw7j72cZ6t4Rj7d+NhBPjsAoMhb4m3Nsu55EAZVRJ7llVCcmGBf5uMKwwOUcFUy
wwl1L6zxpSEYf8fpPpLssOktsJ0HFVoT8raQ5Fx9nsozG0IWqP/Imkw3jba0XKsdE9DZ+prRbJue
Syx4gMrtTRwTMcm14ENr0eNz5BDvsKtIxkAUmat4+CrfmQTcz2COsYo3aTAiZTP9ZXj66qYuk25b
cYQzZ225JQlpByd0kjVcYYKyXoxeqK3MSPh6Q0rTRMV3OA0SJNwY5hUW2uFis0V4ASIg3XvtY/D2
rADgrBWUxvQZrYs/W3LDQ5+pv4iG4KeVVZZ/PBM7qhRBDo/Hz97uO35uPzPIaUlgQSqqBrwllswx
0wTfZCJt9GDblCX+fS5pAhYtUGNkJ2B8VGEbrTHketnatol8v5e0ErkE9FVI5L3KktV0R0MrDngs
v7omqXzk89+2u7PtqktE/LDkPiWcM/6sTZBDYo4OLXz2Ep6p+U5qNskP6lgpH8ndWD447GxCLQ0z
Ltg3iUHrDQBMhIG6nVBH+yLf+rqwuMuJUi3icmpN1N3zsdV9N8/i++kYDUEXJrGcEVU7JNub2Xiw
79AXgnW19sJZLzMfX6qqFHrF8MbvsSj2IPrg4A9myj1WOvb5wh+gGZ+nP/6eM8qVqCn2Rc7yGbEx
tP5hjGcMEtscUCP5SkcP6JlatK7qDtvIrei1Z6TRdS0kw2GLt1MZCI+7G0vGgw7vbx9IxjocFfDV
QMgvDTuWtfMvw0oKD9U9xYyPjRWl/GrvzqM7tpHYW9C9w3se/afl2+2eB/BXNm3zYvCQZqjUY7gP
LlqJ0D7gerj8/yRp/g4/e1avMm6E7FduRpW1qLmca6xJ+8+7KCvhUX4uCDIlSVWq1+GnGzK/l1K3
gp1AUU8yE1Q2XT1rML0p3k7tM3DbXV1DkNoB7wcLW12QIkVWD/vOoYEVn7mJH+7uH/Ra8lc+N6EF
uYnoLh6gWBxXoDn57bkXgFyU6rO4wB1qTClmVJwEKw01jprdX6ZEp/uDSTfUYWcvtIW7v757XqXY
RAJSV7GQA0b+R28lr3W9l+veKlIIr35PjGQgbYhJRrSK4R14G74h9B0TMxiWi/eQcppXutNuZ2pk
hm2B2T58H2kCI0JLz9avWcPIrvc7kf852U2kgKXrcd9c8e5Y4EEuB1XmCP96c9DncDgpJWMH7CrX
+2ypabbeo8FPADugVQHH3qGx0UBIF8JUjgmER49K/Y9sjgw2AnESfjp2mGukr0P+m3jI9w2YVvXA
8+mi6zXgmiTcUoNjTAXpLTmkNx9iV+E4oTh1Hpw2WVTReuci1H/weKJKqy5C1wmtaNWNyCNumwW5
YpXC0AAMhqx2VXW7NXlafbVS71svfeZIPXkGKnW0HDZbCJuOgYfpXwIwfLyKQ+vDXA7H2ArW2s1E
+nJhpbXZrKzlBfGs4JEFUytHQ186oXOLawxh9olhEMPVxWXapv2/1UXospbqtXp0EkPD5zcSTilr
P5BkG8xCbpaL3f3yG+gZ1mKxkrnXk2Xg/wUGkcy+9pPGWutqCZH+l9THS3VjFLPn9VekkuE5ZMYH
O/+5anbLJ4i/LEqrtJ3vTORiURFd+7iXYxTOxWmNVhNQIYu+vFEOOJTzcJpxQHEsbs/SZtLoIdVT
Dm8OA88hSlrmwFsV0TORsRHTGux4cxiJO22H1hGr32z6akRURBGS6S7x4OqhQjxKoXwdt2X8zGfW
oPZ1RS2S90TYX9Znc1cayOsxlOPLCPcWP+b0PmmoPkZC1VzqFOSHiMX13oA+Ue+1b0Ik6eQdr04Q
ZSoEGsovtNQ7VzmLORLYMovKflNUF68mzIgQ+WBjTij15sfO5C2kJJmwt0+1rfvlMPFeebVQcv5u
ychakYWLWOX47qHxN2iyX4ZSjAcPaoaT12fh8sgeWVb+4A5MSuNHPrwEhvZh2bV3KO5zOkmv/TRH
6gtOsutJY7RsxevKi68Kh2TN449Zqt3PLxLHs7M/NeyPHuyVBj7bsIkxHhkqfGNoMKoPQCGC77Hx
krhczyfpwbY204iRGXlVP1MQXtANXdVCP3JV22FHetNhbAwpcnik2LUUSdXzcX6dVQy8QwQ3VMp/
k9mlm7+6cIZVaNSPa5g8vtM7YzCoGS4WZG++vr9If7wJnrGlR4hD7OeaoHSDfd7M/UhHSMyCVHm6
vBV80JSSJn/WKsk8VaB/uInab626Pzh7eFDMQ2MlopvrvufFKmsGJFDPiSC4/ZLfgUNmidKNA98e
xKqaF/hTsMXvVsJkxc/lYUlDy85lrJlWXF9ttwUPNmI4kPBowCjmjlnh58AEHaj/YXBzyU2uYHje
B+el9wT/9pdvEL9cVLXjyWZQ/N1rHbJVunYlMCicsdxzvEdkq7yjVrERQPqTyg0VyVLcHvpDGs56
fH5XFAWrCxU7diqr69PdsmUDVdfFBlgQ6TZXZRQhHS7q/AeRaSy8SO8RL7mjm66UHNQWeat0Hghj
gMQMqWjWHmi7nPd8azGjL2Hx6K9iaybDNgSmJl9D0Y2+Sdj/Tb1y6oPX88N66ljmSshYDGOxGRgv
PklW5qmBYuL4Fol74bzAec6R9fthtZAHP2enjw9EmSDXPrHhtitrEHqRY6szvNDxc1pSk/ujhFdO
zJX218cP3v/ZLIKp1hTfk/jEvm/78/eJhAqko0CC1CSBzhtr5A0of3bwAxaKvvBH8Dm6Vaw2jvD6
LWPNd5pEvct1eKW4+V5lozaizmJqEt7rr8Xjq3llDq27xGRxqdFzNMv0PsWp5bUom3hdQCIr4GXJ
U04XGcvsZlKqMFL4j5ZuPkZvH89diP3YWhEFXFH+Krav7EAepGroJa41YfeaEVQbeiUe4D4+HwbS
NKLNdgXo/9TE7w3Q5fK+pIikTR4txeJkn7z+sEmPaHNz+fxv8drJ17BaOF3GQ2gIUcTsafhBYzPy
KUtaCzVbOKIC8Z/BjwgDmUVJLP9gdYQcYVGCHD/oI0lKEzmNjVSeuywi8Yyr0X+kaLxBfeiqOGd3
zeIHApW2mujIq+YbrPW+K+/ONbE5hThedPiSjW4CN06D2953vnGMru0A+FfOJQN/ElFgW2WVx+tz
aUHPbpC9P3+G7OrUmhpPqk78NCaaauBVCEuwyut3wOCRYP5D/oj4BiAh6cS9RInhmvOdDLsRyXHu
bLdDuIXiCeEI9E9NCDkGDAX0Frcuo6XtXpVKyJISgQDDcIoWasl616nBX0FBWAVcS4ejF7imzHPs
HcanNljwJXSmFxrOVwvNEm9hG9a1Piw3D6FflTH42zofU629VsUxfsx4G3JziJddGPbQMsoR7207
Hjgve8U29UBJCpdqwuJl1IL4VlRRN+nmbicrio2s+bQXHeBnVEpi/eVZ/+gepMdsuE9OeRoGiJOF
Vi/TzfJw+3+vdSCas1bG6ir5SOYs3IUqZotg2lXzC15qX/LHnNVpwrC6bv0R7HlYaNZXKRboRdjz
MqwmI+5sSsHvMlvSoGispOV8pWF/vKkzmcv+r6lop7PujS1cVMHaGCki668b2OvP9Kzy/gxzEZjK
HpKothCvRw13Y1njf5qc2FffZke6cvz5ZD9eicKIy6PsTu3KTEF8CJyDjDncMuLuT/48XUA1F+h5
06+tTj5RRCr6MQAoZqFyRW7+ySgSCLAVJ1u5lp1vlerKQoObURzbPdLE/OxZ7zcfRWkIc4fOSDAC
cye5zS+dHBENEb1gHNfbA8dm8wrhU8puB0W/F8QfAVrvdS+hVPu9SKdaqp327wNvL8Eahb9A72D/
4E/qhTzBGfzwCBe4NlORre3XHRL7oU3S98Sc+cmkH3xyZMeubedRyR9itEAKQ48nudxUAQ39g5tY
AefDiMuZJb2WArN3sZrtZbB3NJoYVnNbAoaPSyWOm5oFRb2OEUY+jh4ZAW5Ayo4JcapcK1uc2cwO
dOpj4IyU/G1Fhsld6Y4oxyMXT9pbc6udk7FYu3oSITkyjogO3Q9WFuDrC8F1dnA06935bQXis/lU
Qsi8SXYW//LsuTrhJGkEbxmsoS/qIFSSCj9WMHg3U1gHyY+rUDaGBSvBQxvwA+FZNug0uSrdRFa7
RXLs+vmTwdvl1/tiRYcE4TPhUDDjlygKGAyEcAT2xBd2Yb+s+UishIu3Rkw2Zl6VjJRnqgyxv8mZ
e2DEowtL56TCLQa4p3npXpQKutAYLiJ6/fUQU6jlA3RAje1CvFtVtmqLdSSginGQxierKa5fsyoD
bPxaPUDx4MhBAipOJNKpeRaOoUpPCC26NAhjLZ0JmRLmtoFLeYhajlhxUE7FR2V4WB34zozyzlfI
RWxZkQvJNtroFMOXRrzytD3vhP1S9fL+IQA9a3jypabBvaPEKwpKjsO2koP1JVwBZE1vi7RcLs1m
3hbSzEbhb8MIdliR+n4xoNx8VzQZjzoahktsx6RTA5iL2w0asiL2g/LnXgBjACndx7R6kI6Gq65+
Y1/ABTveHJ1t6HInFMcY16cdLcdyT0vZNqqull/mXWeFdoTuJZm7kznuyeh/dsCT2MwYIYFbWgf3
j+kbfLTH6bZlp25KhvDwKETuT9r9YmHMyKDMEqN+DXLtGR5w3OB4JdvppMmRTOFStdUI7UYnuuxa
WC1Ys2UlGNrHXXjJfB+PK0yPUNChhj0CkPNMQgBCNTdc1gWgL7FjSVTtN4u3GXDmletm8pvLZUyq
vnIzssa4jCSpZkmcPJulb8kM6HZE4zjfZE7R82zKHNNYUxiLuWhLbUMuKZ4IRoleF2gI39mdFnXP
rAERenbGTmplZ/rq/EvS9tcq6mkCd9/Qf9FL4C6tnVcBVfVtRHIjy+s6M6U4PRr/tOpuJ0ZDW+kz
DDlml4idDcrJM/LQUFamR1rXqN5Pm+nnVnzNKxt+CUmtC44qMZGxuglIpW9p+ryruwGq8cAIJfzC
XoeD20MmSa3AHx6FSdY4ej2q5pR6QjVteVNS8fiCvEo8hEsKbFJ2sPNjk+xzkJnM+UHeemSDMZim
V9MsoKSKDFEHjCV2x5cEWwW7M9bxqr7vdfkC6hn1oDpJBbOcJV6SD/7Ykrp4clfMG5JW7Xy+6usc
AEqeHCKK4Rpts4FdRxQVdOQaXxJ9B8EKSPRbOHSaJJ7W44uuDV7PfYMHPujGumQmp7o5jOEr2Qsm
J+RXXYqCKsubdpF05EvmQX8xMFG2wa+zv0jhQkGJbvoNUDcpC4ImYsy0E1IppRikFq5jOJGiznR6
0M9dq7Q5n3ZWpJ0+lU2Fhywpb0X52eQOTTdPcqdXs9H0d4DD1axrUjDKO8994+sf1GgXLM+hZCNV
IX7AYzpnHDG9xT8uh7l0i8Jl9EWCUgnRzT63bysOFEnrCpgcNWxZqjMZhPbz8EQgN6mMzu+BWZgk
jsRprPVGAdsalK+yaQgQfmMcgoMeywbq/Tod8AxmrOrnZUVzADyxpF2ow6Kj2EPOrvYoNHzl7Vl4
6YxwgASYyGyXr5MxowGYjf6K7BDWg2WI0R4OH4vm4lL8IFyHlhzqGUVikPvLsMptDWMg4UEfO1ax
3+xC48rkT5wya/FPW35sNJJS9GOGTD89q6Ffwr0F2yZyczmefG1lyfiekczm5rEmXxZxfAIUGO79
B1kFw/xicLDKXXVYbDsp1pSslbwJW7lsj1lVix95GhG1n3tg+7KQPA60eHnDV4Sm5FjmmwR9kf+2
H42/Mm6oeLXd1ePQT/QL8Mz9ugHMBwguhlgro1Yzt1qNeH5YX0NayT+6JbW91cZlJU4ySjIIbxVY
XREzYdtuyvD+T0m6mw+y+qjMxauRd8yNyJGyqO6jnL8YSDfIOrF5svDjinbKY9fVo+vez/up+mst
9jSC4VWBV4zt7Ikq3n63RgvNt9d1IfGG1YH2oi00SnG3JFUz41FggHK0uEgpcWBAZoSvrbVfs+it
CJ5FmLGTw6BUCtCfzndInyo49/0/eaLcS9ildSKfrBTHEVitW11PLuiiLtNb3YJqfn6S20ghqiWO
1QfBuJATCM4MCApdOumQI9ZbYzxAFFxD8yUM7I7K6lO6bLJZCeD8/EMvi00SkWZ/MYit+Febc5VL
G4KnSs+zlP5TC3IOePYMu35sATviDIgytPA=
`protect end_protected

