

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HkvkoCL0GWrNz7UZveLW08/L6sfDm0zZGNFYNcAn/nN//DPdCiitkWZaJWtNOusOSxOuhl+sv0z+
p1lz7dl//g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
krz6nWvdzbpcwbTOZlkbRdRmwRVOtCA4XeulIVQdqRCh46kKaQ1Az7t++QIQaaeY+GuPXRG5f+RT
/lT23OvjNTfUf7qRgYm7gawbEeSl7iLfiLygAHoLsmNj+AH8gs8Hs0aW+rBlNMkW1CiYm18CYdKe
BMk1gzJz99beaH3xgaI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S0rVRcgWQWVr47wX9qwnY6bNCk5yWX3QNuIUM8LuaX8hn/SFQmfJmPcNes8Folei/+/6+LEFm6Vx
Qdmf/pAXoMlDqA6Tk9J6e0EI5j98K8SO2xXJ+gzU3YFj+q4fP4roFCd0CsvGnNVnvR9QSY67D4GT
hyqra7o7wYbpUx2mTiv2gaLMwnoWnT5ZzsGdEf59HajWnwkeRTiguJpFlA2id/NPwWgZgHvKZ76o
YSHOqyB8zjfPqIPDhrl7blVRoBZvXmfF2bfsq19DFJHfG7UvY7EZPYFBD6y+qNjbBLb+5dGFTo4R
zppTZwWHLFQj7AvvDn7yqC0n1LpKK7npCeJwig==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FWYznElFJatYtjlAAT1QGN7C2Fn0bGHYIFjGBmEoLmnBxd4gbSui3fgk6xjK9rjjplTgHc9C9c6z
TaKY9/4GWl/7UJ0kugef7sQQoHIeQF6ee7w50lZjl/t7MzkZrTP5lkQthyugzPF6QCmhskF1nRLh
8U809RlH8O1td9E+1vzWR95+g13/K5/hcQtfJV6eMA0T69sJUMfVXf9ZGpdTEe+8VgstiL0bspGh
nonmspk+8f3Lj48HEmy9cJWNiF23grWiYEzGAr2f3JfUuscQoAvyNZKmszKrqZ+SsW18FBFVcMMR
aHTvY8YDuc/AQzYbOqTYkc0p9ROnWPSlq9UfKQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l2MUNe3fletgp7klnltItrRM3tzG4+89OKOcJcVRFyluXO3yMDNdtTkvc/SDua4RluI8ntOM03dS
viHFsuwjhwYJedBAb33tsrvwg7rG9tbt/LEG/pDQgEQsMWzKwbaNYxt96yL1pqBTCXrawJRgzhDf
3V9E64J00EAhc+Oi7ns=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OwI84vg3qgYuEbxZTTdCAx7VKjyk9xG5pPpZRLX9rHBXg1TaS1COb9wYAyuUkiMaNfwU+43FnUYR
zPr+xswATVVwp9fQM0Trz2CcY0oNj9FQu4CbQMbwQTnIOsyvnJwIujdxNq8gsEGemveYYjxPfj8o
WumIWJs8TCPZgcTg7V/Igr2IkCv5OUXoa1wEoiQnNS8hgrskPdguRrE0QQRg0ky2cZtAABfuiBng
oKj2VdTugfxBQIi1J4RVAb74Pk9k9CVJDv80IQ0VWrPTk5H0XM/u7z1dp2SYZUzGAyorho9pm3D+
vSFM5cFHGC5DCvaNPak36o3DJ+oTWzbx/S2Y9g==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1lsEBCKB2sqDzwDdv+Ksc4XOO4/Mx6iEV4rMgINzaVZhDq0geGva7klDVIzj0wbmLz8Oy6aAf2gm
jnjEr0kr4HwkpIFY6bw4gHSiuL42715ss8LC/IamaJMz1UyvyuflZZ5+w3WnVQUVJyFbnT6PcbiJ
iJr3kzP3kvqWO8h1atovR6OTQ2AeF0M57F5iLaipkXR/+ybFxvyZ9/Mn/qb/hckXmTrKdKyWjYzq
82ZZ7bsguLRLWbUGJAR1Xf2ACffKjcMtafkrD7fm3SKeBuj4CCaR/XIqBQ/Vqh0CD2XwAVxA4CgU
ZEl5yQsW3u3xjQa/H8EYOKX4ui7vrtobcsVM+Q==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JbNe8kbb6DVzM+tMySGJicqHJ/6WO4jSB3NMMp+SwRzyNOEwlfByQCraQ3Y3nQHUREYyNsKKEufK
sUjuV46dEokHCsNIUkveT8nCh+SboPES01C1eQx0/AR8CKBy6y/sWYwi+cSgLOC//wf4MVo0NRlr
eZ0/T4NrY4XEQRt4OBnbRuWmVqhfEtKNwQR7xNIqFBEeEC2O+ol58Gdq0+YRgeRtdKiHyAVVSxa0
bMzI/T9jTTCNMKv0ckDJ1cbw9LGyoLwKGWSWrxLIFXUBt+xE59mdFcCOcJdPGespM1nKJzWzlXnO
JERLLXL5nt7hTwByS9AR0qDsi72yUzO0FxCuRg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nIxk7DmB875soFV2AQWrZMt/6MixO4JJ3i54+8Qs3fBsH6g4tDNCPbpBqLlDed6dueueFUP0dHHM
RB9QdEjaoRsDWcLMgii2yco/P0MgRA4zsSUGcovzMhypbrSuZvmaTEzWy52XWlXwmKs7YM96nPq/
+TMw/n+G5Le6vtVfxveHYs+NHPeqVuCWg70NBSzkoShfjtC742vBlPPhAT4TNTPpDbQjcMK5+KMb
7KckSUrXtTbN2R3+5LJhQ0B7eVbv4QRxFhX3jgi+lsX0cRB3GokzHZJA8SZkAZj38gyTfEqTEmuh
NTect/sqzLJU6IZH233HF6Qn0DElnGjCYm/NQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
D0rl/DV2cnttRkRjmu+s9NzOBrUgyC+EJt7OrxzWrKZamdicpRkcpBIEHIJV65Nq8B17iN7ClzBI
chWctq9HfP3IfYh1QFBwe1Z4BHjeoWydYy3/uXwuajylz53dvBpMtmqcvMP0LUli4qN5PvwJfeWX
1V5rLtnVq85/s/Gp6/9n1YgBqnKuuTHJL7eg3NYDHSVcWR4jAC6VqXPJO6fUla+CSzuu3lCxDoZJ
9m8xBQkdSLEAtGzInvAczjtlri6iOgIKrRFpFDE9K1RB2XcWYHTFiDrvTpPvXEDV+CiPhcSs+0Hn
/jk8DAnoCADyResjFPCmbAUFnz6Ij69QyARd+nZOcLOpd9Qd6ibZOXC1eRw+iR5JEcz8FTzg0TXk
kUnSptoL5HHAyvYtPBVJpwkHsuRbytXDJ/pJovVShtdGPuiQMhEa4PRHKoJ80WhRR63PlFzR1our
D3L5aT8U6CbmSg6gmqsVYOwmetS9kET6vRHSpdNItIN/0FBu7mdKrxW0VJQfvBK2iWRAniOydHII
zI70Yz3+YYKz10wfP/1+tZkLcy0D/As7n7a7F3VTKpYcD+lsO7t6SfPpOJz0MeWsFeGu+JqayzAS
7htuqywwBetM1i3TQGoz1rZRt3i391tBavgJAIDJBUkdCqi1v64cYcim/GCMeG8a15/7KMNOP8Mi
Ys+EnO+ra/wk/vV8ZYh8+sIN8wUUpd1QVk3nFzElENsSK1WlSlWEzrCDlTHathyKwJWe9nOqoku9
L3OkialOFP9XyZSKTLfxTgj5AO6YEzD3qOY6/0iIR7srrri3sgb5FY5DYIB/31xPG1drnpYYmYYQ
WmQKtSUn4/pjGbs9AZoHQ4PrhXRfmGm+0JWEMp7DYjv2PqhgrE7Xx2U0wtq+y41g08DEOoI2jl4K
A2t/2BFaxPG+W8gMjroDmrw1ZewEPsGmUS0/FqsvIsSn8p2slWaBtX/mkZL/X5N4IIkdlQJRjpbJ
0GmcKptA0Ld4nqD4m6HyVww9MaR1GQmX/bDy95sAtkAe7EkOe5MpJypMR7SRHVxbr0mUmSM9YRAw
bq8RIjUiwZeN9Dudk0+ILKl/fdn45GF1xdm0ljZBadkzv9iIEz0GCdw5h9AIo/HLCTVrLd7vn44M
CUT2j88IEj9vc4P9V804oz1PurAlrhzUkTmi8Uro+pRcvM6D+Ni26ebQ/+rDRMmZyUMPwQ+EP51d
mLZzXRDUq6zMx5RArFKfOerzbkHpSQsgxIk9MCJMP5l2/1BsLr2DSn5OjuHDatsVQuPecqHo1ner
QpWyC93d8GbektmL2qfUO0VJ9s/iUk2Z3ogh9t0amSL2+cNRpTfJRJEIN/uQH4C9Kfg/ZaDk6eCv
JVAxmJYsunqVRfivv5cPI2CZ6hb0BvpzEEGAP2hxSjz7r6gCwZVL41+/qlnvY3j5TP5DSn2GZvr4
2halpgHg8895AMiiMFrW16CQRHLhEylbKQEx+8hBiDNjcAnagrHkTRjbUE5EI8WCKW3Jn0obivu7
v2JTzS74zrQW9uocyeebaXmrfee5Ayl6JuKBXPzhNu7ARChHuWy74dSq6WRF/27VWwnKFZOmp7Tb
MX15HdOSlwCo1bXx7D4rXcqjsVAGn7ThS8ndzwpfcc1BUIt32JrJYOdO1C7O1GqAowyXh4rTk2JZ
b5HymF2bEcugXrpki5z4br+6OUmSfgLpowFSqO/FVcshLL6GYx9xHtc1EFuWPDZJ4VZ1RM+iKMAD
Sy1BZhtUbVROsdQdb9fChUFysc6ZCTwLRki5WZxe4pgJydNg3LzF+QhoFRYQeVcYLDUKTbOnbdkx
fKfXS8X8kBaZwjMgtL6owrmIlh6HGxpAw+5Sdl1Ao2QZ3OQZQxkAO5TLgRVTQyyJiIEm2c9Bfiz3
RIx/yfzhWToG5QY65CMdMWrlqbRie28OYGLteQ4DU89RrbJ4yt3Hot0wRPO2WFJikmOQqlyPdsZD
GMEdX2NONss59jWF8mtyqyLapA/kuTE8OHczmvrMl9m2RKcG1qWda15jfW6Pb0tp490Xw5n2aldT
TyGk8DvzObdbMlJ+5CmqTWui3+QPWl3xCWDErIDq9i7+XRGEndQwngTyCYyQxWcaYtIffLZgoeqK
pdVXwzwj/0WuP0iCbqs4CQhpOtEBDijrADfJs6gjYjtn+sHj6wTzYhRKR4Ab8eqUv5pXGcAGHiyj
D92M1Xrr3j7cbYB+o2agkK7qlHMzKbnm+J6fKWorkNYR5t7b1pa2i0cIy7PJdechZIFRRiNWzeLC
/Qh7/HWYFGALzckTL+1Ci5upWIqCRd+hLdHOaYw0+8pO34d2a7uvo1vCsneqI84QgyF7MDJmgoRM
Bq6oQub4AO9sohpEa8ceoWdB7UddSHKHLFK7k7DoYCqjSAymHLtJV7OXxLoXIi1TrXEuBADwX1q6
BMrrdW57PbWi7Q3aOcFChSrF+W+FEwr9aFnpwmt9858CVnWn9c+D69HCmn4ikNyYz39VsApo1EmZ
KpTVkGYFE4eZP2Lmf+utKIT1Q/x4kbiPuMGLb7w1HhNzf8mLPwvLBCbwyiMjKRylJSjwCC70/EtT
WNcQhcAAzQwTBJcv/KK5iTR3bY2Fr7x1UMBsBZd//DI8WikinkaZVlepYJfq5ZetOZd/dQb/vj7o
xgspKEM0dk5dIAF5GhbQFqNWBU5H8zsPejrhwyYIsK/MITaT4GWy179AZXhyZPW3Qd8pwU0B1A+m
Hb85M9/mbXIgmtkW5nEq1bvBm9myY224XQUd8sxjxeVPqh3VA7xO+6IPVc+rKfch6Rrv+EW2o6pt
miMoMWxtisyQvuXgbm7edd0iZQUW/3TvtNPkZBqdrOYXvB+uHWz5/dzo9fOsP70Q14xOyf7Jz+C7
pei5UuqjYVMkGXxLjNN+MuoZWVrkQy3JRuBvuaa1ONlfbISkwKWHgc/isfWsDnd8wSfiTNjNUYSx
KnKIWPU42O/iv8Nv2nSM7HsUgyBYDL01/n4zSzmkSVmSK+F/HtC7czcGQQMaRaLhfQ2cUcGXy+AX
oetHD0yd6mScp08jDq9fk06Ksi0bKp7RCyXPo2tpckQgfiHd5pVBPLtJ1YUHkx2cVZEB2iOYRv1w
BXtyl+F7DSKXh4cfb5luyre0CsAw96z+JJLgsAiQBQYdA1LiMOeSIUP9ThWXszNQzqMhFHJ91mZB
dIreNCnG/McmV+NLu6ipRVhTm3euogRKDXDHkSW+a/9tbcnYC62U0ILwytwu8idktEO/WgzbwVy4
SlP+j5Cvv05Ro3mkwbSJT9vGufGakh9IIUaHaF4Lz8EvjpcdW1gfiuVM5OZhLOn544jOdG7tKZUe
PsnL8AFn1Z5IX3f/moqDJk6/WLBA94LVxZqvRDaBpD8mP0nIOrS/na5qb3/9gSJJ0e6SQaHFDrzA
3JGn6XIqGgI6ySXmgxVtD1mDCNIqScYhiXGwhOB650ywIaMd4VDVexiB9U01F2pk27We9kljAvU4
wsgspe8Z4SvYuUWvKJCiIt5tca2h0+LEiPLER8e2aZ9ypV+9LXGZ9HALVbL64PY6WMJTmW+JRldU
KKDSOLwQqZbV+yDYuDx6fuPv+QmofCn5Zw7y+dwkan+et7bxVIw5RmZc1ad+q6jDvZtEBQOaPxsp
RbmiXU7YALkiMDQm2a6mSRJcETg+oHUi92/cci9Th2aNSPgMyXx49jhcSyA/7RS5cYmj1JcVZrC9
3wSaolVr1CGEVMsxyqXPCa+9RgXZBgBV6nOvl4xS3uN3NvP4ayCaT/G+X2xJ45yI4rZaADFLRUGI
nN8pYsD6QCV54wBvz99GfN6nFwFzXuIT1VTOMLCVNctLU5ZQufmlVh/pc2z/Et3gO0e0mAqdbLpH
7w6/8F10z5gzEF58heuIDP3kvfxgiZWi/2RjU5YXdyp3WhdZ9mBxsF9yPq53Blb0qo6lDeGGlywx
3pYYiR0VA4YtDDh+4I4PYoYj5ALXsPrPHlRifMSY8YbR6l+n4uEDNbrT9bWPQ36mhXlgo6NHt5ic
uY5B/L05ecT1/6pXX25HBXaRrBY8/IZOa0aX8cBn4caMS4ATT+m5EAT4WxyDzeDZwme/ign8v90Q
/ZN5RB8u5nIDwat162rvP+XNZ2EYlKppBmfHtDcuoedlUHuWsp9WY/2/SsrcpkaW4cJ9rNus/0KF
Y52J8QlRVDXir4aPgRjLjD19aKJhqcGx3063VOAwWJTCZfXY/n4dncCP5eUwEfN1Fk47gV85Bwmd
8S0VBRIFydjSLZ4tvDfxqZ15vdqzfRcMLbVyoAQpFy1qLGAWieslQnXuq69xQB6K+pW4tZsBcdMp
ghW3zoeTwJNdDz02ZROFAZWDfOOSssCH4z9W2xAcl2hakGVmU9U8xYWD8ukpz4dUN55S73D8OfAk
1aJ4lovifEv+qpnFjmrIzhf0U2RQvpUcF/i6GaBw7ObTpsMoUe0DGUi1fwzla2sUiHIgBajKR66X
fficVFdoTJZX93IgX6i/e1Tnu6wwoPkRmcIY99mQsyJPsxJyqNWcRar9sxKJ2k+y0UyO2XB1ZGoY
QIEuhH02mDU3xh2bPIA/YXR/Dpasu58T8LCktAnkwLRa0jRc8mQCVC87JNIT8tHQq9ZXZHnpE+dT
OAScf7HSuaygU+xpGZEeWQnyGzbnXpO+UiCclNOIlZKoOSRgc6ZJkS0iVy5S05Ezebkr4qQ2VIPT
QE+OenDKAdjlQrwOTjNEidepsHa9ACN50NPJ22uc/jhKb1C4YIizlWNArBd93d5mvX9SrhnzqM04
ho84CSBdvuTku9tBbYlobrE/JqvchizeBvk8VLc1kCF4lgObzGcKM3A2XZuvcm/foybbWjZHLNmG
QOjwlmhRTjA3cXmDJF02wivK5YOY/niMGXD2Nht/qVIYD/u+wHeCshmZT6FSJsqUxqDGSwrRk/K6
/eWjxeKoJSfRB1G1A/Zu5Z4pueo4ZrvdTqzRqaEs54HxX2sH91g7yKIo4o8pSbONHyyzNxnDO8pD
wGgyoYnUdpKukOgV/ehtosPncem8RS0qB+R9fJ03j06CDpFP/StqZw3dr8/uQZ0nEW3x7S0avX3i
2PrDIf1xFncsRPyrjjpw9DQfxFR2/4gxz2XIZlnDIhq2dOwk8StmRY/Mu2fFQWzcN5Lz6WcU2R6I
AoWXJm7Pu0tSgQoQFpVMr5P04cAseo6+utlPVM2bOmGLNZrKo0NcKpZEOkx/pBeRAoqEpm1Ztcvh
uvIMlcU1nPy9NvOqDhqx6jmbnV6OPXDX1ViKyKoBjE1X9YovjmBAAQsh+HdqY83akN9rwgcMkivd
gODARRY6oIAnlgB022Lp0fNwrtist1DBwifCBTuN5G1Kp2bbtBlD2G+B/C83602ujMFBP7E8Nc3x
WiV04prq3fmH5ZXf3QTb5gufOuw1cTSygGy/r0Exjn6acUP/fVTlBgpkCV30Q3i88VsfcanUFJ+p
OTtWxfVnmIuSdSRaDX1dDaJpOOqFi+3fHkaynDLf/cKy8SmmfW1Zoio0DiHMGT+VjPe9AbfQ2AkG
mOBFKfHbv9JLmSr6+upj80K0iBq+j+tj989GavIeA/9pf1DzOK9LHKDYCuPxgODAn6EYU7E8zX6p
MB8Ytu9ZPou/QlaO4H7heBN6aVhnbnw/SRoFhsmlRORmsWTD6EuDCnim5sNECBIuhrPW0g19m8Eb
jkw/XqK7IjeM0YNQpE8xnNdgsZhNV6pNs+rKHWsNSuf6/MBR7NMN1e7aDt33FuCFfsfGvjczvh1Q
ROlI8+5a9rqcpYReE4Uuca34TtMbajO309UVxuFY6MJXe5Os46V0uc1GplRp9kGf8DGLsE5Hau25
bs/jJCr507Xn8vufpWhZHs+kqVj/vxOBqyBr6TG6D4CKFK6h6Kc9cacf/pNVZ6V4K97LAW/7ktgx
hOf2AA2bQFujaBlzDz6xqGD9oZZM98pmQb3J0J9g1M0aZU5CiwsoFtI02bIT4iZ6YleA0yMvUSvf
B8Wbhc4CBNmSSdGXiuI1xRsbSMGezRStaVGFn9WGhkNhE+Jw3+CP/T+IzzkB8sXg2UKcl8xy4Cmy
JXGp/SBEK9ZrOWICgScLHdi8AgTi43BuMDUkxOYPLzcRKL39WPE0558uKJNP5xH+RDCVzMT8RoK1
zaJpEvMRYZvENT/MstuEQezg0pOX17SKiq4VaWpuVKBoNHTWt8Kv8ClgaOeWcfwWHNpMiIjqhQjk
PhmWyy247fteAwqae0klkgc5O+BeoWdCWe1W93r3x46Nk82YmP1rqAY69IQtQIPmxIZ4KmzQiGX0
Fp1+QxLKBTBZS0tWCFppY2Sjro/bp7TuSoVFGWRFXTZMkEzA4jSYJ1WsXORGWZ4tlgJaUoyIaFX/
sg5MUxuAOEvlVhPChrn+SIbHz/Mq9zZyMs6Gp5oq/Zc/nn1p94kQ414sB7X7XvYIaFgJcqGK4ufb
rjH8G9jRF/+70aozCuUgmqiB8WzGEUsgP8l3DgSugXf3icH1/jP3OYRqZIHrA5KClRX1ojFZGo0n
J5vcm080MLSWoZgIGYqEshxaFZ/tBxIlcFTwXzagvVPcVEA4kQzkdXVxsrEDahik83DScIJ4dJb1
Nn1JNsXmzBt771WxllbQmi1ZGbs9AZl9kot4HKjk4+Qxnr5jiXGcMleLWnBgpaXlgJJfB+CPinUX
n/CbdR5Z8guWK51RVDB2mUva2u7ecBF9YBwT4SFyJW6cunbqB27I+UQcHvA6i0XUaF23vbmiLCyT
kGm2XT5RWBQu138c/aUqYFjXH8bPpBwjHEUZh95l99Eq3xU8yYQlH5+AkqtRlzAS0cqb16cdzDBL
pMze3uDjoqY209QoydbKq5bXdPNQDuv0CFrwcL8Zmh6xV5feKfwNS+7HD7eL1lUPU5zZSSQ8dSTm
guPYm13A/Dt1YinqsEqA7WO0ndnyCshRDYtCvnFXtEnPacEcAWrngsZJcuGGEAUbmt0VJveTmPr9
NkKSWCaLROEwR6oylC3fX2MNilnwn0JwyRES8sN8/3aQwNI2QJvAphn8FVHVf6NpJLLMMnf09jJT
h6gTe7RsZvcGwdrcqm67+krpmjhBRdDoIPUOaHm+WJNKAUGJ2QfT3O/RF9B+euZ6UEuU40tpFt3W
78MOPObUU4UeW4x9oLM4s/9IxiBeax75LyTG79+Ps7Th42t0uTPxGEYo/pV1TOOcBdBdtSVHIZZQ
5vbDHQwaNpHiyV8ZR8x5lRoMFC3/Luy60Dg7P3McNjezX7xSd+7h+ACq8C84jjsBTS0lJOBtu9VA
EKYCuv12BP4mOjUt+9HinK7t1LbD9DedVaHVDpbOuVEB/r4VTKHu6SWaj45YSJfuySdbnIXs/5+v
HopjojX+HDJWFDYEwgUJpJKlXxizKkSLzWFsCHKphmU1dUegMNYdwDjEsIJ1SwO9cU1W76o9sw8W
4aPRaGSn8gZXrDEGtLNsdV+vamUXM3b5CLM7dLTqyWaKyzKUKjxArCoa2ycp9/o99fmq8pXhjMsT
9X6ReOdF8KYAj3SQSH51NQHsJOlZY2aHenbP7ynNHmz6LJFsyRS6sOWhsGs2PcDWEJprJmx2Uvgi
nt77K+UMMgzUeHgXyEfy/BGAiQnV6STw60fX2NTArsq59tlz2tEyW1EL/TIkU+xjte4DACsKCa2i
jQsEykKG0LzPRtoMD4Q1KB4qH7xGPePFFHvjPaYyt7RfC6NJw4Qf86Gumduk7GFUdjujsDeP30GY
em1SyifZ9P4PiXM1s0SB+uLjMidmCwIMPOW/v9ssYiNCuRXgF51Fat8Tu3STg9M5Wgr6skj3rKO/
c/Bwcm6q3qPl8U5Gs+/i4xz99xQclcJytO03zxU3e7cv3EVzHS/WP7TqGsa4ZKMf6mtrPCjY6XFw
X4NeRBvzhuogdtEGhkHMNRMvua/qN2G4TNA86pSArbnLw1PE+eYc/hNzRVxXB2A7RlkDYAqVtNW6
zySuEJV0J6m+75yv3MduH8b2q7F6Ezc1Pz+vB+aVuc2tP5AhidWOOnk+k5QItvzNdybhrEBogZXV
vWCkzgRu11hE9k7WMeRBkZT4lBLvbWfca5NseKAIVfxvFdQHfpnm8TMTm4tUwGrdmA7oyCfDV6aW
JruGRtXgW7ROFkEefTZX9Tdz5+CxLqgIj33f1Jhm0dq2y+vWqs2WOpNGH/J6syYe0Ti9h9k8nRjb
BZMCzoMeJkAyPSYMxhkP4yBbzMOwAWcQqjrA4eG+JVbgLraJKXzkUoXn6wRzl8Qyl4leL8G11pur
XyETcjuzxrfVS3ms3WJ6TGh6zRCDVGAQvEX91/RU6nOkXIfK+7xoUrdVc+KnNATw6XhlsR6xhrI0
x9i31r9dPSHSKFQ17X01OxK/I1yI4lLKTvk9G6wsh5st4N4sKgsPjNWJnDNjqzcrqpzqIzdXk+Y8
/CQYOpIu1cmqDehUWPseWI4WwJSueVleyReNGuUr+LUKnA87ounwkSgm1Wy9KgIWhHfSjGDTNwR/
Az9JSpLMylxC63xM4ZXXeneZM+yLXjEOi/RJqu6I3ivw+tUl7BvD6H0BzQ26xlssnZgY4cKe7bev
RXLGBc0QHBy9F1kXW5kmxGyllwer+8pNV4W2erJSl4cQ3dOg590EvZR8HTAsRY3Dk7dTNVuqynK2
nCLD5gVJ1Qhqs3z4OGcHsymiXIwspl+wmprDgMaz76pNu11AKXe/NQ5EdNt9papCH4+ir9lTAer8
MGDq17bRAwa9l2g3cpQ9YsctbdGBDQCXlUepogP+zL+4EreAd19mUEv7+ssRpqhgzh7++mLnUh3k
fz9AeMiYBC5vIFItTfLHWu/3ZO1WU1Ev6mY22wsWPpMx0gyQd5FnHeIc6V9/aXrnZpNjdBbTFFnu
8oWhC0BZhQqhuyvIsimHLSIU+WvyfrNLQFh17X3XMayO1wGYWWJVrPnagmm6RRDnNo3gmurjwMn0
wNB4kS+SxwtkaccOkqGFRO6xjF2aE8hExPzXrgdMskGsr7YkeEQM6n973VyVnxj8EyxPRZQ9X89i
ck+HgBOhT0wggJw5ZqmlS8aTXSCGplMSji7kKX0qord26MbkBo9y9wQSTRPgO8PQIYaFUjKFwrPn
GaJ45qmX99iq626nlfsYfW+QvJgs3zqJTXIyAheT3UTJlRaZaXA84ohzNWstp6oKvN4H8TTQvnJb
0huOfrCGk6RB9F3R6+AUxa7DqVNVAsFeXBHlc9zSg2TtKSqjnHjOLZ9N8QjEHnsjdIrpjJwThhqF
328JHk7SK7PbJcImCNFBMTXIiyo4Psv9SJtmXuX6rUl4m1CESWfAcYVS2Rnl+2x8xPy2B+ihI3er
TFc40rcL55JOPtmn7yM6CRF5OO3DbkafuNcOUcX92na2rfKK5zTcEk/8O7XZW2MO4+YTlEbMBUJX
anugEBBXoj1ee96gEW+770OqP9azI+2od91YVlq/syFVYSdxitonOnldnQYh3FRdFTuJ4xe6pUpl
0YWBRiyQhcXQYjLfwq0WMzwcdHkCbNCPP5m0ohavkvaZwlz5mkn68535MEzDPBOG+fiPr4BxWfDS
CDGfSqPCSvzlWKAnCyFromdaTINTKg1+WvzOO5W2awNUuPk9NmHgfPif3/ZgbV+jauVnOCBlyK7W
rLiLO2Dr8J5cc1EOOXQHFqxHVxrvF/h80Y1jplzFn+XwV+gAt0v6o26zKf91TxxUT+ygdtsnKZMe
0DFY+BQ8HTHb9XZMRoEjx/InThdsrrBz3BCe1PVi0Jjjk36x1+hNpFMQrWVwpQBGuNPanIGnwbMh
dGL8GKKL/7937FJZC0l8AvnyhGIHZo307yc9U/xUQR12AfzhVxmwu04/C06glBX1Uxu2PFKl0wPx
CfB88JZnirq8uGJljfcx7M68lo0/JE0i9b1xEi/7Lkr0IFU2+JMjUloZOyjDnP6mYi4hSat7q1vS
6iS+36lwVGz54+Lq0vNNIxL+1bhww5eVsBgd5nHW89hp+kW8qkXOX9T4+FmRxo+4cV48jLldgY+1
7/w9E2yTKx97UDQEqnt/NWmMPkDtBCxPPlvduL46a/DrBX8OIhE/PlcjA5WDnc4q5IOwhdar9wMP
xRpNmBAFQX3UBiQjq7TaYm1M05gNiIGSQvt5kuC24tqxdXupG7ixBuv1LMVUaYusdonlGildz9X+
nNHx6lbpa7QLYYc+hFrOIcXDaMbimydJktS5jeqAYCiY9sa63p0u8V3u53R82E3hw+xK0ndhQjaR
HAOZERUNFvSb1EaSrcAyBHG3sVPcgYx983VtlVFjsOYvqZkZXFO/tZLs6ZmHw3VSeinTjI5Pfe9P
2eTiqv2FL0kjk8UEj9XRj+nC+6elN80Co6c5A4bet42IDbA/hdcVZcnPZcpq8vewx8GZkCo7NUe/
hoPriKLaMnLWrkzDBvQj7nMefQ3q2907s13E6D1XAGx4n1N0vPVP4hDTQbfVkGg27J724loT5TXf
89ReIrAsV/don2BdRts4DPtRMK4bnqzzNWuuA7mbU7EpO0S2upFNNaKuy7njGAGkdkxk+kMzLXUm
OD+AYQomFOakE+hZPFvgZ6v6UN85a3joAoguG1MebG9EhJF9nxdHvkQWVxsY7kVOsM3cR8mh1/SI
CUdV4GkMdILq1E8rakhki9URqvvCQofILSgjgz5bfFsohMe3nTarseao6nz5/uEYsvDIEgGVMdYQ
0ISmX3UA3MWWpIRGNv6nsnlKrDYHknTz6ilZpzA1c3WH0HjRaymChh1XryImvVenW32P1IKjpaKd
9RHhsRZvuCXo/ZdeZgwnYBEDG7eZ1ouThGSyK8AQJKjV6F61xrTFtyZ2SLaowrKmsgU3wYFDCtcM
PyT5cK3Hx1RJpjq8+IPeIRh5QSHbRWQreoaZGbXQvDZ4uVJ3PdCnkZ+nmwAznNyzFKafRl0Ukkm/
nlI8zNBkqeWfFJsQfa5XwYWfPNLXX53IrXKn3JlcCGd4k3GOFCzvllhAqnRvMmMyvyy8ez8ve6S6
+4rBSvWMeMIgQJGHI9QIALaGC+uPAZgibrZ0QaK1zJF+Vo0Ht+ydkVoAg6QyXO3sAm7Pe3GeOQOw
xNPUgmqmj2PZhtaSY0goQFzynhEUf/EKtPNRN2ktesAzuYbuJxqXAzFn4C/hB/nRMhfCQ3bReScA
pbQZVd/L1NKlfd94Ha4gExFnGAqx/EokqueBOtfWZHxD5x4HXZVGYAX1IZsPrV9B3/64RmJjI0FB
l0R9RYZroheasI1Nu9h6n6Kngj1UIO0SO32aaVPFng+00aFMvJNQgJP1SNmMmvKChes90YvnJoTX
A6OryqSkVDjweJgfHOwGBAQQCKm+4+2Q0JqdiI5Rt2URCWqb9xKYJ5/a45DsK/n76ZOLf6Dtoyqm
zbp/NCTX4LJHOYrJVQ5hyg/PTytwzeWk+mQ5Q/9pMHF+TQitpnSXPBhLF+NSSxbldmpxNEZlHPHH
HFM+F3L7SiM8sMXSBAw+d/qdGWj5dAw9tCUmRBToVL8cA0zElStDVFLO3+g5zvXHpD5kqGH5oxpl
BMYM1lLn0i53Hsipu+66o/JN8XnfiOIiUD4ikT2BFY829P3i1vCLYSnn/w4XPIYXg4vFa+nTuWz5
tfvUrcqTXY7/xfZWnWgI49HO6Ay9ujUsVpzIliFNBcFdMgaIWnYlt4v31fqDUL96BqDkCv+6+P/v
DZrh29CQrPOMH7YHyb/vXUraFZj5RSYzYk2F/fIZEHm6Up02NMVGHBO/ddyxRTGWqw3qMsXOlvRD
fDX8FY7IKVKNJcylaV4645H2vq6lK9uDN2ocYfV5e09QdXTDulQkXhEYz4jaxBbQH2uv8u/c8R6n
ujVCJraqUjAZDxJL6GuLqyji/pHr8RyFsmYRgWS2r5dcXVURmF5OY9QpGT7lh/GQ1HocN0Y3xcL7
bmjbSx11bsvqIRlSZVlhDN1LBdZyfqYlzK7snaqFO3MnB8uBf12xjWSQ+yLhK/ZZFxt0hAtoFWib
vBuqtmuzWSkSkGyB7R8By8HaJzts+gSqdWDVS9CEVO8BW+9FS+Xet+Qxs7Q2PVOdm6oBz4sSwGyN
1Uq6nJXHDeEjK9oG7n5/758YlftdI3YX1o+FwbSD2IYTbGe9U5qgLEMquZhuZfKiX/VBmjVrHHjS
y7LkkiRbHXiA07R69rgxS8cERKJtQUT/LzBLkXyBeqKOmI2n5KyGAsZ8adkVuiK14rBGuGC4Z7cy
XCXVTDn0oNl3XLYXd6jBy2ZYmCxacBSLNHKDfG3WLx6ixbCYf0H+7PtUjcUUZEmGHauEjgdgcAun
gcFtS7sIt9qH+l3OKiQHjdAiiLSQ0cziuW7jVwu3qAW8DdPNS3fUIKXVWQCAwxo2nLX6lh28lm4w
V6iizGUq1amNneOnX2s7vNCIdo5mxXyqJLnOX5/SIlozEW0h9dZmQ7MZMv+gsfKnQe4VwdqlWDT1
Rb2+1Awi22mFUfhsyOsQ9vvH0RhR3rjeiBU5H4fSqnMvsPHqYAIHphv5Dbfl1lj7mXCNr6715Bv4
NWJJm/57y2X/Sez/YzdDUxJVTggKR/z6MJ6yvRdar0w75b1/y6FjMf+9FKsedxgxy9ZSI8JzI55P
H7ShYUHFHyMzrzB6pAAITYHTJ1CX0mtJYwJi/ez66oX/ej7W3MRe0wN498djeu2/dVkeRoF00KF2
5pDFHFBuCtq1uVgAM6B9MHeEf1sdbt6PKa2WUv3wm4N4+adlkIxiGKq3oROGBNwlbP2QnBBh8sYr
f40Cx1uWh7aD1/N7mXvYo4ESwJzuwvsY24+99bwjZ+qD80oELsNsN0Bun88nxXOgupIJQsgUwBZT
gp3Z3Wx05OnVMWYbNEZZe+zd62nLCSj+O6PohS63iDMbVyi0qi/aJahH5ataYLzJe91LPxMS7Mi7
5sUq5jSPSzTO7XnOtPr4CLKaYGP0Nyo3x0affhkiMXCYuHHuxWrSdoDurRAhEY+dcd7mmZWzKJH/
QOJ44kUyUsN72LxE+hdmmse+1dOkPVt9iLS9PIF1c+v9PRMZeFLWRWKkfA2RYuLr4vHTf/O/AVPN
SpfRJ6lX93gLy63BufdAPcJANpTSz65+KYbFHMmSH7EGgR6xWWLF5qlHa3MBxA13UHiBhmpRhhnC
Yl5Mvoj5AZEsQeGJFM9tw6L+2tHH6RMLuR3/hMME8KrIqOw194qFuBQh0TfrFfanBhrVYuLnMbSf
2J4IbnSPBNqiARRDN2esqhqjyydZZJQT8Oo0U5+q9w34DJ4kTuTtyG49GN4DxxIMJrG3s88zOg7f
635We7onHxjwY+8zKUhdourwSHVIUyBEFfRhHlQ0EUkrHojLX7u6o8sGy++gVpRrucXO4osP06fv
RkvIahDaYsDuIqGymc+WLPSQJSPctuBPbvjzgl8q+YbA/y9O/xbtneeEOPazT8JypGU2u5HkLZe1
uARCTTenm5AnFbLmpmK9eUuLr36db7siSSgxz9UpH+6XSnZbTctGGN2Ayidn6kcwFDUk8RDlQn3u
a3/g3eox2wMpWejK0ylSZmBkDJXZBrmyg9uMSGnJHPDflDTjMxX2f82UKuuRfNKbscNUXatIJR41
3uyICOFCDxOG+zUyIkWTcj+Ttx6qO2TMP0xU2FA2I5hl5Xj0t3NWq7+3XROtLeSRCWKZfzJjCAku
KyYSw4KeOEwK0YD5GlHGYS24H/OwhgiyWpiDnK1RgkJK4lJjjr63hYzI6S++bbsC2tdMzqJ3HwRz
4RWlWQm4pCJZpiRmPLK/BCYrbLC/dj57iIur+iS78ax0gficETXiE68F/Codgf18nfKarDLkyBt5
fs3oD4UsXSR9TJO6ByW8StttPwxqUdlPRtI3vTblm9qaKD3V+6HjhETV+UXNyZfoh04ZNZwZsdut
bFzzbIVMOWBTaaTqiyg1cjtjxisEDQP1WbhjosKzHJiBCW03hgxIIV234yCgZEJLbnptANaTQFNw
cWwsyMkf0IVgbEMYT+/smMpP+3al0aOuxSCJF2o6Ude6ok+i1O+V3DYmzb5mY0+3P+iME5p6PclI
HJ6WNTXNtnBg6Qgq0yj5Bs6Z+gyns+VCgkgSlpb1XH8/UMcp7GUhhYWGg/nVKSobMMKZodeL/2iW
N48DTiPfQIpGnywW1BWpXIOmDGVrduo0W+fYrpuiXNIWGszhjMeCx1mboVZUMNk2AHwEw8Gr4QBN
kT5idQ1B2YzZ77bPhZ5RoTZXZZ+v02YAdHd1EctDRFPXEWb2l4U2i3aB8eLTsBlMNDK0nX+m74qY
xbxpvsUnRmcsW+1wbHDvmKVGhqLSMNPDMQ2q3ORzHrS2SdP1XH1Fu39xojbxbzgakTn63rgcnZTW
cg0TdEcs559YlgkeZ6qp+A4Y0BCj1DPXJlseABD9BqPsNXc4ANPo/9cPapfUte9rhLpcflrn4rRN
bVg6reC70a5H2VEyBTBSua/PVjJJNBw8Gur9INILg4xRA1l5KZ567OQm+GKVKBMpMx9FsXXt+euc
nxppbRJkZjLUwAnNk3eeYvfso8Itm5mS3Pfy1rjnLlkYVdYWGjzb/W9PkZGS2focf42aDWtGTvep
4djxypNAx1R69n3T5mNCCThQADYZsUbbrhCEIcySXoqFZswfvSLGpMIVS8tEnnuiHcHq/17VxDg6
2pnxIGvA2CNB3rP22xJZtd3+dpR/VjMaHJr8FugoJCxH5qgZldKEcspHvvWBvdjs719pAQhsa6J6
qEdiCUUNCbeRi41fzURUvRmEnYoTPmOedf2/sG0PzaJAuZAjuf3DkR/MQaVUFpd5VvBAOPtVbF2w
WDoBigKV794H+dnZIpFOO43okPzVu3FwEV6BpsPTyhCQe0sBEDTzuKeoNoKb3wl/p57ZCzjSp3MF
izEz0JET0mi9wnQyoqfrwgG1qPnZshJvAH/F9nbL8+uilbvQ0mR+BjJXwK2xn2fA+aMf+NiNR96v
5VEEfI+sRScO3HRC+IRAGQi6E9TFfAEVn0WjNLrAk7YlfOOKCYu1J57PxnAeooK4KF2OMMOX/FED
yFXNj12yoyCb0KdP0aqLm6hoD581Ppg9/LnTJMd9Y9eJa2MtZd+ajED2QAPeSFysq1/FettLSdjp
JT7NvgH9EHrGAVK2MW9ixFqQSqiMLVIzumeT/sISLXyxdWg65+uac6uU3L2O0+XY3BtB4e2xt0Ix
6uxUDtB6t32bZehHe7INE2Lxgmaq9ci1g9Sy7DyMpu89S5Ih3kG4LfhMGZTJ5ERg2uoI7fehtNcA
Y+L15z9kPSKMOmWCFcZcWUovf5uxNoBF+5erR3F+Gf7KtTjOM10OYVp7YDbG0JTaTGopmQA4LG6Z
WPqaQ0N092TeQhm4zq3hCkIqPHIJBCc9ZNTIirfPMBlQR/UyRDvFRkCnOQQwg9i/OQJpRLqXQids
o8q2QQJi7PIReXsHXmOzatOPNVtM9pCcr7qwt5ty29dSlumMG0pEexR6nkKnokQzji6d4I4RGgQt
dhCuDAssQRpTKUE+ifzatlbHNVRb9tsDL9gTl0ypxznDm7aL6o0WUrfkUBaiUac+KwZTdepNJuQj
riBSffA/H6gRRAIi84P0xE4Bsh3WT2pwTfprO2ErPz3EUpPtHuslOQRJHvYw7e7E/y/EPzx5G4IL
LVJoDXEZAPzHt1x0QyXuMtp3IguUtK52kbBFBqRc8obR+7QY7LafSuBsC/JwDcp9cPdrVVnIXFj5
y5TxYjM9dfT0bbGmkpWhP1eeIclRx2O0XlY15T+zPabaNcnC6PMCp2/PfQ5A2ke1hatILzwHCSqE
Sn0TF/XIRQW5Ldu0H3WLQiYApHJP9z45uqJPP5OOcp5moygq7LJeocb5b7P+lNM09/xgpcJ/6Plw
7s0f/KG2c/hbmyX3U+Ixh8Ahi+vqa7PF3x4/3g9GXxiyzGSCxktvTuYxsyqyHCUysjJhU7XaW21b
ZuZNPwMTUPYVMeJYo26+7UmXUaCtTqRN1PbqByLqkgcGXYKeBrfwFJOpNtr1XiPvwFvAEtdYRhhI
v09EIrUZJDIF1UDZXeNY45u0UITOFwSpZCuYmxW+IPidiVUzFaLfggQFVCe80QaFgxMlw74HG4Vy
k/7hSh8mLGz+0kcGGKmEO+Ee7HErGXz3XEUh3HZjfAiDUTrBRbgd9rCE2uCg/f3PTsYBc7BkqjRk
usfBUHbzyAnmXfFMTNADsq6YxtDC3Gy00c7pliT3UNCvHNPuw8ZcmVmxaGQ8u+UGnBuuPXTsVlWF
kWSssZueNr/AHpsemIziEiqUq+q8tHvamb5tXtH8c0fj2Ohefl9RWC5dKrAGHqEZQyKp4u+e7kvS
KQB5QduRF1+LMC5NEP4oZHrmQCWcm5fJQZ3cmh4y2b7TWFpVz75w/0ku2i/HM/2X/30I6pweqnY8
WoRA5GgLtxC7kxslTQXOcaavwtKomM9o7lXh7cxW3AFMNY8HWxeadQ859sZeY8uln7UJOboF2Ato
ruA1gFAK0Q3yWNOFPgMjDdpWLaHnppckrqbqrhxWA2p/3JvmCuOm8vtfMOCupiZjT3yZcSya3m6U
tgENokPLj0Vade5AnSZt9suIJ71h4h6lDyGGYVotHrJi/VLKIm3ka2Ru91DOHmmeljBwIv7+WXdd
ThgLDoIHsB8pub7ua5RmmLpWu6qwyZEy8KQijoP/KzWvCw8e34DPgUjFhKFHUWYPvoTegfhgKROZ
zqe9E6wvnFzV2gPbUBnHnPX8AMCaCVLa2IeD8mN8qvTFF0gyflDoyeliS82n9DbDg/oX+ZbT9Owy
HkDWBcBxk927nvGoX6v4T1jRKZ3wzLS6AogrJas0pU/aYvHnJvjIXlc/H+Tyg8jxapA6reCxbEwo
VTbxURn0C/xCxNXfQmSfvXwOdUDGfAOXxn2V8RKqn7qmRnyP5ts9Avh7qOJz/LhpkQS66I3qGFld
KOYFAQjbcbqyzFDZIgttzv1ggvQGRjC+5Q3pCHFcIZ2oz1Kx2zV2r8ElVsouG4VgkOKzB4IAgWRh
HkCalCCGzrlQMobqPmLZqrXhjThIV+tmgxLPD6ebrY80YMc5+KrYFZO8AplOIexeMxdxLM8elwzK
3Eo2slq6XHgDtEgHzFSOtq+md7hR+P4vpGX0t/e04985/Rdit+UVxr6eg5RF2Ai9vI7rY+9Uvxkg
MKIdwnSc3HIFs+priSJo7j1G28X6tdCAM5MITd5uRK5cmsgAO4UHLF8Ck+a1ufc+B3tzxfR1Nzwt
jH9DpIMEx/Ezoz9O7pGzPCvLCDm3xJPHSSsNwlrGp5qeOvgFrmGLLmLjbZTsTv2kRb2xz7caYOv6
K2tZMm8g6T69Gl71tJyO8LDhn8l0NLI9xiLX5rwPHtR4iP2INh23wNIv1V/7c1EQBdEARvzWJP2n
CjxAq26nf3SzE0KhHnamLT6ibq8Q6gY4qBig8ha0ZwbRO2jwGGMryPy4b2mDDvATyhSD0s4VVIkS
dnppVW+j7LiXPdVBhMiqxIqfpwalmT7fKCYLvmpyhTw8LQKK8Xr3kYg7/Cxu2ug3WG7SxjYPhzxC
s93end8MxjbBAVyTu4rsDd3oXwsTf+5iIkuLQ9h7eZT66lktydmPiKY8Zs6BfOYhhViD/0qoAPfH
9rzoQD9bC7uixzCtaxgfU+2uPHQN+ZtFeJGgtG7tteC5XunBtpECJuzIsjEXH7b7ObQqn10lQufv
l8WPhxiQcNOXW8vkBxCf38w8A8i92yo7iOtHCLWgtBB5zIV1A8BToKM8tgxURmtze6LbEtYYxRff
//oljWW/ZtYmKtbAsRJuvKXHfneCypx+eYe41UUDuKeI6XpbKvdQRrBk2dHgluUqUFqlmJSW6wR3
BKS7S+PbuREf3rwWmEZzJwha6ouTFGCrPF6iws0d4MVYvi5m4hQcDJTsjUwr84M0A4nTooSSiKdX
bPHmslSHzedEObxqPvbcfRqBhdmZ/v/LGNJIBzWYH8wRWfNmI0lUVNUBA3p2PYbUlAQ7G6EV1Wqg
6k12KrgMWNpKOGu7xHx/Pcf9wbuBu8dTnxz+6v+X5IcAopY8/FTKpvnDZmxc5F8Prq4fKaPTr/en
K7WXZ0GZ8dSSYDeG7cbljX3huoZZ6PDHwwp5pKuoaGNqgd3jOG8aI7Ou36GULkISGO7pwpkP8ZcY
QdcOLRE00cyO2/3BpYB8m8WMx5hKbKrVRpDm1tI0iIlh1leNYrR3qzhQbLYafCyWhG8BshxHhsZM
iG2PdIq7XrOD2/9D2sWXVbOGsB0sSaJRBgy3c40QfEDWCBY89BLXy6vCXOarOS5D/4H3dSH6xvkc
O/xHduK79tRmUcrZXYSzOUOMFsvHbZzqHFuMOuryCsGIRaMP7OBBnSEQrY0fq4dUVdpIIHKb5iH6
1BdPbV0Ws8Tt7MPL8/7qUbpRuzY0wB248HGVWbVzbQUtEK7g9lhJTQCUKzDYPKUrTsXdExp2QUtg
HBdskpJDrszpJ5UAWoWeWqFcVqkaWFOJ6Wx74VqODYCD1o3+s1nobfe2yv//NLyLlg5Giz7FVPq9
Lb3/6Hyeb4gE5HE+jAZoL33SuFfqFVmCDEsWCvWgbW2R3ZgFx0IR7HhCglEhLgdRS0tjI90Mz1Fq
SHlIjUtWpA5Igp26LEHvRpsgv7SKixh1fThyG9BOw1DWiUbnov0TannZaU6ZYZMNy4DIYIwQwyux
fToJHJ3CpnWtfPA4lQqHFVNCOZMjDB7nZvv4aVBuip4ILME6DJ2dJsYCtOKMeiV4EXjSrukceDXb
dhmv5EKrQr+l+i+YzLfTHZyX3SAoXE+MUKnwBKypfY1YLeO3JrqYFKziWEiljBEpGWAdqZOd4/6Q
WEFrrRDiHUuCXbtiRHeYiXSmbWL4U5nrFhR3byLHRQ+tLqbNuxorwYRRVZol2eqw8/0sfezJQNYs
zr7eYkT/D72jgHuySS0e484QHv6h8mrzJCC1itDe0A1+LRYXBMCqSOkeXWM5JQIRZENJ/Iu+mtIb
aTDw5/QY5AX/JEsPudooWRGoMkrGKnMxPUKt/I0UYYmoaPMzZ/ItEUsImlTMXi/hfTzhOizq6CfB
Fmr9TmpudrapJS9uxeI/JZf2+tKD8TUXYLTZR+Krzysjej+a372wKRhcuum8oyB9+GctYlYPsDlN
rD7Xha8pX89A0dSqWcZbzfKGU6kM8/HEiQQtp1MhpqjsqONOeo4vrbqkGvY4pskAfP/aMCpmsrxN
r4xwD5/ge0DaapDfeYuuxpkHE0ohEOlyPD2j4Svp614EhwIHijCJttRvsj9P68DxFIa2SGRpUGK3
kx3MX7wqXO+09bjAGtnYWnShBVE+TDp1lDpcCzrhGPLS3djH6SfVPClSUM073D9b8FSFH5iX4Z8h
w02CIWEosUp32Cp2dYBFkWYp7/BYSIt5VENsxoF8dN+Z/AUonUFc/fPB3D8r8By0+RD6kq8+KSO8
0rkDklnEd80PdJv1mKXwR9A9QEj7Ta/KY71kYs/2R3RxOT2wQroVP6iy/N4T54wfzWmoL7DIojp8
77j9uqN6AcobIgc1E+pfQMkvYsFQXMLrbMYIU5o7kv9W0+bJZcbzTxsz5gl6g3EeIQ3HnhoHPe50
3UkffdVH8SztE4RiJKcqTPTUD7bKgZkgAFHVfnLB8NO1c3Ro7FL4tP6NsTOZgg4SOzdEFvYKc1ps
JnpfVDzh8y2faNwG9E3wQF6XTkfgvD+kEG1XbhWPZLsQCjNji1Q3LeoFIMTfv4TajSCOFY7A2IvC
Kv+dKj+MrG7PXZXHhkNy5tIq5JfOKoUHj1ZMrivRw3+k+gc88Apd9VOc6ajOL6xe8wXlJ0liXdsD
bp4Oyp8uqVq6KTO/SkCxmYdRSKYq68hSJ9MXxLPB07rLRIFd6soHInIZm3Yme1JUW+8YaYZSRhgi
fA1hD+eTWVI/gQ4tZKp761U1rCmpIYmeR4EbetLMiCL277qjO9gqyt6M/ToiGEdFVnGfi5TxC+Xl
MgBMmWxh/4vqkzIaVL8KTTwlcTry3feDQOwEfJTlRu6sbjl1EP9ekh9Ep8o0WkLXFtGvbPSqQhY0
51o4yWQ53qIY26O9Q5WSoFnIlL/BsaPnVV+xGsdvpHiXHYx1yQrl70axiNDI4T08SgBbg1h15ncp
YM+yzlW6+bvaB0pgWiodghVah4yICcaItHLnD0kYiF4xMjAACHuEPVV4sIsMYt+LihwY686GEsta
yJYcIGSRsN1IB8xTFJ8rC7v+sS9c+YbXA1gOUGp/vAwqgumQVxzNyw3wS03GfHS0onuDvsKBDACg
e7+OzT7SRLPpeEGWEVCW44hgQoYBHnKJ2XkXaMlnBE26gh7atSCDNeTZ9rZitW1knkNtbhzhpQYj
RrksTyy0VSJCsB1Y/MpS3bAVXU5eZfUlmudeoci+p1JEWCtHkGS7WGMOtDCtpZpTarUA1KYdaen3
FtMi88kgJrEJt88z0p5BrK8HEU0U7fBHXPOnge3Eb4gLkY3ED6ZASJm+bDLRluLUy71FzT2PdcMI
/NB7Zhb055wyyQE0/zI8AcuCqIJoknmmFJFt8p4Iazj0vYauq5qntYv3guKxxwoA4oLNMUn+PSBP
L5ep/SUe63Zl/zoVmdsouehtDvU8lqK3xgCS9lFYrcTt67bvZWMH0yNmZjvSv7WRX2iyh1DfVsjF
MSkX8QrvKvEOnKT5+DO0JOrnNC8Jm12SfXFeEUMkJ/PSwYD+C4ZSZfIzBykK96TKuiyYaXosJfwJ
h1CqlDpHkHhJXTsd75L89sLJRaKaEPnlX9v1kS8UFn75ncPtJH5h1Lx0ueiRIyr6xhmJnXHktpzH
xI+eFDt0a2gU2sw78IRzu5/b79rxG6j9+UeaaWSBvccDRel5j/G3TeDdxvvD4TsfCAkDqMNFVC+n
CBNebUSjRmpKaCWGaQ+37kkRDneaV9icA9uUdTEWsOMBaD1XbIlyq9eKSrefV5/epYA+bDI/wlvV
rZ5YVVEEHmy38S5BsmZI/4SpM/WN9pz+4GK8BCSaCwpNN/YG0PiKVZVGqG6hWPKEXv9lbwc0RLmZ
TnFPjwphvEDXjI1gZVlirqjzC60T6NOl+T8JUsY8lfWkhegVUhIV+aAB7VxWV1gMkkCjRborDsFp
3PuTEqsUHNTpN03jgivwxICo2otWqmsO8GkfzFEqZSSKLkhaXCCtBN7gensaaAU1Xge1W/FGi/Qk
r9qnLEAIciWdvRJApDABQg5IiS1MNq/LTGKHvssyNuzUJems+SEM7l57NYYzRxvxPnDPEtHEOkc/
z5ITpdC+EKCKD+4G6xZu87FQy14xV3bhTLBYEN6N467QsqGf2QJk9jMUMFIdC4J8WH9ekm9WmQw5
XnJxHctr44h+MQYYL3jLFG7sPM2Wms+PKKJPx7OHhSNCiQDEqHGCsnjBKO4hiUFfDb20ieyh7nKW
jp3GIlwmpXjY0tI9AeIMdHX+JjE26V+B0yN7Z7fgvB7lfSaB4cQ+1qSLYFxk3Prks+fao4DQygUV
KniIMJ1uEe53Dh6t8s4YSTgBTrZJoAketSbUH6dtASX/W3g336OnhWaA7eel2+HjTNZPMjQOmUUG
XKyaq0tlk/RlCIbaIKSnXHpjvdpjt2Pq8BghD1vKn4YWa72M/f4uIy2CosaavRDQF1GqW0PUoUsD
RAruHQ+57td0WZcM6489jp2JFnf1zSd1p+1GpIgJ40s3G2N+e/OOn4SWnOPCCAPBbYcluphioYbp
dfBW/wQ3Yb+TRuIjv0XCItNGPOVwgUVd24VtHIHz3ePtZcOw/ryqxX1Xmg6Kua1jc1YLXjJ7qIP+
PMZ6/NPIogmV3exrRMB7+InUArx0RTIch95QSnC7neeMmPJfNduV+uVn8wV9NT2IJ7sRp6y5IwXi
QJGousnF2ge8aVIPGbQVhwTJjEyE3usUD1PhsRpXyK1gSkm/mMLO1vD+DzCGDi2Bpi+TJ9r1/qG2
K6x0iQ7AQEX/CeFbMcYkFNHwJHIT9tIZr+P80qEbhvHjRyg7lz65TX5M2b+iH2xywOxGzrt59pha
1IcPsuEMeWcjrUe3J3jVWTRBu6Kb2kjKprxQF/GkdY4GQFCHpXgvbAL5Ds2PCva78I7FIhJyClQ+
yjfdIzHJI2D72UetusNA4ro1ONvsJa2pMAmSijTaSBAi6tkrz8+U06lEldDcfPc8AvcvL52LvNMR
pXmrR3suuOv0fLsJo6AocVU3T8DedOsVxdJjjtslcd4+9xxpjmncXazHbfHo2bWAZB60mgRxmAX9
HSpTDK+8cY1ghZ8AgoVGEBsvGkUclp5opKKvnc4yuPupHzykyjVxp1hVixexPpoKIOiYwu9lpO2C
NtwkrK2YJwVVjgQySI9IEnv7jLmqxMpZ5td2kqIn/MU4Zt+GjSEBqht19SMcFlsqt/zewZnWg022
VdY2ewHInp29ZL+69HwO18uafAxaJCDxtbnrTaRTAngtRXaH8OUf1ZC0VjCganVVlsCA3X7GaaQf
F5x/w2u7O16Akziye8wZH7r5HkDYnT0PpdtrZPNAt6xbVx6jGnVqqwttnhnBKj9sv3WgxE9v3OsG
+gbA5GUhnZUvZP5CCXZSAfDFhn7QJEL/+QwUCrOJru/vflMX53UzUP3Sx77v06A5kX1sXb1PHJHa
0nUWXYC1JTObQagfbNjJ4QVHBj4I0yf+Ln5p4UKY0EnVWdjpkhKVbQp3aKOj+J77npKcTJD+0zyx
MBFRqUsvKk5vRKdUeOUprQBqwc2KvbWF4N7qQRYKklZTFHCG38pshykOw+cQtmt/9/XWHfm9l3An
//BoF1wlFGI9obPMFnEd067lkO1SQKtEb0noQYSL+sE7KTwXFvcwwrbHI7j5UNdH4ZXxOC3ODaIH
1HrikDbiHMk6SzEX4kWPTkJS9YPCic7HWcrcUDEVdyx/qb71fSA8R74OU5iHbuVN6qWPTTgl+utu
tdHt64LGUBuWoHQac383uGWsOs44YtROYK2vwfaJtSRYEWh8siLjJy2YVRJv0qoKvqa1Ca/vRSdr
4gw1+BrXBLpox8Iupi6HbK9ybGtwobgs3c8JLMwg1vU8Mgr3jAvTCj+l/vEYVdMLjjXBX16m1b1h
hckuuWpz+GEG1vHfbVwuIotXIq3VVldou8piqyDLp5Sl3nAwIo5OZTBUl7c6u5gc7h8I24IY0PoS
FGVUg1rFwpgzOjjPvfnFn8xkkLUvecBXkDbMnNfscJF3iLuRVUCJO4F/5pGlFfTF4/q63GjFqb5v
0AA4HakxopiarUeuiNP3ODxCPtdjxrKvyFoS1ZwwLoEhOEgxg/VCqKvvCxClbRXOsyJNfqV5zoCM
UxZQ0nfRJdFl9rswJNj4Cy7frdY3Op8ZYZH7z+CcDmHbGS3qXa2z8xNa4d+uGvnPtJFS4xtcKM+3
lgOaTq41XtPYdsCLmg5SSTJzJ1gqQjp3daRnvGJd7xLPyz7J1sJxpXP4fEtVYXP52Zlb0+3bXir5
E9/Co+/wiQvm/DM9JXJaPMqhyK3an2Ac8wM1hHY8vN8HzlaggbiQe/WMg2c+TN7mvwaKV/LTGHeY
xSMJn6XHwzJBM22gsRX5U97svsofXxQikuaDlo7nIHq132XIIDlIaDa2ppLo9kL39VsBMgYvGxzK
kNUUzDckzexSK1TGnJEE+1PS+BjMulafOEE6cYiZygN69QERLFoONfxKF2mVppFUX630Pmugq5fu
W2HSLCH2vyHHwgjDWvw7RRzB+TgsZsc30H6ZiifDGqzulB9mWrszFsS8yTM1MI+M/25gMLUAdOPh
2+A4nTBJ2bawcObRr4hHgoFU5MuivoAU7wPwJbyDqEUM74mGtiY3rlgB9Wjj76GfcebcLkqBcRDB
W9PYDj0ON0bIwOpM1mjuq8ZkjKbhgqOo3BxMUy4o+olpClMKuIIxZ2J8pA1bGjnluwIGrZGeNRrD
nzsgozSWDpcFD7WMrrXqdAJXaFawnaMXVmI1wZz10GQ8HkK6Qd9bTkFuuBVjjifak4/PJwL9MieN
5rT7dFWKVb2tS/NeFzpIB/oxkFpS62N+31S1MtMvNgJKornyj4ThRldcoh1rK79cLpFh8lT/zVGU
9ll8Rw7e4aRX1NYIT1ibkyEamKPVtCYUWq8UbyPksy1+zMhN1PHgWCANs5Dn2nlopY4h9M82Wuc8
/16EFtBgtGwoPsfDereD1zYIICLZmYBb8P6zI1ntJ1jDpY+ZCy6Q/Sx+9RdPVYGzTO0tlhAifo3k
ceMrZo0HZVgDQox6n55gEi61mksqBgy04esF5mcHMqJWGsR68G3rXKOA0UwnrU+nCKdQc3dVEPZI
GT7N/nlKDnghPci9KgqQ7knff4KrBxxjRp3ppCq4vPhaVexGRY7H/Gxen0ib6r7ztzwXNTYJLCYh
7RzS4pieIwS/mVgn7c5NaD1LqUPesnqGcaIi10fnUm17XeMIXpdvCKOxhXZb1PhxsR7mkO3b1BWE
gyP1r9A9+W4Itvav3igb/bFgSzwH05+F6DbkuaeDt3daRrHcoxmP6s/fqq1c8LmVJbminnGLu660
BszzNo/bfjiOphMAXAtuWyzGmJ/2Nqxn/13xtyXgYpMj7koX5p1XFYszwMjm+oh3HN+IinwpWKdb
6505fgybTIiQFR9nfxKJl14DfTCMJe2xomZo9COWQrZeDBluU8wyVx9jm5C1pc7wAua7His5hFGj
EH5ZSz2oMvQmgEXGPS7v+WuItPTEdY2Le0jl9gamxkfATH2e/pO1XoZcuuVZzMgxhXC/DhPYAh3x
GFXsRXkRSxTGCatdLGZfGGpEIw05RetFjhvFuDM5xC3Ooo/Le0gQJnjlGNLB7xUBHf2IdBoY2Jdt
Sqag5OTfZXazTg0KqS29yo/+5YtPBNR4fyZf4/6s9Lq8W7IBokgdU0ECO1Rl5dkQj20BNbdoBM/w
TWQrwLI5EOmtotvQvbTiC4ecazqmc1rBBAyo81pRZPGri+V+tppMxDnRQxWyf1yTeCQHKxl/99Oo
NCJQpNrh16DAUcOvZW10dM8qr2auoT88k/wldLki9MOtahZ6nU9e0Taf3h2NNxRFgT60q1QWsPcl
he+TS2L4pi6zzf8/BwLZqYVE/klcMojOm2zSOXXP6yRHjLrPgvuhaZbaXSnYAH7MGrz7LuHpdnqu
tg2SvT2s9rIabj/Rg7cUNtfV8NX8DpynCXK/IqLW0fKzAFgbRAHGo0t68A7pROE/ALeGjGfS6AFs
+8t8gwalGMOiOkKeGUvgY9dQn7AhFAxbjg9Nyvo48bDn8Z3MyeRuazzBA6PbkRi2bR/piqy7PaBd
fERiBCdbFuB94VY7g/SKJeGIqddIandNEXW9YfOSXcaEm620QFdTOLJouVhK2W441jF4+KWKfmy2
kJIb89WqFvw+9CPXDO+kO6pJIrRhUwPz79jhJqKWyNJIfY6YB5Qj/2b9R5WV2Jk5pLbBKPc/J+EY
vMa5r5+MAVFpcEobLzuyX96flmAy50O/JD/ZqiCYIDf+GZF5poPhWmIKeYFZvYi335YhHGrTbswE
ncFmnfdQOYTQl89AxX2cEf+tDTSFyHeJ54hJCP90o7Yla6sAqS2Fm0SIUp36rPkZlRFIumvuwDWi
ex6UH0qpA1XGWUP6Jgna9P85W2gKfE72Gpw/zUqQhu7ytCs3tpQxAwvO8n8GXe8S6wjd8vjDw8Zm
uRNDCorm+EQpMUk4eZKRqV7lFA4+OtsKuRrH4qL2NuxW7HybO+HC9r7GnhCOjPkLRzvGmc0mEP20
S5bG2LJCha3QYw7JNnYa/ljEUos/PQIHwQOIbRiTr26bFAkcCnfHsSefZ1VIUpy0hy0M6rnbPd1o
ws9MPrFSt+bK0esLWN8TyCzu1qDLmD6zeECG9Yj512OjunqcoVV2M40FcTP5yxx9I5GXQ1Sz/WkS
8S+GzLBCzwqCpo+dwnDJFKwyyfmT/OnkLKefCC3dvY162Iubixc+vq4J8F9P33nrx7a328WU4kxE
eerbaiWVmoD5ki4/VrjYftqr8ZBwolY4Eq3D9Y3oZcZl6YmXHErn7UXruqMuuTVQvrapFQfBiclq
HOE4lZmVUNPFWGqirzRRM2aOlgRCLbhWOEataDsglpL8vYcTh91tRuCcDRfJasM2aHyP9aT/UJTP
wDIq+g3WY4tUB0ZqmdntTlxviY2Ve91sSA1puRtN8FY1WGmlpmzI469eyAyuZPGVdJr+H9J4cdNo
MM6pf661k1J4ff0UaGVKz64225LQjAaeTWOfaigmmZ98tMulGXCkZiBxk3ri30QrVMK3xqjuMX0a
CrO9TVxaxWvpzvP5Lp0vOe+D7Z1q5yJECWyZNpVn69KsvCSWEyHwH5YOqAhV4jNvIziki9/061Va
h9DreeEST5ivofVh6aw8R+0c9/0lbBjmxCU8AwZG01vL5xQfjBqezd/gTLMZpy803tgSBQbg/ZXG
u98boghpK1qvuv5AIaosBVxiVD2YTQgXBAK5IPIoeYoFh/5pERLJw1fW9qL0JK2BJrkNMwK0DPZx
MYvWZLD2OUoLbnucBIvfhuFJZTxHJc2QbH4zWDtjAfuNsM+Db34ZLVQ/YohPWVg+cnTQU7klw7y7
sMNFc7EtZKrx2eg+LRA3iURN2kopwGEqp4uTAv1IbzXDE2t45zdcLvL2n1TB3cw1s1rD3c7gXXKu
Ny38MbCZE/HTsLu63fl5xYqlinUmQnGCMo+cKcw0weI/BYAKznxeCZBZwbtOdm89l+fnq79qz5+j
o/AoDcjp4XOn0BXk5P4bJZZeEZxp/oPYY6MpuVcDHQfPVZji6wBvPfJpleouS7T/lWkno6sWyarp
f8zZeVFl8w==
`protect end_protected

